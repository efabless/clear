module fpga_core (IO_ISOL_N,
    Test_en,
    ccff_head,
    ccff_tail,
    clk,
    prog_clk,
    sc_head,
    sc_tail,
    VPWR,
    VGND,
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR,
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN,
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT);
 input IO_ISOL_N;
 input Test_en;
 input ccff_head;
 output ccff_tail;
 input clk;
 input prog_clk;
 input sc_head;
 output sc_tail;
 input VPWR;
 input VGND;
 output [95:0] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
 input [95:0] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
 output [95:0] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;

 cbx_1__0_ cbx_1__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[17] ),
    .SC_OUT_BOT(\scff_Wires[18] ),
    .bottom_grid_pin_0_(cbx_1__0__0_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__0_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__0_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__0_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__0_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__0_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__0_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__0_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__0_bottom_grid_pin_8_),
    .ccff_head(sb_1__0__0_ccff_tail),
    .ccff_tail(grid_io_bottom_7_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[0] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[5] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__0_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__0_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_7_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_7_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__0_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_7_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_7_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__0_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_7_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_7_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__0_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_7_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_7_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_7_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_7_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__0_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_7_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_7_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__0_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_7_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_7_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__0_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_7_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_7_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__0_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_7_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_7_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__0__0_chanx_right_out[0] ,
    \sb_0__0__0_chanx_right_out[1] ,
    \sb_0__0__0_chanx_right_out[2] ,
    \sb_0__0__0_chanx_right_out[3] ,
    \sb_0__0__0_chanx_right_out[4] ,
    \sb_0__0__0_chanx_right_out[5] ,
    \sb_0__0__0_chanx_right_out[6] ,
    \sb_0__0__0_chanx_right_out[7] ,
    \sb_0__0__0_chanx_right_out[8] ,
    \sb_0__0__0_chanx_right_out[9] ,
    \sb_0__0__0_chanx_right_out[10] ,
    \sb_0__0__0_chanx_right_out[11] ,
    \sb_0__0__0_chanx_right_out[12] ,
    \sb_0__0__0_chanx_right_out[13] ,
    \sb_0__0__0_chanx_right_out[14] ,
    \sb_0__0__0_chanx_right_out[15] ,
    \sb_0__0__0_chanx_right_out[16] ,
    \sb_0__0__0_chanx_right_out[17] ,
    \sb_0__0__0_chanx_right_out[18] ,
    \sb_0__0__0_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__0_chanx_left_out[0] ,
    \cbx_1__0__0_chanx_left_out[1] ,
    \cbx_1__0__0_chanx_left_out[2] ,
    \cbx_1__0__0_chanx_left_out[3] ,
    \cbx_1__0__0_chanx_left_out[4] ,
    \cbx_1__0__0_chanx_left_out[5] ,
    \cbx_1__0__0_chanx_left_out[6] ,
    \cbx_1__0__0_chanx_left_out[7] ,
    \cbx_1__0__0_chanx_left_out[8] ,
    \cbx_1__0__0_chanx_left_out[9] ,
    \cbx_1__0__0_chanx_left_out[10] ,
    \cbx_1__0__0_chanx_left_out[11] ,
    \cbx_1__0__0_chanx_left_out[12] ,
    \cbx_1__0__0_chanx_left_out[13] ,
    \cbx_1__0__0_chanx_left_out[14] ,
    \cbx_1__0__0_chanx_left_out[15] ,
    \cbx_1__0__0_chanx_left_out[16] ,
    \cbx_1__0__0_chanx_left_out[17] ,
    \cbx_1__0__0_chanx_left_out[18] ,
    \cbx_1__0__0_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__0__0_chanx_left_out[0] ,
    \sb_1__0__0_chanx_left_out[1] ,
    \sb_1__0__0_chanx_left_out[2] ,
    \sb_1__0__0_chanx_left_out[3] ,
    \sb_1__0__0_chanx_left_out[4] ,
    \sb_1__0__0_chanx_left_out[5] ,
    \sb_1__0__0_chanx_left_out[6] ,
    \sb_1__0__0_chanx_left_out[7] ,
    \sb_1__0__0_chanx_left_out[8] ,
    \sb_1__0__0_chanx_left_out[9] ,
    \sb_1__0__0_chanx_left_out[10] ,
    \sb_1__0__0_chanx_left_out[11] ,
    \sb_1__0__0_chanx_left_out[12] ,
    \sb_1__0__0_chanx_left_out[13] ,
    \sb_1__0__0_chanx_left_out[14] ,
    \sb_1__0__0_chanx_left_out[15] ,
    \sb_1__0__0_chanx_left_out[16] ,
    \sb_1__0__0_chanx_left_out[17] ,
    \sb_1__0__0_chanx_left_out[18] ,
    \sb_1__0__0_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__0_chanx_right_out[0] ,
    \cbx_1__0__0_chanx_right_out[1] ,
    \cbx_1__0__0_chanx_right_out[2] ,
    \cbx_1__0__0_chanx_right_out[3] ,
    \cbx_1__0__0_chanx_right_out[4] ,
    \cbx_1__0__0_chanx_right_out[5] ,
    \cbx_1__0__0_chanx_right_out[6] ,
    \cbx_1__0__0_chanx_right_out[7] ,
    \cbx_1__0__0_chanx_right_out[8] ,
    \cbx_1__0__0_chanx_right_out[9] ,
    \cbx_1__0__0_chanx_right_out[10] ,
    \cbx_1__0__0_chanx_right_out[11] ,
    \cbx_1__0__0_chanx_right_out[12] ,
    \cbx_1__0__0_chanx_right_out[13] ,
    \cbx_1__0__0_chanx_right_out[14] ,
    \cbx_1__0__0_chanx_right_out[15] ,
    \cbx_1__0__0_chanx_right_out[16] ,
    \cbx_1__0__0_chanx_right_out[17] ,
    \cbx_1__0__0_chanx_right_out[18] ,
    \cbx_1__0__0_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]}));
 cbx_1__1_ cbx_1__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[0] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[0] ),
    .SC_IN_TOP(\scff_Wires[14] ),
    .SC_OUT_BOT(\scff_Wires[15] ),
    .bottom_grid_pin_0_(cbx_1__1__0_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__0_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__0_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__0_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__0_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__0_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__0_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__0_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__0_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__0_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__0_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__0_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__0_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__0_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__0_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__0_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__0_ccff_tail),
    .ccff_tail(cbx_1__1__0_ccff_tail),
    .clk_1_N_out(\clk_1_wires[3] ),
    .clk_1_S_out(\clk_1_wires[4] ),
    .clk_1_W_in(\clk_1_wires[2] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[6] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[4] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[3] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[4] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[2] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__1__0_chanx_right_out[0] ,
    \sb_0__1__0_chanx_right_out[1] ,
    \sb_0__1__0_chanx_right_out[2] ,
    \sb_0__1__0_chanx_right_out[3] ,
    \sb_0__1__0_chanx_right_out[4] ,
    \sb_0__1__0_chanx_right_out[5] ,
    \sb_0__1__0_chanx_right_out[6] ,
    \sb_0__1__0_chanx_right_out[7] ,
    \sb_0__1__0_chanx_right_out[8] ,
    \sb_0__1__0_chanx_right_out[9] ,
    \sb_0__1__0_chanx_right_out[10] ,
    \sb_0__1__0_chanx_right_out[11] ,
    \sb_0__1__0_chanx_right_out[12] ,
    \sb_0__1__0_chanx_right_out[13] ,
    \sb_0__1__0_chanx_right_out[14] ,
    \sb_0__1__0_chanx_right_out[15] ,
    \sb_0__1__0_chanx_right_out[16] ,
    \sb_0__1__0_chanx_right_out[17] ,
    \sb_0__1__0_chanx_right_out[18] ,
    \sb_0__1__0_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__0_chanx_left_out[0] ,
    \cbx_1__1__0_chanx_left_out[1] ,
    \cbx_1__1__0_chanx_left_out[2] ,
    \cbx_1__1__0_chanx_left_out[3] ,
    \cbx_1__1__0_chanx_left_out[4] ,
    \cbx_1__1__0_chanx_left_out[5] ,
    \cbx_1__1__0_chanx_left_out[6] ,
    \cbx_1__1__0_chanx_left_out[7] ,
    \cbx_1__1__0_chanx_left_out[8] ,
    \cbx_1__1__0_chanx_left_out[9] ,
    \cbx_1__1__0_chanx_left_out[10] ,
    \cbx_1__1__0_chanx_left_out[11] ,
    \cbx_1__1__0_chanx_left_out[12] ,
    \cbx_1__1__0_chanx_left_out[13] ,
    \cbx_1__1__0_chanx_left_out[14] ,
    \cbx_1__1__0_chanx_left_out[15] ,
    \cbx_1__1__0_chanx_left_out[16] ,
    \cbx_1__1__0_chanx_left_out[17] ,
    \cbx_1__1__0_chanx_left_out[18] ,
    \cbx_1__1__0_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__0_chanx_left_out[0] ,
    \sb_1__1__0_chanx_left_out[1] ,
    \sb_1__1__0_chanx_left_out[2] ,
    \sb_1__1__0_chanx_left_out[3] ,
    \sb_1__1__0_chanx_left_out[4] ,
    \sb_1__1__0_chanx_left_out[5] ,
    \sb_1__1__0_chanx_left_out[6] ,
    \sb_1__1__0_chanx_left_out[7] ,
    \sb_1__1__0_chanx_left_out[8] ,
    \sb_1__1__0_chanx_left_out[9] ,
    \sb_1__1__0_chanx_left_out[10] ,
    \sb_1__1__0_chanx_left_out[11] ,
    \sb_1__1__0_chanx_left_out[12] ,
    \sb_1__1__0_chanx_left_out[13] ,
    \sb_1__1__0_chanx_left_out[14] ,
    \sb_1__1__0_chanx_left_out[15] ,
    \sb_1__1__0_chanx_left_out[16] ,
    \sb_1__1__0_chanx_left_out[17] ,
    \sb_1__1__0_chanx_left_out[18] ,
    \sb_1__1__0_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__0_chanx_right_out[0] ,
    \cbx_1__1__0_chanx_right_out[1] ,
    \cbx_1__1__0_chanx_right_out[2] ,
    \cbx_1__1__0_chanx_right_out[3] ,
    \cbx_1__1__0_chanx_right_out[4] ,
    \cbx_1__1__0_chanx_right_out[5] ,
    \cbx_1__1__0_chanx_right_out[6] ,
    \cbx_1__1__0_chanx_right_out[7] ,
    \cbx_1__1__0_chanx_right_out[8] ,
    \cbx_1__1__0_chanx_right_out[9] ,
    \cbx_1__1__0_chanx_right_out[10] ,
    \cbx_1__1__0_chanx_right_out[11] ,
    \cbx_1__1__0_chanx_right_out[12] ,
    \cbx_1__1__0_chanx_right_out[13] ,
    \cbx_1__1__0_chanx_right_out[14] ,
    \cbx_1__1__0_chanx_right_out[15] ,
    \cbx_1__1__0_chanx_right_out[16] ,
    \cbx_1__1__0_chanx_right_out[17] ,
    \cbx_1__1__0_chanx_right_out[18] ,
    \cbx_1__1__0_chanx_right_out[19] }));
 cbx_1__1_ cbx_1__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[1] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[1] ),
    .SC_IN_TOP(\scff_Wires[12] ),
    .SC_OUT_BOT(\scff_Wires[13] ),
    .bottom_grid_pin_0_(cbx_1__1__1_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__1_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__1_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__1_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__1_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__1_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__1_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__1_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__1_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__1_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__1_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__1_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__1_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__1_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__1_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__1_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__1_ccff_tail),
    .ccff_tail(cbx_1__1__1_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[11] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[10] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__1__1_chanx_right_out[0] ,
    \sb_0__1__1_chanx_right_out[1] ,
    \sb_0__1__1_chanx_right_out[2] ,
    \sb_0__1__1_chanx_right_out[3] ,
    \sb_0__1__1_chanx_right_out[4] ,
    \sb_0__1__1_chanx_right_out[5] ,
    \sb_0__1__1_chanx_right_out[6] ,
    \sb_0__1__1_chanx_right_out[7] ,
    \sb_0__1__1_chanx_right_out[8] ,
    \sb_0__1__1_chanx_right_out[9] ,
    \sb_0__1__1_chanx_right_out[10] ,
    \sb_0__1__1_chanx_right_out[11] ,
    \sb_0__1__1_chanx_right_out[12] ,
    \sb_0__1__1_chanx_right_out[13] ,
    \sb_0__1__1_chanx_right_out[14] ,
    \sb_0__1__1_chanx_right_out[15] ,
    \sb_0__1__1_chanx_right_out[16] ,
    \sb_0__1__1_chanx_right_out[17] ,
    \sb_0__1__1_chanx_right_out[18] ,
    \sb_0__1__1_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__1_chanx_left_out[0] ,
    \cbx_1__1__1_chanx_left_out[1] ,
    \cbx_1__1__1_chanx_left_out[2] ,
    \cbx_1__1__1_chanx_left_out[3] ,
    \cbx_1__1__1_chanx_left_out[4] ,
    \cbx_1__1__1_chanx_left_out[5] ,
    \cbx_1__1__1_chanx_left_out[6] ,
    \cbx_1__1__1_chanx_left_out[7] ,
    \cbx_1__1__1_chanx_left_out[8] ,
    \cbx_1__1__1_chanx_left_out[9] ,
    \cbx_1__1__1_chanx_left_out[10] ,
    \cbx_1__1__1_chanx_left_out[11] ,
    \cbx_1__1__1_chanx_left_out[12] ,
    \cbx_1__1__1_chanx_left_out[13] ,
    \cbx_1__1__1_chanx_left_out[14] ,
    \cbx_1__1__1_chanx_left_out[15] ,
    \cbx_1__1__1_chanx_left_out[16] ,
    \cbx_1__1__1_chanx_left_out[17] ,
    \cbx_1__1__1_chanx_left_out[18] ,
    \cbx_1__1__1_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__1_chanx_left_out[0] ,
    \sb_1__1__1_chanx_left_out[1] ,
    \sb_1__1__1_chanx_left_out[2] ,
    \sb_1__1__1_chanx_left_out[3] ,
    \sb_1__1__1_chanx_left_out[4] ,
    \sb_1__1__1_chanx_left_out[5] ,
    \sb_1__1__1_chanx_left_out[6] ,
    \sb_1__1__1_chanx_left_out[7] ,
    \sb_1__1__1_chanx_left_out[8] ,
    \sb_1__1__1_chanx_left_out[9] ,
    \sb_1__1__1_chanx_left_out[10] ,
    \sb_1__1__1_chanx_left_out[11] ,
    \sb_1__1__1_chanx_left_out[12] ,
    \sb_1__1__1_chanx_left_out[13] ,
    \sb_1__1__1_chanx_left_out[14] ,
    \sb_1__1__1_chanx_left_out[15] ,
    \sb_1__1__1_chanx_left_out[16] ,
    \sb_1__1__1_chanx_left_out[17] ,
    \sb_1__1__1_chanx_left_out[18] ,
    \sb_1__1__1_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__1_chanx_right_out[0] ,
    \cbx_1__1__1_chanx_right_out[1] ,
    \cbx_1__1__1_chanx_right_out[2] ,
    \cbx_1__1__1_chanx_right_out[3] ,
    \cbx_1__1__1_chanx_right_out[4] ,
    \cbx_1__1__1_chanx_right_out[5] ,
    \cbx_1__1__1_chanx_right_out[6] ,
    \cbx_1__1__1_chanx_right_out[7] ,
    \cbx_1__1__1_chanx_right_out[8] ,
    \cbx_1__1__1_chanx_right_out[9] ,
    \cbx_1__1__1_chanx_right_out[10] ,
    \cbx_1__1__1_chanx_right_out[11] ,
    \cbx_1__1__1_chanx_right_out[12] ,
    \cbx_1__1__1_chanx_right_out[13] ,
    \cbx_1__1__1_chanx_right_out[14] ,
    \cbx_1__1__1_chanx_right_out[15] ,
    \cbx_1__1__1_chanx_right_out[16] ,
    \cbx_1__1__1_chanx_right_out[17] ,
    \cbx_1__1__1_chanx_right_out[18] ,
    \cbx_1__1__1_chanx_right_out[19] }));
 cbx_1__1_ cbx_1__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[2] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[2] ),
    .SC_IN_TOP(\scff_Wires[10] ),
    .SC_OUT_BOT(\scff_Wires[11] ),
    .bottom_grid_pin_0_(cbx_1__1__2_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__2_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__2_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__2_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__2_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__2_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__2_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__2_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__2_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__2_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__2_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__2_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__2_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__2_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__2_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__2_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__2_ccff_tail),
    .ccff_tail(cbx_1__1__2_ccff_tail),
    .clk_1_N_out(\clk_1_wires[10] ),
    .clk_1_S_out(\clk_1_wires[11] ),
    .clk_1_W_in(\clk_1_wires[9] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[16] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[15] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[10] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[11] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[9] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__1__2_chanx_right_out[0] ,
    \sb_0__1__2_chanx_right_out[1] ,
    \sb_0__1__2_chanx_right_out[2] ,
    \sb_0__1__2_chanx_right_out[3] ,
    \sb_0__1__2_chanx_right_out[4] ,
    \sb_0__1__2_chanx_right_out[5] ,
    \sb_0__1__2_chanx_right_out[6] ,
    \sb_0__1__2_chanx_right_out[7] ,
    \sb_0__1__2_chanx_right_out[8] ,
    \sb_0__1__2_chanx_right_out[9] ,
    \sb_0__1__2_chanx_right_out[10] ,
    \sb_0__1__2_chanx_right_out[11] ,
    \sb_0__1__2_chanx_right_out[12] ,
    \sb_0__1__2_chanx_right_out[13] ,
    \sb_0__1__2_chanx_right_out[14] ,
    \sb_0__1__2_chanx_right_out[15] ,
    \sb_0__1__2_chanx_right_out[16] ,
    \sb_0__1__2_chanx_right_out[17] ,
    \sb_0__1__2_chanx_right_out[18] ,
    \sb_0__1__2_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__2_chanx_left_out[0] ,
    \cbx_1__1__2_chanx_left_out[1] ,
    \cbx_1__1__2_chanx_left_out[2] ,
    \cbx_1__1__2_chanx_left_out[3] ,
    \cbx_1__1__2_chanx_left_out[4] ,
    \cbx_1__1__2_chanx_left_out[5] ,
    \cbx_1__1__2_chanx_left_out[6] ,
    \cbx_1__1__2_chanx_left_out[7] ,
    \cbx_1__1__2_chanx_left_out[8] ,
    \cbx_1__1__2_chanx_left_out[9] ,
    \cbx_1__1__2_chanx_left_out[10] ,
    \cbx_1__1__2_chanx_left_out[11] ,
    \cbx_1__1__2_chanx_left_out[12] ,
    \cbx_1__1__2_chanx_left_out[13] ,
    \cbx_1__1__2_chanx_left_out[14] ,
    \cbx_1__1__2_chanx_left_out[15] ,
    \cbx_1__1__2_chanx_left_out[16] ,
    \cbx_1__1__2_chanx_left_out[17] ,
    \cbx_1__1__2_chanx_left_out[18] ,
    \cbx_1__1__2_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__2_chanx_left_out[0] ,
    \sb_1__1__2_chanx_left_out[1] ,
    \sb_1__1__2_chanx_left_out[2] ,
    \sb_1__1__2_chanx_left_out[3] ,
    \sb_1__1__2_chanx_left_out[4] ,
    \sb_1__1__2_chanx_left_out[5] ,
    \sb_1__1__2_chanx_left_out[6] ,
    \sb_1__1__2_chanx_left_out[7] ,
    \sb_1__1__2_chanx_left_out[8] ,
    \sb_1__1__2_chanx_left_out[9] ,
    \sb_1__1__2_chanx_left_out[10] ,
    \sb_1__1__2_chanx_left_out[11] ,
    \sb_1__1__2_chanx_left_out[12] ,
    \sb_1__1__2_chanx_left_out[13] ,
    \sb_1__1__2_chanx_left_out[14] ,
    \sb_1__1__2_chanx_left_out[15] ,
    \sb_1__1__2_chanx_left_out[16] ,
    \sb_1__1__2_chanx_left_out[17] ,
    \sb_1__1__2_chanx_left_out[18] ,
    \sb_1__1__2_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__2_chanx_right_out[0] ,
    \cbx_1__1__2_chanx_right_out[1] ,
    \cbx_1__1__2_chanx_right_out[2] ,
    \cbx_1__1__2_chanx_right_out[3] ,
    \cbx_1__1__2_chanx_right_out[4] ,
    \cbx_1__1__2_chanx_right_out[5] ,
    \cbx_1__1__2_chanx_right_out[6] ,
    \cbx_1__1__2_chanx_right_out[7] ,
    \cbx_1__1__2_chanx_right_out[8] ,
    \cbx_1__1__2_chanx_right_out[9] ,
    \cbx_1__1__2_chanx_right_out[10] ,
    \cbx_1__1__2_chanx_right_out[11] ,
    \cbx_1__1__2_chanx_right_out[12] ,
    \cbx_1__1__2_chanx_right_out[13] ,
    \cbx_1__1__2_chanx_right_out[14] ,
    \cbx_1__1__2_chanx_right_out[15] ,
    \cbx_1__1__2_chanx_right_out[16] ,
    \cbx_1__1__2_chanx_right_out[17] ,
    \cbx_1__1__2_chanx_right_out[18] ,
    \cbx_1__1__2_chanx_right_out[19] }));
 cbx_1__1_ cbx_1__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[3] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[3] ),
    .SC_IN_TOP(\scff_Wires[8] ),
    .SC_OUT_BOT(\scff_Wires[9] ),
    .bottom_grid_pin_0_(cbx_1__1__3_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__3_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__3_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__3_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__3_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__3_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__3_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__3_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__3_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__3_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__3_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__3_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__3_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__3_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__3_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__3_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__3_ccff_tail),
    .ccff_tail(cbx_1__1__3_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[21] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[20] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__1__3_chanx_right_out[0] ,
    \sb_0__1__3_chanx_right_out[1] ,
    \sb_0__1__3_chanx_right_out[2] ,
    \sb_0__1__3_chanx_right_out[3] ,
    \sb_0__1__3_chanx_right_out[4] ,
    \sb_0__1__3_chanx_right_out[5] ,
    \sb_0__1__3_chanx_right_out[6] ,
    \sb_0__1__3_chanx_right_out[7] ,
    \sb_0__1__3_chanx_right_out[8] ,
    \sb_0__1__3_chanx_right_out[9] ,
    \sb_0__1__3_chanx_right_out[10] ,
    \sb_0__1__3_chanx_right_out[11] ,
    \sb_0__1__3_chanx_right_out[12] ,
    \sb_0__1__3_chanx_right_out[13] ,
    \sb_0__1__3_chanx_right_out[14] ,
    \sb_0__1__3_chanx_right_out[15] ,
    \sb_0__1__3_chanx_right_out[16] ,
    \sb_0__1__3_chanx_right_out[17] ,
    \sb_0__1__3_chanx_right_out[18] ,
    \sb_0__1__3_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__3_chanx_left_out[0] ,
    \cbx_1__1__3_chanx_left_out[1] ,
    \cbx_1__1__3_chanx_left_out[2] ,
    \cbx_1__1__3_chanx_left_out[3] ,
    \cbx_1__1__3_chanx_left_out[4] ,
    \cbx_1__1__3_chanx_left_out[5] ,
    \cbx_1__1__3_chanx_left_out[6] ,
    \cbx_1__1__3_chanx_left_out[7] ,
    \cbx_1__1__3_chanx_left_out[8] ,
    \cbx_1__1__3_chanx_left_out[9] ,
    \cbx_1__1__3_chanx_left_out[10] ,
    \cbx_1__1__3_chanx_left_out[11] ,
    \cbx_1__1__3_chanx_left_out[12] ,
    \cbx_1__1__3_chanx_left_out[13] ,
    \cbx_1__1__3_chanx_left_out[14] ,
    \cbx_1__1__3_chanx_left_out[15] ,
    \cbx_1__1__3_chanx_left_out[16] ,
    \cbx_1__1__3_chanx_left_out[17] ,
    \cbx_1__1__3_chanx_left_out[18] ,
    \cbx_1__1__3_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__3_chanx_left_out[0] ,
    \sb_1__1__3_chanx_left_out[1] ,
    \sb_1__1__3_chanx_left_out[2] ,
    \sb_1__1__3_chanx_left_out[3] ,
    \sb_1__1__3_chanx_left_out[4] ,
    \sb_1__1__3_chanx_left_out[5] ,
    \sb_1__1__3_chanx_left_out[6] ,
    \sb_1__1__3_chanx_left_out[7] ,
    \sb_1__1__3_chanx_left_out[8] ,
    \sb_1__1__3_chanx_left_out[9] ,
    \sb_1__1__3_chanx_left_out[10] ,
    \sb_1__1__3_chanx_left_out[11] ,
    \sb_1__1__3_chanx_left_out[12] ,
    \sb_1__1__3_chanx_left_out[13] ,
    \sb_1__1__3_chanx_left_out[14] ,
    \sb_1__1__3_chanx_left_out[15] ,
    \sb_1__1__3_chanx_left_out[16] ,
    \sb_1__1__3_chanx_left_out[17] ,
    \sb_1__1__3_chanx_left_out[18] ,
    \sb_1__1__3_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__3_chanx_right_out[0] ,
    \cbx_1__1__3_chanx_right_out[1] ,
    \cbx_1__1__3_chanx_right_out[2] ,
    \cbx_1__1__3_chanx_right_out[3] ,
    \cbx_1__1__3_chanx_right_out[4] ,
    \cbx_1__1__3_chanx_right_out[5] ,
    \cbx_1__1__3_chanx_right_out[6] ,
    \cbx_1__1__3_chanx_right_out[7] ,
    \cbx_1__1__3_chanx_right_out[8] ,
    \cbx_1__1__3_chanx_right_out[9] ,
    \cbx_1__1__3_chanx_right_out[10] ,
    \cbx_1__1__3_chanx_right_out[11] ,
    \cbx_1__1__3_chanx_right_out[12] ,
    \cbx_1__1__3_chanx_right_out[13] ,
    \cbx_1__1__3_chanx_right_out[14] ,
    \cbx_1__1__3_chanx_right_out[15] ,
    \cbx_1__1__3_chanx_right_out[16] ,
    \cbx_1__1__3_chanx_right_out[17] ,
    \cbx_1__1__3_chanx_right_out[18] ,
    \cbx_1__1__3_chanx_right_out[19] }));
 cbx_1__1_ cbx_1__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[4] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[4] ),
    .SC_IN_TOP(\scff_Wires[6] ),
    .SC_OUT_BOT(\scff_Wires[7] ),
    .bottom_grid_pin_0_(cbx_1__1__4_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__4_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__4_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__4_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__4_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__4_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__4_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__4_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__4_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__4_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__4_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__4_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__4_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__4_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__4_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__4_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__4_ccff_tail),
    .ccff_tail(cbx_1__1__4_ccff_tail),
    .clk_1_N_out(\clk_1_wires[17] ),
    .clk_1_S_out(\clk_1_wires[18] ),
    .clk_1_W_in(\clk_1_wires[16] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[26] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[25] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[17] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[18] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[16] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__1__4_chanx_right_out[0] ,
    \sb_0__1__4_chanx_right_out[1] ,
    \sb_0__1__4_chanx_right_out[2] ,
    \sb_0__1__4_chanx_right_out[3] ,
    \sb_0__1__4_chanx_right_out[4] ,
    \sb_0__1__4_chanx_right_out[5] ,
    \sb_0__1__4_chanx_right_out[6] ,
    \sb_0__1__4_chanx_right_out[7] ,
    \sb_0__1__4_chanx_right_out[8] ,
    \sb_0__1__4_chanx_right_out[9] ,
    \sb_0__1__4_chanx_right_out[10] ,
    \sb_0__1__4_chanx_right_out[11] ,
    \sb_0__1__4_chanx_right_out[12] ,
    \sb_0__1__4_chanx_right_out[13] ,
    \sb_0__1__4_chanx_right_out[14] ,
    \sb_0__1__4_chanx_right_out[15] ,
    \sb_0__1__4_chanx_right_out[16] ,
    \sb_0__1__4_chanx_right_out[17] ,
    \sb_0__1__4_chanx_right_out[18] ,
    \sb_0__1__4_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__4_chanx_left_out[0] ,
    \cbx_1__1__4_chanx_left_out[1] ,
    \cbx_1__1__4_chanx_left_out[2] ,
    \cbx_1__1__4_chanx_left_out[3] ,
    \cbx_1__1__4_chanx_left_out[4] ,
    \cbx_1__1__4_chanx_left_out[5] ,
    \cbx_1__1__4_chanx_left_out[6] ,
    \cbx_1__1__4_chanx_left_out[7] ,
    \cbx_1__1__4_chanx_left_out[8] ,
    \cbx_1__1__4_chanx_left_out[9] ,
    \cbx_1__1__4_chanx_left_out[10] ,
    \cbx_1__1__4_chanx_left_out[11] ,
    \cbx_1__1__4_chanx_left_out[12] ,
    \cbx_1__1__4_chanx_left_out[13] ,
    \cbx_1__1__4_chanx_left_out[14] ,
    \cbx_1__1__4_chanx_left_out[15] ,
    \cbx_1__1__4_chanx_left_out[16] ,
    \cbx_1__1__4_chanx_left_out[17] ,
    \cbx_1__1__4_chanx_left_out[18] ,
    \cbx_1__1__4_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__4_chanx_left_out[0] ,
    \sb_1__1__4_chanx_left_out[1] ,
    \sb_1__1__4_chanx_left_out[2] ,
    \sb_1__1__4_chanx_left_out[3] ,
    \sb_1__1__4_chanx_left_out[4] ,
    \sb_1__1__4_chanx_left_out[5] ,
    \sb_1__1__4_chanx_left_out[6] ,
    \sb_1__1__4_chanx_left_out[7] ,
    \sb_1__1__4_chanx_left_out[8] ,
    \sb_1__1__4_chanx_left_out[9] ,
    \sb_1__1__4_chanx_left_out[10] ,
    \sb_1__1__4_chanx_left_out[11] ,
    \sb_1__1__4_chanx_left_out[12] ,
    \sb_1__1__4_chanx_left_out[13] ,
    \sb_1__1__4_chanx_left_out[14] ,
    \sb_1__1__4_chanx_left_out[15] ,
    \sb_1__1__4_chanx_left_out[16] ,
    \sb_1__1__4_chanx_left_out[17] ,
    \sb_1__1__4_chanx_left_out[18] ,
    \sb_1__1__4_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__4_chanx_right_out[0] ,
    \cbx_1__1__4_chanx_right_out[1] ,
    \cbx_1__1__4_chanx_right_out[2] ,
    \cbx_1__1__4_chanx_right_out[3] ,
    \cbx_1__1__4_chanx_right_out[4] ,
    \cbx_1__1__4_chanx_right_out[5] ,
    \cbx_1__1__4_chanx_right_out[6] ,
    \cbx_1__1__4_chanx_right_out[7] ,
    \cbx_1__1__4_chanx_right_out[8] ,
    \cbx_1__1__4_chanx_right_out[9] ,
    \cbx_1__1__4_chanx_right_out[10] ,
    \cbx_1__1__4_chanx_right_out[11] ,
    \cbx_1__1__4_chanx_right_out[12] ,
    \cbx_1__1__4_chanx_right_out[13] ,
    \cbx_1__1__4_chanx_right_out[14] ,
    \cbx_1__1__4_chanx_right_out[15] ,
    \cbx_1__1__4_chanx_right_out[16] ,
    \cbx_1__1__4_chanx_right_out[17] ,
    \cbx_1__1__4_chanx_right_out[18] ,
    \cbx_1__1__4_chanx_right_out[19] }));
 cbx_1__1_ cbx_1__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[5] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[5] ),
    .SC_IN_TOP(\scff_Wires[4] ),
    .SC_OUT_BOT(\scff_Wires[5] ),
    .bottom_grid_pin_0_(cbx_1__1__5_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__5_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__5_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__5_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__5_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__5_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__5_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__5_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__5_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__5_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__5_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__5_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__5_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__5_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__5_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__5_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__5_ccff_tail),
    .ccff_tail(cbx_1__1__5_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[31] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[30] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__1__5_chanx_right_out[0] ,
    \sb_0__1__5_chanx_right_out[1] ,
    \sb_0__1__5_chanx_right_out[2] ,
    \sb_0__1__5_chanx_right_out[3] ,
    \sb_0__1__5_chanx_right_out[4] ,
    \sb_0__1__5_chanx_right_out[5] ,
    \sb_0__1__5_chanx_right_out[6] ,
    \sb_0__1__5_chanx_right_out[7] ,
    \sb_0__1__5_chanx_right_out[8] ,
    \sb_0__1__5_chanx_right_out[9] ,
    \sb_0__1__5_chanx_right_out[10] ,
    \sb_0__1__5_chanx_right_out[11] ,
    \sb_0__1__5_chanx_right_out[12] ,
    \sb_0__1__5_chanx_right_out[13] ,
    \sb_0__1__5_chanx_right_out[14] ,
    \sb_0__1__5_chanx_right_out[15] ,
    \sb_0__1__5_chanx_right_out[16] ,
    \sb_0__1__5_chanx_right_out[17] ,
    \sb_0__1__5_chanx_right_out[18] ,
    \sb_0__1__5_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__5_chanx_left_out[0] ,
    \cbx_1__1__5_chanx_left_out[1] ,
    \cbx_1__1__5_chanx_left_out[2] ,
    \cbx_1__1__5_chanx_left_out[3] ,
    \cbx_1__1__5_chanx_left_out[4] ,
    \cbx_1__1__5_chanx_left_out[5] ,
    \cbx_1__1__5_chanx_left_out[6] ,
    \cbx_1__1__5_chanx_left_out[7] ,
    \cbx_1__1__5_chanx_left_out[8] ,
    \cbx_1__1__5_chanx_left_out[9] ,
    \cbx_1__1__5_chanx_left_out[10] ,
    \cbx_1__1__5_chanx_left_out[11] ,
    \cbx_1__1__5_chanx_left_out[12] ,
    \cbx_1__1__5_chanx_left_out[13] ,
    \cbx_1__1__5_chanx_left_out[14] ,
    \cbx_1__1__5_chanx_left_out[15] ,
    \cbx_1__1__5_chanx_left_out[16] ,
    \cbx_1__1__5_chanx_left_out[17] ,
    \cbx_1__1__5_chanx_left_out[18] ,
    \cbx_1__1__5_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__5_chanx_left_out[0] ,
    \sb_1__1__5_chanx_left_out[1] ,
    \sb_1__1__5_chanx_left_out[2] ,
    \sb_1__1__5_chanx_left_out[3] ,
    \sb_1__1__5_chanx_left_out[4] ,
    \sb_1__1__5_chanx_left_out[5] ,
    \sb_1__1__5_chanx_left_out[6] ,
    \sb_1__1__5_chanx_left_out[7] ,
    \sb_1__1__5_chanx_left_out[8] ,
    \sb_1__1__5_chanx_left_out[9] ,
    \sb_1__1__5_chanx_left_out[10] ,
    \sb_1__1__5_chanx_left_out[11] ,
    \sb_1__1__5_chanx_left_out[12] ,
    \sb_1__1__5_chanx_left_out[13] ,
    \sb_1__1__5_chanx_left_out[14] ,
    \sb_1__1__5_chanx_left_out[15] ,
    \sb_1__1__5_chanx_left_out[16] ,
    \sb_1__1__5_chanx_left_out[17] ,
    \sb_1__1__5_chanx_left_out[18] ,
    \sb_1__1__5_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__5_chanx_right_out[0] ,
    \cbx_1__1__5_chanx_right_out[1] ,
    \cbx_1__1__5_chanx_right_out[2] ,
    \cbx_1__1__5_chanx_right_out[3] ,
    \cbx_1__1__5_chanx_right_out[4] ,
    \cbx_1__1__5_chanx_right_out[5] ,
    \cbx_1__1__5_chanx_right_out[6] ,
    \cbx_1__1__5_chanx_right_out[7] ,
    \cbx_1__1__5_chanx_right_out[8] ,
    \cbx_1__1__5_chanx_right_out[9] ,
    \cbx_1__1__5_chanx_right_out[10] ,
    \cbx_1__1__5_chanx_right_out[11] ,
    \cbx_1__1__5_chanx_right_out[12] ,
    \cbx_1__1__5_chanx_right_out[13] ,
    \cbx_1__1__5_chanx_right_out[14] ,
    \cbx_1__1__5_chanx_right_out[15] ,
    \cbx_1__1__5_chanx_right_out[16] ,
    \cbx_1__1__5_chanx_right_out[17] ,
    \cbx_1__1__5_chanx_right_out[18] ,
    \cbx_1__1__5_chanx_right_out[19] }));
 cbx_1__1_ cbx_1__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[6] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[6] ),
    .SC_IN_TOP(\scff_Wires[2] ),
    .SC_OUT_BOT(\scff_Wires[3] ),
    .bottom_grid_pin_0_(cbx_1__1__6_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__6_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__6_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__6_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__6_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__6_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__6_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__6_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__6_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__6_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__6_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__6_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__6_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__6_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__6_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__6_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__6_ccff_tail),
    .ccff_tail(cbx_1__1__6_ccff_tail),
    .clk_1_N_out(\clk_1_wires[24] ),
    .clk_1_S_out(\clk_1_wires[25] ),
    .clk_1_W_in(\clk_1_wires[23] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[36] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[35] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[24] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[25] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[23] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__1__6_chanx_right_out[0] ,
    \sb_0__1__6_chanx_right_out[1] ,
    \sb_0__1__6_chanx_right_out[2] ,
    \sb_0__1__6_chanx_right_out[3] ,
    \sb_0__1__6_chanx_right_out[4] ,
    \sb_0__1__6_chanx_right_out[5] ,
    \sb_0__1__6_chanx_right_out[6] ,
    \sb_0__1__6_chanx_right_out[7] ,
    \sb_0__1__6_chanx_right_out[8] ,
    \sb_0__1__6_chanx_right_out[9] ,
    \sb_0__1__6_chanx_right_out[10] ,
    \sb_0__1__6_chanx_right_out[11] ,
    \sb_0__1__6_chanx_right_out[12] ,
    \sb_0__1__6_chanx_right_out[13] ,
    \sb_0__1__6_chanx_right_out[14] ,
    \sb_0__1__6_chanx_right_out[15] ,
    \sb_0__1__6_chanx_right_out[16] ,
    \sb_0__1__6_chanx_right_out[17] ,
    \sb_0__1__6_chanx_right_out[18] ,
    \sb_0__1__6_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__6_chanx_left_out[0] ,
    \cbx_1__1__6_chanx_left_out[1] ,
    \cbx_1__1__6_chanx_left_out[2] ,
    \cbx_1__1__6_chanx_left_out[3] ,
    \cbx_1__1__6_chanx_left_out[4] ,
    \cbx_1__1__6_chanx_left_out[5] ,
    \cbx_1__1__6_chanx_left_out[6] ,
    \cbx_1__1__6_chanx_left_out[7] ,
    \cbx_1__1__6_chanx_left_out[8] ,
    \cbx_1__1__6_chanx_left_out[9] ,
    \cbx_1__1__6_chanx_left_out[10] ,
    \cbx_1__1__6_chanx_left_out[11] ,
    \cbx_1__1__6_chanx_left_out[12] ,
    \cbx_1__1__6_chanx_left_out[13] ,
    \cbx_1__1__6_chanx_left_out[14] ,
    \cbx_1__1__6_chanx_left_out[15] ,
    \cbx_1__1__6_chanx_left_out[16] ,
    \cbx_1__1__6_chanx_left_out[17] ,
    \cbx_1__1__6_chanx_left_out[18] ,
    \cbx_1__1__6_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__6_chanx_left_out[0] ,
    \sb_1__1__6_chanx_left_out[1] ,
    \sb_1__1__6_chanx_left_out[2] ,
    \sb_1__1__6_chanx_left_out[3] ,
    \sb_1__1__6_chanx_left_out[4] ,
    \sb_1__1__6_chanx_left_out[5] ,
    \sb_1__1__6_chanx_left_out[6] ,
    \sb_1__1__6_chanx_left_out[7] ,
    \sb_1__1__6_chanx_left_out[8] ,
    \sb_1__1__6_chanx_left_out[9] ,
    \sb_1__1__6_chanx_left_out[10] ,
    \sb_1__1__6_chanx_left_out[11] ,
    \sb_1__1__6_chanx_left_out[12] ,
    \sb_1__1__6_chanx_left_out[13] ,
    \sb_1__1__6_chanx_left_out[14] ,
    \sb_1__1__6_chanx_left_out[15] ,
    \sb_1__1__6_chanx_left_out[16] ,
    \sb_1__1__6_chanx_left_out[17] ,
    \sb_1__1__6_chanx_left_out[18] ,
    \sb_1__1__6_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__6_chanx_right_out[0] ,
    \cbx_1__1__6_chanx_right_out[1] ,
    \cbx_1__1__6_chanx_right_out[2] ,
    \cbx_1__1__6_chanx_right_out[3] ,
    \cbx_1__1__6_chanx_right_out[4] ,
    \cbx_1__1__6_chanx_right_out[5] ,
    \cbx_1__1__6_chanx_right_out[6] ,
    \cbx_1__1__6_chanx_right_out[7] ,
    \cbx_1__1__6_chanx_right_out[8] ,
    \cbx_1__1__6_chanx_right_out[9] ,
    \cbx_1__1__6_chanx_right_out[10] ,
    \cbx_1__1__6_chanx_right_out[11] ,
    \cbx_1__1__6_chanx_right_out[12] ,
    \cbx_1__1__6_chanx_right_out[13] ,
    \cbx_1__1__6_chanx_right_out[14] ,
    \cbx_1__1__6_chanx_right_out[15] ,
    \cbx_1__1__6_chanx_right_out[16] ,
    \cbx_1__1__6_chanx_right_out[17] ,
    \cbx_1__1__6_chanx_right_out[18] ,
    \cbx_1__1__6_chanx_right_out[19] }));
 cbx_1__2_ cbx_1__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[0] ),
    .SC_OUT_BOT(\scff_Wires[1] ),
    .bottom_grid_pin_0_(cbx_1__8__0_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__0_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__0_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__0_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__0_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__0_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__0_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__0_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__0_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__0_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__0_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__0_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__0_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__0_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__0_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__0_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__0_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_0_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_0_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_1__8__0_ccff_tail),
    .ccff_tail(grid_io_top_0_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]),
    .prog_clk_0_S_in(\prog_clk_0_wires[39] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[42] ),
    .top_grid_pin_0_(cbx_1__8__0_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_0__8__0_chanx_right_out[0] ,
    \sb_0__8__0_chanx_right_out[1] ,
    \sb_0__8__0_chanx_right_out[2] ,
    \sb_0__8__0_chanx_right_out[3] ,
    \sb_0__8__0_chanx_right_out[4] ,
    \sb_0__8__0_chanx_right_out[5] ,
    \sb_0__8__0_chanx_right_out[6] ,
    \sb_0__8__0_chanx_right_out[7] ,
    \sb_0__8__0_chanx_right_out[8] ,
    \sb_0__8__0_chanx_right_out[9] ,
    \sb_0__8__0_chanx_right_out[10] ,
    \sb_0__8__0_chanx_right_out[11] ,
    \sb_0__8__0_chanx_right_out[12] ,
    \sb_0__8__0_chanx_right_out[13] ,
    \sb_0__8__0_chanx_right_out[14] ,
    \sb_0__8__0_chanx_right_out[15] ,
    \sb_0__8__0_chanx_right_out[16] ,
    \sb_0__8__0_chanx_right_out[17] ,
    \sb_0__8__0_chanx_right_out[18] ,
    \sb_0__8__0_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__0_chanx_left_out[0] ,
    \cbx_1__8__0_chanx_left_out[1] ,
    \cbx_1__8__0_chanx_left_out[2] ,
    \cbx_1__8__0_chanx_left_out[3] ,
    \cbx_1__8__0_chanx_left_out[4] ,
    \cbx_1__8__0_chanx_left_out[5] ,
    \cbx_1__8__0_chanx_left_out[6] ,
    \cbx_1__8__0_chanx_left_out[7] ,
    \cbx_1__8__0_chanx_left_out[8] ,
    \cbx_1__8__0_chanx_left_out[9] ,
    \cbx_1__8__0_chanx_left_out[10] ,
    \cbx_1__8__0_chanx_left_out[11] ,
    \cbx_1__8__0_chanx_left_out[12] ,
    \cbx_1__8__0_chanx_left_out[13] ,
    \cbx_1__8__0_chanx_left_out[14] ,
    \cbx_1__8__0_chanx_left_out[15] ,
    \cbx_1__8__0_chanx_left_out[16] ,
    \cbx_1__8__0_chanx_left_out[17] ,
    \cbx_1__8__0_chanx_left_out[18] ,
    \cbx_1__8__0_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__8__0_chanx_left_out[0] ,
    \sb_1__8__0_chanx_left_out[1] ,
    \sb_1__8__0_chanx_left_out[2] ,
    \sb_1__8__0_chanx_left_out[3] ,
    \sb_1__8__0_chanx_left_out[4] ,
    \sb_1__8__0_chanx_left_out[5] ,
    \sb_1__8__0_chanx_left_out[6] ,
    \sb_1__8__0_chanx_left_out[7] ,
    \sb_1__8__0_chanx_left_out[8] ,
    \sb_1__8__0_chanx_left_out[9] ,
    \sb_1__8__0_chanx_left_out[10] ,
    \sb_1__8__0_chanx_left_out[11] ,
    \sb_1__8__0_chanx_left_out[12] ,
    \sb_1__8__0_chanx_left_out[13] ,
    \sb_1__8__0_chanx_left_out[14] ,
    \sb_1__8__0_chanx_left_out[15] ,
    \sb_1__8__0_chanx_left_out[16] ,
    \sb_1__8__0_chanx_left_out[17] ,
    \sb_1__8__0_chanx_left_out[18] ,
    \sb_1__8__0_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__0_chanx_right_out[0] ,
    \cbx_1__8__0_chanx_right_out[1] ,
    \cbx_1__8__0_chanx_right_out[2] ,
    \cbx_1__8__0_chanx_right_out[3] ,
    \cbx_1__8__0_chanx_right_out[4] ,
    \cbx_1__8__0_chanx_right_out[5] ,
    \cbx_1__8__0_chanx_right_out[6] ,
    \cbx_1__8__0_chanx_right_out[7] ,
    \cbx_1__8__0_chanx_right_out[8] ,
    \cbx_1__8__0_chanx_right_out[9] ,
    \cbx_1__8__0_chanx_right_out[10] ,
    \cbx_1__8__0_chanx_right_out[11] ,
    \cbx_1__8__0_chanx_right_out[12] ,
    \cbx_1__8__0_chanx_right_out[13] ,
    \cbx_1__8__0_chanx_right_out[14] ,
    \cbx_1__8__0_chanx_right_out[15] ,
    \cbx_1__8__0_chanx_right_out[16] ,
    \cbx_1__8__0_chanx_right_out[17] ,
    \cbx_1__8__0_chanx_right_out[18] ,
    \cbx_1__8__0_chanx_right_out[19] }));
 cbx_1__0_ cbx_2__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[19] ),
    .SC_OUT_TOP(\scff_Wires[20] ),
    .bottom_grid_pin_0_(cbx_1__0__1_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__1_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__1_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__1_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__1_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__1_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__1_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__1_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__1_bottom_grid_pin_8_),
    .ccff_head(sb_1__0__1_ccff_tail),
    .ccff_tail(grid_io_bottom_6_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[43] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__1_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__1_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_6_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_6_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__1_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_6_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_6_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__1_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_6_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_6_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__1_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_6_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_6_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_6_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_6_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__1_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_6_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_6_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__1_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_6_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_6_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__1_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_6_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_6_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__1_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_6_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_6_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__0__0_chanx_right_out[0] ,
    \sb_1__0__0_chanx_right_out[1] ,
    \sb_1__0__0_chanx_right_out[2] ,
    \sb_1__0__0_chanx_right_out[3] ,
    \sb_1__0__0_chanx_right_out[4] ,
    \sb_1__0__0_chanx_right_out[5] ,
    \sb_1__0__0_chanx_right_out[6] ,
    \sb_1__0__0_chanx_right_out[7] ,
    \sb_1__0__0_chanx_right_out[8] ,
    \sb_1__0__0_chanx_right_out[9] ,
    \sb_1__0__0_chanx_right_out[10] ,
    \sb_1__0__0_chanx_right_out[11] ,
    \sb_1__0__0_chanx_right_out[12] ,
    \sb_1__0__0_chanx_right_out[13] ,
    \sb_1__0__0_chanx_right_out[14] ,
    \sb_1__0__0_chanx_right_out[15] ,
    \sb_1__0__0_chanx_right_out[16] ,
    \sb_1__0__0_chanx_right_out[17] ,
    \sb_1__0__0_chanx_right_out[18] ,
    \sb_1__0__0_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__1_chanx_left_out[0] ,
    \cbx_1__0__1_chanx_left_out[1] ,
    \cbx_1__0__1_chanx_left_out[2] ,
    \cbx_1__0__1_chanx_left_out[3] ,
    \cbx_1__0__1_chanx_left_out[4] ,
    \cbx_1__0__1_chanx_left_out[5] ,
    \cbx_1__0__1_chanx_left_out[6] ,
    \cbx_1__0__1_chanx_left_out[7] ,
    \cbx_1__0__1_chanx_left_out[8] ,
    \cbx_1__0__1_chanx_left_out[9] ,
    \cbx_1__0__1_chanx_left_out[10] ,
    \cbx_1__0__1_chanx_left_out[11] ,
    \cbx_1__0__1_chanx_left_out[12] ,
    \cbx_1__0__1_chanx_left_out[13] ,
    \cbx_1__0__1_chanx_left_out[14] ,
    \cbx_1__0__1_chanx_left_out[15] ,
    \cbx_1__0__1_chanx_left_out[16] ,
    \cbx_1__0__1_chanx_left_out[17] ,
    \cbx_1__0__1_chanx_left_out[18] ,
    \cbx_1__0__1_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__0__1_chanx_left_out[0] ,
    \sb_1__0__1_chanx_left_out[1] ,
    \sb_1__0__1_chanx_left_out[2] ,
    \sb_1__0__1_chanx_left_out[3] ,
    \sb_1__0__1_chanx_left_out[4] ,
    \sb_1__0__1_chanx_left_out[5] ,
    \sb_1__0__1_chanx_left_out[6] ,
    \sb_1__0__1_chanx_left_out[7] ,
    \sb_1__0__1_chanx_left_out[8] ,
    \sb_1__0__1_chanx_left_out[9] ,
    \sb_1__0__1_chanx_left_out[10] ,
    \sb_1__0__1_chanx_left_out[11] ,
    \sb_1__0__1_chanx_left_out[12] ,
    \sb_1__0__1_chanx_left_out[13] ,
    \sb_1__0__1_chanx_left_out[14] ,
    \sb_1__0__1_chanx_left_out[15] ,
    \sb_1__0__1_chanx_left_out[16] ,
    \sb_1__0__1_chanx_left_out[17] ,
    \sb_1__0__1_chanx_left_out[18] ,
    \sb_1__0__1_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__1_chanx_right_out[0] ,
    \cbx_1__0__1_chanx_right_out[1] ,
    \cbx_1__0__1_chanx_right_out[2] ,
    \cbx_1__0__1_chanx_right_out[3] ,
    \cbx_1__0__1_chanx_right_out[4] ,
    \cbx_1__0__1_chanx_right_out[5] ,
    \cbx_1__0__1_chanx_right_out[6] ,
    \cbx_1__0__1_chanx_right_out[7] ,
    \cbx_1__0__1_chanx_right_out[8] ,
    \cbx_1__0__1_chanx_right_out[9] ,
    \cbx_1__0__1_chanx_right_out[10] ,
    \cbx_1__0__1_chanx_right_out[11] ,
    \cbx_1__0__1_chanx_right_out[12] ,
    \cbx_1__0__1_chanx_right_out[13] ,
    \cbx_1__0__1_chanx_right_out[14] ,
    \cbx_1__0__1_chanx_right_out[15] ,
    \cbx_1__0__1_chanx_right_out[16] ,
    \cbx_1__0__1_chanx_right_out[17] ,
    \cbx_1__0__1_chanx_right_out[18] ,
    \cbx_1__0__1_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]}));
 cbx_1__1_ cbx_2__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[7] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[7] ),
    .SC_IN_BOT(\scff_Wires[21] ),
    .SC_OUT_TOP(\scff_Wires[22] ),
    .bottom_grid_pin_0_(cbx_1__1__7_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__7_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__7_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__7_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__7_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__7_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__7_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__7_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__7_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__7_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__7_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__7_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__7_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__7_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__7_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__7_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__7_ccff_tail),
    .ccff_tail(cbx_1__1__7_ccff_tail),
    .clk_1_N_out(\clk_1_wires[5] ),
    .clk_1_S_out(\clk_1_wires[6] ),
    .clk_1_W_in(\clk_1_wires[1] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[46] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[5] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[6] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[1] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__0_chanx_right_out[0] ,
    \sb_1__1__0_chanx_right_out[1] ,
    \sb_1__1__0_chanx_right_out[2] ,
    \sb_1__1__0_chanx_right_out[3] ,
    \sb_1__1__0_chanx_right_out[4] ,
    \sb_1__1__0_chanx_right_out[5] ,
    \sb_1__1__0_chanx_right_out[6] ,
    \sb_1__1__0_chanx_right_out[7] ,
    \sb_1__1__0_chanx_right_out[8] ,
    \sb_1__1__0_chanx_right_out[9] ,
    \sb_1__1__0_chanx_right_out[10] ,
    \sb_1__1__0_chanx_right_out[11] ,
    \sb_1__1__0_chanx_right_out[12] ,
    \sb_1__1__0_chanx_right_out[13] ,
    \sb_1__1__0_chanx_right_out[14] ,
    \sb_1__1__0_chanx_right_out[15] ,
    \sb_1__1__0_chanx_right_out[16] ,
    \sb_1__1__0_chanx_right_out[17] ,
    \sb_1__1__0_chanx_right_out[18] ,
    \sb_1__1__0_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__7_chanx_left_out[0] ,
    \cbx_1__1__7_chanx_left_out[1] ,
    \cbx_1__1__7_chanx_left_out[2] ,
    \cbx_1__1__7_chanx_left_out[3] ,
    \cbx_1__1__7_chanx_left_out[4] ,
    \cbx_1__1__7_chanx_left_out[5] ,
    \cbx_1__1__7_chanx_left_out[6] ,
    \cbx_1__1__7_chanx_left_out[7] ,
    \cbx_1__1__7_chanx_left_out[8] ,
    \cbx_1__1__7_chanx_left_out[9] ,
    \cbx_1__1__7_chanx_left_out[10] ,
    \cbx_1__1__7_chanx_left_out[11] ,
    \cbx_1__1__7_chanx_left_out[12] ,
    \cbx_1__1__7_chanx_left_out[13] ,
    \cbx_1__1__7_chanx_left_out[14] ,
    \cbx_1__1__7_chanx_left_out[15] ,
    \cbx_1__1__7_chanx_left_out[16] ,
    \cbx_1__1__7_chanx_left_out[17] ,
    \cbx_1__1__7_chanx_left_out[18] ,
    \cbx_1__1__7_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__7_chanx_left_out[0] ,
    \sb_1__1__7_chanx_left_out[1] ,
    \sb_1__1__7_chanx_left_out[2] ,
    \sb_1__1__7_chanx_left_out[3] ,
    \sb_1__1__7_chanx_left_out[4] ,
    \sb_1__1__7_chanx_left_out[5] ,
    \sb_1__1__7_chanx_left_out[6] ,
    \sb_1__1__7_chanx_left_out[7] ,
    \sb_1__1__7_chanx_left_out[8] ,
    \sb_1__1__7_chanx_left_out[9] ,
    \sb_1__1__7_chanx_left_out[10] ,
    \sb_1__1__7_chanx_left_out[11] ,
    \sb_1__1__7_chanx_left_out[12] ,
    \sb_1__1__7_chanx_left_out[13] ,
    \sb_1__1__7_chanx_left_out[14] ,
    \sb_1__1__7_chanx_left_out[15] ,
    \sb_1__1__7_chanx_left_out[16] ,
    \sb_1__1__7_chanx_left_out[17] ,
    \sb_1__1__7_chanx_left_out[18] ,
    \sb_1__1__7_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__7_chanx_right_out[0] ,
    \cbx_1__1__7_chanx_right_out[1] ,
    \cbx_1__1__7_chanx_right_out[2] ,
    \cbx_1__1__7_chanx_right_out[3] ,
    \cbx_1__1__7_chanx_right_out[4] ,
    \cbx_1__1__7_chanx_right_out[5] ,
    \cbx_1__1__7_chanx_right_out[6] ,
    \cbx_1__1__7_chanx_right_out[7] ,
    \cbx_1__1__7_chanx_right_out[8] ,
    \cbx_1__1__7_chanx_right_out[9] ,
    \cbx_1__1__7_chanx_right_out[10] ,
    \cbx_1__1__7_chanx_right_out[11] ,
    \cbx_1__1__7_chanx_right_out[12] ,
    \cbx_1__1__7_chanx_right_out[13] ,
    \cbx_1__1__7_chanx_right_out[14] ,
    \cbx_1__1__7_chanx_right_out[15] ,
    \cbx_1__1__7_chanx_right_out[16] ,
    \cbx_1__1__7_chanx_right_out[17] ,
    \cbx_1__1__7_chanx_right_out[18] ,
    \cbx_1__1__7_chanx_right_out[19] }));
 cbx_1__1_ cbx_2__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[8] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[8] ),
    .SC_IN_BOT(\scff_Wires[23] ),
    .SC_OUT_TOP(\scff_Wires[24] ),
    .bottom_grid_pin_0_(cbx_1__1__8_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__8_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__8_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__8_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__8_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__8_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__8_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__8_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__8_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__8_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__8_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__8_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__8_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__8_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__8_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__8_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__8_ccff_tail),
    .ccff_tail(cbx_1__1__8_ccff_tail),
    .clk_2_W_in(\clk_2_wires[3] ),
    .clk_2_W_out(\clk_2_wires[4] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[49] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[3] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[4] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__1_chanx_right_out[0] ,
    \sb_1__1__1_chanx_right_out[1] ,
    \sb_1__1__1_chanx_right_out[2] ,
    \sb_1__1__1_chanx_right_out[3] ,
    \sb_1__1__1_chanx_right_out[4] ,
    \sb_1__1__1_chanx_right_out[5] ,
    \sb_1__1__1_chanx_right_out[6] ,
    \sb_1__1__1_chanx_right_out[7] ,
    \sb_1__1__1_chanx_right_out[8] ,
    \sb_1__1__1_chanx_right_out[9] ,
    \sb_1__1__1_chanx_right_out[10] ,
    \sb_1__1__1_chanx_right_out[11] ,
    \sb_1__1__1_chanx_right_out[12] ,
    \sb_1__1__1_chanx_right_out[13] ,
    \sb_1__1__1_chanx_right_out[14] ,
    \sb_1__1__1_chanx_right_out[15] ,
    \sb_1__1__1_chanx_right_out[16] ,
    \sb_1__1__1_chanx_right_out[17] ,
    \sb_1__1__1_chanx_right_out[18] ,
    \sb_1__1__1_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__8_chanx_left_out[0] ,
    \cbx_1__1__8_chanx_left_out[1] ,
    \cbx_1__1__8_chanx_left_out[2] ,
    \cbx_1__1__8_chanx_left_out[3] ,
    \cbx_1__1__8_chanx_left_out[4] ,
    \cbx_1__1__8_chanx_left_out[5] ,
    \cbx_1__1__8_chanx_left_out[6] ,
    \cbx_1__1__8_chanx_left_out[7] ,
    \cbx_1__1__8_chanx_left_out[8] ,
    \cbx_1__1__8_chanx_left_out[9] ,
    \cbx_1__1__8_chanx_left_out[10] ,
    \cbx_1__1__8_chanx_left_out[11] ,
    \cbx_1__1__8_chanx_left_out[12] ,
    \cbx_1__1__8_chanx_left_out[13] ,
    \cbx_1__1__8_chanx_left_out[14] ,
    \cbx_1__1__8_chanx_left_out[15] ,
    \cbx_1__1__8_chanx_left_out[16] ,
    \cbx_1__1__8_chanx_left_out[17] ,
    \cbx_1__1__8_chanx_left_out[18] ,
    \cbx_1__1__8_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__8_chanx_left_out[0] ,
    \sb_1__1__8_chanx_left_out[1] ,
    \sb_1__1__8_chanx_left_out[2] ,
    \sb_1__1__8_chanx_left_out[3] ,
    \sb_1__1__8_chanx_left_out[4] ,
    \sb_1__1__8_chanx_left_out[5] ,
    \sb_1__1__8_chanx_left_out[6] ,
    \sb_1__1__8_chanx_left_out[7] ,
    \sb_1__1__8_chanx_left_out[8] ,
    \sb_1__1__8_chanx_left_out[9] ,
    \sb_1__1__8_chanx_left_out[10] ,
    \sb_1__1__8_chanx_left_out[11] ,
    \sb_1__1__8_chanx_left_out[12] ,
    \sb_1__1__8_chanx_left_out[13] ,
    \sb_1__1__8_chanx_left_out[14] ,
    \sb_1__1__8_chanx_left_out[15] ,
    \sb_1__1__8_chanx_left_out[16] ,
    \sb_1__1__8_chanx_left_out[17] ,
    \sb_1__1__8_chanx_left_out[18] ,
    \sb_1__1__8_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__8_chanx_right_out[0] ,
    \cbx_1__1__8_chanx_right_out[1] ,
    \cbx_1__1__8_chanx_right_out[2] ,
    \cbx_1__1__8_chanx_right_out[3] ,
    \cbx_1__1__8_chanx_right_out[4] ,
    \cbx_1__1__8_chanx_right_out[5] ,
    \cbx_1__1__8_chanx_right_out[6] ,
    \cbx_1__1__8_chanx_right_out[7] ,
    \cbx_1__1__8_chanx_right_out[8] ,
    \cbx_1__1__8_chanx_right_out[9] ,
    \cbx_1__1__8_chanx_right_out[10] ,
    \cbx_1__1__8_chanx_right_out[11] ,
    \cbx_1__1__8_chanx_right_out[12] ,
    \cbx_1__1__8_chanx_right_out[13] ,
    \cbx_1__1__8_chanx_right_out[14] ,
    \cbx_1__1__8_chanx_right_out[15] ,
    \cbx_1__1__8_chanx_right_out[16] ,
    \cbx_1__1__8_chanx_right_out[17] ,
    \cbx_1__1__8_chanx_right_out[18] ,
    \cbx_1__1__8_chanx_right_out[19] }));
 cbx_1__1_ cbx_2__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[9] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[9] ),
    .SC_IN_BOT(\scff_Wires[25] ),
    .SC_OUT_TOP(\scff_Wires[26] ),
    .bottom_grid_pin_0_(cbx_1__1__9_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__9_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__9_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__9_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__9_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__9_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__9_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__9_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__9_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__9_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__9_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__9_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__9_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__9_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__9_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__9_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__9_ccff_tail),
    .ccff_tail(cbx_1__1__9_ccff_tail),
    .clk_1_N_out(\clk_1_wires[12] ),
    .clk_1_S_out(\clk_1_wires[13] ),
    .clk_1_W_in(\clk_1_wires[8] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[52] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[12] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[13] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[8] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__2_chanx_right_out[0] ,
    \sb_1__1__2_chanx_right_out[1] ,
    \sb_1__1__2_chanx_right_out[2] ,
    \sb_1__1__2_chanx_right_out[3] ,
    \sb_1__1__2_chanx_right_out[4] ,
    \sb_1__1__2_chanx_right_out[5] ,
    \sb_1__1__2_chanx_right_out[6] ,
    \sb_1__1__2_chanx_right_out[7] ,
    \sb_1__1__2_chanx_right_out[8] ,
    \sb_1__1__2_chanx_right_out[9] ,
    \sb_1__1__2_chanx_right_out[10] ,
    \sb_1__1__2_chanx_right_out[11] ,
    \sb_1__1__2_chanx_right_out[12] ,
    \sb_1__1__2_chanx_right_out[13] ,
    \sb_1__1__2_chanx_right_out[14] ,
    \sb_1__1__2_chanx_right_out[15] ,
    \sb_1__1__2_chanx_right_out[16] ,
    \sb_1__1__2_chanx_right_out[17] ,
    \sb_1__1__2_chanx_right_out[18] ,
    \sb_1__1__2_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__9_chanx_left_out[0] ,
    \cbx_1__1__9_chanx_left_out[1] ,
    \cbx_1__1__9_chanx_left_out[2] ,
    \cbx_1__1__9_chanx_left_out[3] ,
    \cbx_1__1__9_chanx_left_out[4] ,
    \cbx_1__1__9_chanx_left_out[5] ,
    \cbx_1__1__9_chanx_left_out[6] ,
    \cbx_1__1__9_chanx_left_out[7] ,
    \cbx_1__1__9_chanx_left_out[8] ,
    \cbx_1__1__9_chanx_left_out[9] ,
    \cbx_1__1__9_chanx_left_out[10] ,
    \cbx_1__1__9_chanx_left_out[11] ,
    \cbx_1__1__9_chanx_left_out[12] ,
    \cbx_1__1__9_chanx_left_out[13] ,
    \cbx_1__1__9_chanx_left_out[14] ,
    \cbx_1__1__9_chanx_left_out[15] ,
    \cbx_1__1__9_chanx_left_out[16] ,
    \cbx_1__1__9_chanx_left_out[17] ,
    \cbx_1__1__9_chanx_left_out[18] ,
    \cbx_1__1__9_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__9_chanx_left_out[0] ,
    \sb_1__1__9_chanx_left_out[1] ,
    \sb_1__1__9_chanx_left_out[2] ,
    \sb_1__1__9_chanx_left_out[3] ,
    \sb_1__1__9_chanx_left_out[4] ,
    \sb_1__1__9_chanx_left_out[5] ,
    \sb_1__1__9_chanx_left_out[6] ,
    \sb_1__1__9_chanx_left_out[7] ,
    \sb_1__1__9_chanx_left_out[8] ,
    \sb_1__1__9_chanx_left_out[9] ,
    \sb_1__1__9_chanx_left_out[10] ,
    \sb_1__1__9_chanx_left_out[11] ,
    \sb_1__1__9_chanx_left_out[12] ,
    \sb_1__1__9_chanx_left_out[13] ,
    \sb_1__1__9_chanx_left_out[14] ,
    \sb_1__1__9_chanx_left_out[15] ,
    \sb_1__1__9_chanx_left_out[16] ,
    \sb_1__1__9_chanx_left_out[17] ,
    \sb_1__1__9_chanx_left_out[18] ,
    \sb_1__1__9_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__9_chanx_right_out[0] ,
    \cbx_1__1__9_chanx_right_out[1] ,
    \cbx_1__1__9_chanx_right_out[2] ,
    \cbx_1__1__9_chanx_right_out[3] ,
    \cbx_1__1__9_chanx_right_out[4] ,
    \cbx_1__1__9_chanx_right_out[5] ,
    \cbx_1__1__9_chanx_right_out[6] ,
    \cbx_1__1__9_chanx_right_out[7] ,
    \cbx_1__1__9_chanx_right_out[8] ,
    \cbx_1__1__9_chanx_right_out[9] ,
    \cbx_1__1__9_chanx_right_out[10] ,
    \cbx_1__1__9_chanx_right_out[11] ,
    \cbx_1__1__9_chanx_right_out[12] ,
    \cbx_1__1__9_chanx_right_out[13] ,
    \cbx_1__1__9_chanx_right_out[14] ,
    \cbx_1__1__9_chanx_right_out[15] ,
    \cbx_1__1__9_chanx_right_out[16] ,
    \cbx_1__1__9_chanx_right_out[17] ,
    \cbx_1__1__9_chanx_right_out[18] ,
    \cbx_1__1__9_chanx_right_out[19] }));
 cbx_1__1_ cbx_2__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[10] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[10] ),
    .SC_IN_BOT(\scff_Wires[27] ),
    .SC_OUT_TOP(\scff_Wires[28] ),
    .bottom_grid_pin_0_(cbx_1__1__10_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__10_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__10_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__10_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__10_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__10_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__10_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__10_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__10_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__10_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__10_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__10_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__10_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__10_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__10_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__10_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__10_ccff_tail),
    .ccff_tail(cbx_1__1__10_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[55] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__3_chanx_right_out[0] ,
    \sb_1__1__3_chanx_right_out[1] ,
    \sb_1__1__3_chanx_right_out[2] ,
    \sb_1__1__3_chanx_right_out[3] ,
    \sb_1__1__3_chanx_right_out[4] ,
    \sb_1__1__3_chanx_right_out[5] ,
    \sb_1__1__3_chanx_right_out[6] ,
    \sb_1__1__3_chanx_right_out[7] ,
    \sb_1__1__3_chanx_right_out[8] ,
    \sb_1__1__3_chanx_right_out[9] ,
    \sb_1__1__3_chanx_right_out[10] ,
    \sb_1__1__3_chanx_right_out[11] ,
    \sb_1__1__3_chanx_right_out[12] ,
    \sb_1__1__3_chanx_right_out[13] ,
    \sb_1__1__3_chanx_right_out[14] ,
    \sb_1__1__3_chanx_right_out[15] ,
    \sb_1__1__3_chanx_right_out[16] ,
    \sb_1__1__3_chanx_right_out[17] ,
    \sb_1__1__3_chanx_right_out[18] ,
    \sb_1__1__3_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__10_chanx_left_out[0] ,
    \cbx_1__1__10_chanx_left_out[1] ,
    \cbx_1__1__10_chanx_left_out[2] ,
    \cbx_1__1__10_chanx_left_out[3] ,
    \cbx_1__1__10_chanx_left_out[4] ,
    \cbx_1__1__10_chanx_left_out[5] ,
    \cbx_1__1__10_chanx_left_out[6] ,
    \cbx_1__1__10_chanx_left_out[7] ,
    \cbx_1__1__10_chanx_left_out[8] ,
    \cbx_1__1__10_chanx_left_out[9] ,
    \cbx_1__1__10_chanx_left_out[10] ,
    \cbx_1__1__10_chanx_left_out[11] ,
    \cbx_1__1__10_chanx_left_out[12] ,
    \cbx_1__1__10_chanx_left_out[13] ,
    \cbx_1__1__10_chanx_left_out[14] ,
    \cbx_1__1__10_chanx_left_out[15] ,
    \cbx_1__1__10_chanx_left_out[16] ,
    \cbx_1__1__10_chanx_left_out[17] ,
    \cbx_1__1__10_chanx_left_out[18] ,
    \cbx_1__1__10_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__10_chanx_left_out[0] ,
    \sb_1__1__10_chanx_left_out[1] ,
    \sb_1__1__10_chanx_left_out[2] ,
    \sb_1__1__10_chanx_left_out[3] ,
    \sb_1__1__10_chanx_left_out[4] ,
    \sb_1__1__10_chanx_left_out[5] ,
    \sb_1__1__10_chanx_left_out[6] ,
    \sb_1__1__10_chanx_left_out[7] ,
    \sb_1__1__10_chanx_left_out[8] ,
    \sb_1__1__10_chanx_left_out[9] ,
    \sb_1__1__10_chanx_left_out[10] ,
    \sb_1__1__10_chanx_left_out[11] ,
    \sb_1__1__10_chanx_left_out[12] ,
    \sb_1__1__10_chanx_left_out[13] ,
    \sb_1__1__10_chanx_left_out[14] ,
    \sb_1__1__10_chanx_left_out[15] ,
    \sb_1__1__10_chanx_left_out[16] ,
    \sb_1__1__10_chanx_left_out[17] ,
    \sb_1__1__10_chanx_left_out[18] ,
    \sb_1__1__10_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__10_chanx_right_out[0] ,
    \cbx_1__1__10_chanx_right_out[1] ,
    \cbx_1__1__10_chanx_right_out[2] ,
    \cbx_1__1__10_chanx_right_out[3] ,
    \cbx_1__1__10_chanx_right_out[4] ,
    \cbx_1__1__10_chanx_right_out[5] ,
    \cbx_1__1__10_chanx_right_out[6] ,
    \cbx_1__1__10_chanx_right_out[7] ,
    \cbx_1__1__10_chanx_right_out[8] ,
    \cbx_1__1__10_chanx_right_out[9] ,
    \cbx_1__1__10_chanx_right_out[10] ,
    \cbx_1__1__10_chanx_right_out[11] ,
    \cbx_1__1__10_chanx_right_out[12] ,
    \cbx_1__1__10_chanx_right_out[13] ,
    \cbx_1__1__10_chanx_right_out[14] ,
    \cbx_1__1__10_chanx_right_out[15] ,
    \cbx_1__1__10_chanx_right_out[16] ,
    \cbx_1__1__10_chanx_right_out[17] ,
    \cbx_1__1__10_chanx_right_out[18] ,
    \cbx_1__1__10_chanx_right_out[19] }));
 cbx_1__1_ cbx_2__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[11] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[11] ),
    .SC_IN_BOT(\scff_Wires[29] ),
    .SC_OUT_TOP(\scff_Wires[30] ),
    .bottom_grid_pin_0_(cbx_1__1__11_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__11_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__11_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__11_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__11_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__11_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__11_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__11_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__11_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__11_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__11_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__11_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__11_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__11_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__11_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__11_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__11_ccff_tail),
    .ccff_tail(cbx_1__1__11_ccff_tail),
    .clk_1_N_out(\clk_1_wires[19] ),
    .clk_1_S_out(\clk_1_wires[20] ),
    .clk_1_W_in(\clk_1_wires[15] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[58] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[19] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[20] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[15] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__4_chanx_right_out[0] ,
    \sb_1__1__4_chanx_right_out[1] ,
    \sb_1__1__4_chanx_right_out[2] ,
    \sb_1__1__4_chanx_right_out[3] ,
    \sb_1__1__4_chanx_right_out[4] ,
    \sb_1__1__4_chanx_right_out[5] ,
    \sb_1__1__4_chanx_right_out[6] ,
    \sb_1__1__4_chanx_right_out[7] ,
    \sb_1__1__4_chanx_right_out[8] ,
    \sb_1__1__4_chanx_right_out[9] ,
    \sb_1__1__4_chanx_right_out[10] ,
    \sb_1__1__4_chanx_right_out[11] ,
    \sb_1__1__4_chanx_right_out[12] ,
    \sb_1__1__4_chanx_right_out[13] ,
    \sb_1__1__4_chanx_right_out[14] ,
    \sb_1__1__4_chanx_right_out[15] ,
    \sb_1__1__4_chanx_right_out[16] ,
    \sb_1__1__4_chanx_right_out[17] ,
    \sb_1__1__4_chanx_right_out[18] ,
    \sb_1__1__4_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__11_chanx_left_out[0] ,
    \cbx_1__1__11_chanx_left_out[1] ,
    \cbx_1__1__11_chanx_left_out[2] ,
    \cbx_1__1__11_chanx_left_out[3] ,
    \cbx_1__1__11_chanx_left_out[4] ,
    \cbx_1__1__11_chanx_left_out[5] ,
    \cbx_1__1__11_chanx_left_out[6] ,
    \cbx_1__1__11_chanx_left_out[7] ,
    \cbx_1__1__11_chanx_left_out[8] ,
    \cbx_1__1__11_chanx_left_out[9] ,
    \cbx_1__1__11_chanx_left_out[10] ,
    \cbx_1__1__11_chanx_left_out[11] ,
    \cbx_1__1__11_chanx_left_out[12] ,
    \cbx_1__1__11_chanx_left_out[13] ,
    \cbx_1__1__11_chanx_left_out[14] ,
    \cbx_1__1__11_chanx_left_out[15] ,
    \cbx_1__1__11_chanx_left_out[16] ,
    \cbx_1__1__11_chanx_left_out[17] ,
    \cbx_1__1__11_chanx_left_out[18] ,
    \cbx_1__1__11_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__11_chanx_left_out[0] ,
    \sb_1__1__11_chanx_left_out[1] ,
    \sb_1__1__11_chanx_left_out[2] ,
    \sb_1__1__11_chanx_left_out[3] ,
    \sb_1__1__11_chanx_left_out[4] ,
    \sb_1__1__11_chanx_left_out[5] ,
    \sb_1__1__11_chanx_left_out[6] ,
    \sb_1__1__11_chanx_left_out[7] ,
    \sb_1__1__11_chanx_left_out[8] ,
    \sb_1__1__11_chanx_left_out[9] ,
    \sb_1__1__11_chanx_left_out[10] ,
    \sb_1__1__11_chanx_left_out[11] ,
    \sb_1__1__11_chanx_left_out[12] ,
    \sb_1__1__11_chanx_left_out[13] ,
    \sb_1__1__11_chanx_left_out[14] ,
    \sb_1__1__11_chanx_left_out[15] ,
    \sb_1__1__11_chanx_left_out[16] ,
    \sb_1__1__11_chanx_left_out[17] ,
    \sb_1__1__11_chanx_left_out[18] ,
    \sb_1__1__11_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__11_chanx_right_out[0] ,
    \cbx_1__1__11_chanx_right_out[1] ,
    \cbx_1__1__11_chanx_right_out[2] ,
    \cbx_1__1__11_chanx_right_out[3] ,
    \cbx_1__1__11_chanx_right_out[4] ,
    \cbx_1__1__11_chanx_right_out[5] ,
    \cbx_1__1__11_chanx_right_out[6] ,
    \cbx_1__1__11_chanx_right_out[7] ,
    \cbx_1__1__11_chanx_right_out[8] ,
    \cbx_1__1__11_chanx_right_out[9] ,
    \cbx_1__1__11_chanx_right_out[10] ,
    \cbx_1__1__11_chanx_right_out[11] ,
    \cbx_1__1__11_chanx_right_out[12] ,
    \cbx_1__1__11_chanx_right_out[13] ,
    \cbx_1__1__11_chanx_right_out[14] ,
    \cbx_1__1__11_chanx_right_out[15] ,
    \cbx_1__1__11_chanx_right_out[16] ,
    \cbx_1__1__11_chanx_right_out[17] ,
    \cbx_1__1__11_chanx_right_out[18] ,
    \cbx_1__1__11_chanx_right_out[19] }));
 cbx_1__1_ cbx_2__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[12] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[12] ),
    .SC_IN_BOT(\scff_Wires[31] ),
    .SC_OUT_TOP(\scff_Wires[32] ),
    .bottom_grid_pin_0_(cbx_1__1__12_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__12_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__12_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__12_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__12_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__12_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__12_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__12_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__12_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__12_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__12_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__12_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__12_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__12_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__12_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__12_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__12_ccff_tail),
    .ccff_tail(cbx_1__1__12_ccff_tail),
    .clk_2_W_in(\clk_2_wires[16] ),
    .clk_2_W_out(\clk_2_wires[17] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[61] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[16] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[17] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__5_chanx_right_out[0] ,
    \sb_1__1__5_chanx_right_out[1] ,
    \sb_1__1__5_chanx_right_out[2] ,
    \sb_1__1__5_chanx_right_out[3] ,
    \sb_1__1__5_chanx_right_out[4] ,
    \sb_1__1__5_chanx_right_out[5] ,
    \sb_1__1__5_chanx_right_out[6] ,
    \sb_1__1__5_chanx_right_out[7] ,
    \sb_1__1__5_chanx_right_out[8] ,
    \sb_1__1__5_chanx_right_out[9] ,
    \sb_1__1__5_chanx_right_out[10] ,
    \sb_1__1__5_chanx_right_out[11] ,
    \sb_1__1__5_chanx_right_out[12] ,
    \sb_1__1__5_chanx_right_out[13] ,
    \sb_1__1__5_chanx_right_out[14] ,
    \sb_1__1__5_chanx_right_out[15] ,
    \sb_1__1__5_chanx_right_out[16] ,
    \sb_1__1__5_chanx_right_out[17] ,
    \sb_1__1__5_chanx_right_out[18] ,
    \sb_1__1__5_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__12_chanx_left_out[0] ,
    \cbx_1__1__12_chanx_left_out[1] ,
    \cbx_1__1__12_chanx_left_out[2] ,
    \cbx_1__1__12_chanx_left_out[3] ,
    \cbx_1__1__12_chanx_left_out[4] ,
    \cbx_1__1__12_chanx_left_out[5] ,
    \cbx_1__1__12_chanx_left_out[6] ,
    \cbx_1__1__12_chanx_left_out[7] ,
    \cbx_1__1__12_chanx_left_out[8] ,
    \cbx_1__1__12_chanx_left_out[9] ,
    \cbx_1__1__12_chanx_left_out[10] ,
    \cbx_1__1__12_chanx_left_out[11] ,
    \cbx_1__1__12_chanx_left_out[12] ,
    \cbx_1__1__12_chanx_left_out[13] ,
    \cbx_1__1__12_chanx_left_out[14] ,
    \cbx_1__1__12_chanx_left_out[15] ,
    \cbx_1__1__12_chanx_left_out[16] ,
    \cbx_1__1__12_chanx_left_out[17] ,
    \cbx_1__1__12_chanx_left_out[18] ,
    \cbx_1__1__12_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__12_chanx_left_out[0] ,
    \sb_1__1__12_chanx_left_out[1] ,
    \sb_1__1__12_chanx_left_out[2] ,
    \sb_1__1__12_chanx_left_out[3] ,
    \sb_1__1__12_chanx_left_out[4] ,
    \sb_1__1__12_chanx_left_out[5] ,
    \sb_1__1__12_chanx_left_out[6] ,
    \sb_1__1__12_chanx_left_out[7] ,
    \sb_1__1__12_chanx_left_out[8] ,
    \sb_1__1__12_chanx_left_out[9] ,
    \sb_1__1__12_chanx_left_out[10] ,
    \sb_1__1__12_chanx_left_out[11] ,
    \sb_1__1__12_chanx_left_out[12] ,
    \sb_1__1__12_chanx_left_out[13] ,
    \sb_1__1__12_chanx_left_out[14] ,
    \sb_1__1__12_chanx_left_out[15] ,
    \sb_1__1__12_chanx_left_out[16] ,
    \sb_1__1__12_chanx_left_out[17] ,
    \sb_1__1__12_chanx_left_out[18] ,
    \sb_1__1__12_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__12_chanx_right_out[0] ,
    \cbx_1__1__12_chanx_right_out[1] ,
    \cbx_1__1__12_chanx_right_out[2] ,
    \cbx_1__1__12_chanx_right_out[3] ,
    \cbx_1__1__12_chanx_right_out[4] ,
    \cbx_1__1__12_chanx_right_out[5] ,
    \cbx_1__1__12_chanx_right_out[6] ,
    \cbx_1__1__12_chanx_right_out[7] ,
    \cbx_1__1__12_chanx_right_out[8] ,
    \cbx_1__1__12_chanx_right_out[9] ,
    \cbx_1__1__12_chanx_right_out[10] ,
    \cbx_1__1__12_chanx_right_out[11] ,
    \cbx_1__1__12_chanx_right_out[12] ,
    \cbx_1__1__12_chanx_right_out[13] ,
    \cbx_1__1__12_chanx_right_out[14] ,
    \cbx_1__1__12_chanx_right_out[15] ,
    \cbx_1__1__12_chanx_right_out[16] ,
    \cbx_1__1__12_chanx_right_out[17] ,
    \cbx_1__1__12_chanx_right_out[18] ,
    \cbx_1__1__12_chanx_right_out[19] }));
 cbx_1__1_ cbx_2__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[13] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[13] ),
    .SC_IN_BOT(\scff_Wires[33] ),
    .SC_OUT_TOP(\scff_Wires[34] ),
    .bottom_grid_pin_0_(cbx_1__1__13_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__13_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__13_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__13_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__13_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__13_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__13_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__13_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__13_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__13_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__13_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__13_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__13_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__13_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__13_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__13_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__13_ccff_tail),
    .ccff_tail(cbx_1__1__13_ccff_tail),
    .clk_1_N_out(\clk_1_wires[26] ),
    .clk_1_S_out(\clk_1_wires[27] ),
    .clk_1_W_in(\clk_1_wires[22] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[64] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[26] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[27] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[22] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__6_chanx_right_out[0] ,
    \sb_1__1__6_chanx_right_out[1] ,
    \sb_1__1__6_chanx_right_out[2] ,
    \sb_1__1__6_chanx_right_out[3] ,
    \sb_1__1__6_chanx_right_out[4] ,
    \sb_1__1__6_chanx_right_out[5] ,
    \sb_1__1__6_chanx_right_out[6] ,
    \sb_1__1__6_chanx_right_out[7] ,
    \sb_1__1__6_chanx_right_out[8] ,
    \sb_1__1__6_chanx_right_out[9] ,
    \sb_1__1__6_chanx_right_out[10] ,
    \sb_1__1__6_chanx_right_out[11] ,
    \sb_1__1__6_chanx_right_out[12] ,
    \sb_1__1__6_chanx_right_out[13] ,
    \sb_1__1__6_chanx_right_out[14] ,
    \sb_1__1__6_chanx_right_out[15] ,
    \sb_1__1__6_chanx_right_out[16] ,
    \sb_1__1__6_chanx_right_out[17] ,
    \sb_1__1__6_chanx_right_out[18] ,
    \sb_1__1__6_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__13_chanx_left_out[0] ,
    \cbx_1__1__13_chanx_left_out[1] ,
    \cbx_1__1__13_chanx_left_out[2] ,
    \cbx_1__1__13_chanx_left_out[3] ,
    \cbx_1__1__13_chanx_left_out[4] ,
    \cbx_1__1__13_chanx_left_out[5] ,
    \cbx_1__1__13_chanx_left_out[6] ,
    \cbx_1__1__13_chanx_left_out[7] ,
    \cbx_1__1__13_chanx_left_out[8] ,
    \cbx_1__1__13_chanx_left_out[9] ,
    \cbx_1__1__13_chanx_left_out[10] ,
    \cbx_1__1__13_chanx_left_out[11] ,
    \cbx_1__1__13_chanx_left_out[12] ,
    \cbx_1__1__13_chanx_left_out[13] ,
    \cbx_1__1__13_chanx_left_out[14] ,
    \cbx_1__1__13_chanx_left_out[15] ,
    \cbx_1__1__13_chanx_left_out[16] ,
    \cbx_1__1__13_chanx_left_out[17] ,
    \cbx_1__1__13_chanx_left_out[18] ,
    \cbx_1__1__13_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__13_chanx_left_out[0] ,
    \sb_1__1__13_chanx_left_out[1] ,
    \sb_1__1__13_chanx_left_out[2] ,
    \sb_1__1__13_chanx_left_out[3] ,
    \sb_1__1__13_chanx_left_out[4] ,
    \sb_1__1__13_chanx_left_out[5] ,
    \sb_1__1__13_chanx_left_out[6] ,
    \sb_1__1__13_chanx_left_out[7] ,
    \sb_1__1__13_chanx_left_out[8] ,
    \sb_1__1__13_chanx_left_out[9] ,
    \sb_1__1__13_chanx_left_out[10] ,
    \sb_1__1__13_chanx_left_out[11] ,
    \sb_1__1__13_chanx_left_out[12] ,
    \sb_1__1__13_chanx_left_out[13] ,
    \sb_1__1__13_chanx_left_out[14] ,
    \sb_1__1__13_chanx_left_out[15] ,
    \sb_1__1__13_chanx_left_out[16] ,
    \sb_1__1__13_chanx_left_out[17] ,
    \sb_1__1__13_chanx_left_out[18] ,
    \sb_1__1__13_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__13_chanx_right_out[0] ,
    \cbx_1__1__13_chanx_right_out[1] ,
    \cbx_1__1__13_chanx_right_out[2] ,
    \cbx_1__1__13_chanx_right_out[3] ,
    \cbx_1__1__13_chanx_right_out[4] ,
    \cbx_1__1__13_chanx_right_out[5] ,
    \cbx_1__1__13_chanx_right_out[6] ,
    \cbx_1__1__13_chanx_right_out[7] ,
    \cbx_1__1__13_chanx_right_out[8] ,
    \cbx_1__1__13_chanx_right_out[9] ,
    \cbx_1__1__13_chanx_right_out[10] ,
    \cbx_1__1__13_chanx_right_out[11] ,
    \cbx_1__1__13_chanx_right_out[12] ,
    \cbx_1__1__13_chanx_right_out[13] ,
    \cbx_1__1__13_chanx_right_out[14] ,
    \cbx_1__1__13_chanx_right_out[15] ,
    \cbx_1__1__13_chanx_right_out[16] ,
    \cbx_1__1__13_chanx_right_out[17] ,
    \cbx_1__1__13_chanx_right_out[18] ,
    \cbx_1__1__13_chanx_right_out[19] }));
 cbx_1__2_ cbx_2__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[35] ),
    .SC_OUT_TOP(\scff_Wires[36] ),
    .bottom_grid_pin_0_(cbx_1__8__1_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__1_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__1_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__1_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__1_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__1_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__1_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__1_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__1_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__1_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__1_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__1_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__1_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__1_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__1_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__1_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__1_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_1_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_1_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_1__8__1_ccff_tail),
    .ccff_tail(grid_io_top_1_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]),
    .prog_clk_0_S_in(\prog_clk_0_wires[67] ),
    .top_grid_pin_0_(cbx_1__8__1_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__8__0_chanx_right_out[0] ,
    \sb_1__8__0_chanx_right_out[1] ,
    \sb_1__8__0_chanx_right_out[2] ,
    \sb_1__8__0_chanx_right_out[3] ,
    \sb_1__8__0_chanx_right_out[4] ,
    \sb_1__8__0_chanx_right_out[5] ,
    \sb_1__8__0_chanx_right_out[6] ,
    \sb_1__8__0_chanx_right_out[7] ,
    \sb_1__8__0_chanx_right_out[8] ,
    \sb_1__8__0_chanx_right_out[9] ,
    \sb_1__8__0_chanx_right_out[10] ,
    \sb_1__8__0_chanx_right_out[11] ,
    \sb_1__8__0_chanx_right_out[12] ,
    \sb_1__8__0_chanx_right_out[13] ,
    \sb_1__8__0_chanx_right_out[14] ,
    \sb_1__8__0_chanx_right_out[15] ,
    \sb_1__8__0_chanx_right_out[16] ,
    \sb_1__8__0_chanx_right_out[17] ,
    \sb_1__8__0_chanx_right_out[18] ,
    \sb_1__8__0_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__1_chanx_left_out[0] ,
    \cbx_1__8__1_chanx_left_out[1] ,
    \cbx_1__8__1_chanx_left_out[2] ,
    \cbx_1__8__1_chanx_left_out[3] ,
    \cbx_1__8__1_chanx_left_out[4] ,
    \cbx_1__8__1_chanx_left_out[5] ,
    \cbx_1__8__1_chanx_left_out[6] ,
    \cbx_1__8__1_chanx_left_out[7] ,
    \cbx_1__8__1_chanx_left_out[8] ,
    \cbx_1__8__1_chanx_left_out[9] ,
    \cbx_1__8__1_chanx_left_out[10] ,
    \cbx_1__8__1_chanx_left_out[11] ,
    \cbx_1__8__1_chanx_left_out[12] ,
    \cbx_1__8__1_chanx_left_out[13] ,
    \cbx_1__8__1_chanx_left_out[14] ,
    \cbx_1__8__1_chanx_left_out[15] ,
    \cbx_1__8__1_chanx_left_out[16] ,
    \cbx_1__8__1_chanx_left_out[17] ,
    \cbx_1__8__1_chanx_left_out[18] ,
    \cbx_1__8__1_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__8__1_chanx_left_out[0] ,
    \sb_1__8__1_chanx_left_out[1] ,
    \sb_1__8__1_chanx_left_out[2] ,
    \sb_1__8__1_chanx_left_out[3] ,
    \sb_1__8__1_chanx_left_out[4] ,
    \sb_1__8__1_chanx_left_out[5] ,
    \sb_1__8__1_chanx_left_out[6] ,
    \sb_1__8__1_chanx_left_out[7] ,
    \sb_1__8__1_chanx_left_out[8] ,
    \sb_1__8__1_chanx_left_out[9] ,
    \sb_1__8__1_chanx_left_out[10] ,
    \sb_1__8__1_chanx_left_out[11] ,
    \sb_1__8__1_chanx_left_out[12] ,
    \sb_1__8__1_chanx_left_out[13] ,
    \sb_1__8__1_chanx_left_out[14] ,
    \sb_1__8__1_chanx_left_out[15] ,
    \sb_1__8__1_chanx_left_out[16] ,
    \sb_1__8__1_chanx_left_out[17] ,
    \sb_1__8__1_chanx_left_out[18] ,
    \sb_1__8__1_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__1_chanx_right_out[0] ,
    \cbx_1__8__1_chanx_right_out[1] ,
    \cbx_1__8__1_chanx_right_out[2] ,
    \cbx_1__8__1_chanx_right_out[3] ,
    \cbx_1__8__1_chanx_right_out[4] ,
    \cbx_1__8__1_chanx_right_out[5] ,
    \cbx_1__8__1_chanx_right_out[6] ,
    \cbx_1__8__1_chanx_right_out[7] ,
    \cbx_1__8__1_chanx_right_out[8] ,
    \cbx_1__8__1_chanx_right_out[9] ,
    \cbx_1__8__1_chanx_right_out[10] ,
    \cbx_1__8__1_chanx_right_out[11] ,
    \cbx_1__8__1_chanx_right_out[12] ,
    \cbx_1__8__1_chanx_right_out[13] ,
    \cbx_1__8__1_chanx_right_out[14] ,
    \cbx_1__8__1_chanx_right_out[15] ,
    \cbx_1__8__1_chanx_right_out[16] ,
    \cbx_1__8__1_chanx_right_out[17] ,
    \cbx_1__8__1_chanx_right_out[18] ,
    \cbx_1__8__1_chanx_right_out[19] }));
 cbx_1__0_ cbx_3__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[54] ),
    .SC_OUT_BOT(\scff_Wires[55] ),
    .bottom_grid_pin_0_(cbx_1__0__2_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__2_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__2_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__2_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__2_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__2_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__2_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__2_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__2_bottom_grid_pin_8_),
    .ccff_head(sb_1__0__2_ccff_tail),
    .ccff_tail(grid_io_bottom_5_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[69] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__2_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__2_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_5_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_5_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__2_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_5_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_5_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__2_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_5_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_5_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__2_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_5_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_5_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_5_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_5_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__2_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_5_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_5_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__2_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_5_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_5_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__2_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_5_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_5_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__2_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_5_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_5_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__0__1_chanx_right_out[0] ,
    \sb_1__0__1_chanx_right_out[1] ,
    \sb_1__0__1_chanx_right_out[2] ,
    \sb_1__0__1_chanx_right_out[3] ,
    \sb_1__0__1_chanx_right_out[4] ,
    \sb_1__0__1_chanx_right_out[5] ,
    \sb_1__0__1_chanx_right_out[6] ,
    \sb_1__0__1_chanx_right_out[7] ,
    \sb_1__0__1_chanx_right_out[8] ,
    \sb_1__0__1_chanx_right_out[9] ,
    \sb_1__0__1_chanx_right_out[10] ,
    \sb_1__0__1_chanx_right_out[11] ,
    \sb_1__0__1_chanx_right_out[12] ,
    \sb_1__0__1_chanx_right_out[13] ,
    \sb_1__0__1_chanx_right_out[14] ,
    \sb_1__0__1_chanx_right_out[15] ,
    \sb_1__0__1_chanx_right_out[16] ,
    \sb_1__0__1_chanx_right_out[17] ,
    \sb_1__0__1_chanx_right_out[18] ,
    \sb_1__0__1_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__2_chanx_left_out[0] ,
    \cbx_1__0__2_chanx_left_out[1] ,
    \cbx_1__0__2_chanx_left_out[2] ,
    \cbx_1__0__2_chanx_left_out[3] ,
    \cbx_1__0__2_chanx_left_out[4] ,
    \cbx_1__0__2_chanx_left_out[5] ,
    \cbx_1__0__2_chanx_left_out[6] ,
    \cbx_1__0__2_chanx_left_out[7] ,
    \cbx_1__0__2_chanx_left_out[8] ,
    \cbx_1__0__2_chanx_left_out[9] ,
    \cbx_1__0__2_chanx_left_out[10] ,
    \cbx_1__0__2_chanx_left_out[11] ,
    \cbx_1__0__2_chanx_left_out[12] ,
    \cbx_1__0__2_chanx_left_out[13] ,
    \cbx_1__0__2_chanx_left_out[14] ,
    \cbx_1__0__2_chanx_left_out[15] ,
    \cbx_1__0__2_chanx_left_out[16] ,
    \cbx_1__0__2_chanx_left_out[17] ,
    \cbx_1__0__2_chanx_left_out[18] ,
    \cbx_1__0__2_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__0__2_chanx_left_out[0] ,
    \sb_1__0__2_chanx_left_out[1] ,
    \sb_1__0__2_chanx_left_out[2] ,
    \sb_1__0__2_chanx_left_out[3] ,
    \sb_1__0__2_chanx_left_out[4] ,
    \sb_1__0__2_chanx_left_out[5] ,
    \sb_1__0__2_chanx_left_out[6] ,
    \sb_1__0__2_chanx_left_out[7] ,
    \sb_1__0__2_chanx_left_out[8] ,
    \sb_1__0__2_chanx_left_out[9] ,
    \sb_1__0__2_chanx_left_out[10] ,
    \sb_1__0__2_chanx_left_out[11] ,
    \sb_1__0__2_chanx_left_out[12] ,
    \sb_1__0__2_chanx_left_out[13] ,
    \sb_1__0__2_chanx_left_out[14] ,
    \sb_1__0__2_chanx_left_out[15] ,
    \sb_1__0__2_chanx_left_out[16] ,
    \sb_1__0__2_chanx_left_out[17] ,
    \sb_1__0__2_chanx_left_out[18] ,
    \sb_1__0__2_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__2_chanx_right_out[0] ,
    \cbx_1__0__2_chanx_right_out[1] ,
    \cbx_1__0__2_chanx_right_out[2] ,
    \cbx_1__0__2_chanx_right_out[3] ,
    \cbx_1__0__2_chanx_right_out[4] ,
    \cbx_1__0__2_chanx_right_out[5] ,
    \cbx_1__0__2_chanx_right_out[6] ,
    \cbx_1__0__2_chanx_right_out[7] ,
    \cbx_1__0__2_chanx_right_out[8] ,
    \cbx_1__0__2_chanx_right_out[9] ,
    \cbx_1__0__2_chanx_right_out[10] ,
    \cbx_1__0__2_chanx_right_out[11] ,
    \cbx_1__0__2_chanx_right_out[12] ,
    \cbx_1__0__2_chanx_right_out[13] ,
    \cbx_1__0__2_chanx_right_out[14] ,
    \cbx_1__0__2_chanx_right_out[15] ,
    \cbx_1__0__2_chanx_right_out[16] ,
    \cbx_1__0__2_chanx_right_out[17] ,
    \cbx_1__0__2_chanx_right_out[18] ,
    \cbx_1__0__2_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]}));
 cbx_1__1_ cbx_3__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[14] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[14] ),
    .SC_IN_TOP(\scff_Wires[51] ),
    .SC_OUT_BOT(\scff_Wires[52] ),
    .bottom_grid_pin_0_(cbx_1__1__14_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__14_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__14_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__14_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__14_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__14_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__14_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__14_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__14_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__14_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__14_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__14_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__14_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__14_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__14_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__14_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__14_ccff_tail),
    .ccff_tail(cbx_1__1__14_ccff_tail),
    .clk_1_N_out(\clk_1_wires[31] ),
    .clk_1_S_out(\clk_1_wires[32] ),
    .clk_1_W_in(\clk_1_wires[30] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[72] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[31] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[32] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[30] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__7_chanx_right_out[0] ,
    \sb_1__1__7_chanx_right_out[1] ,
    \sb_1__1__7_chanx_right_out[2] ,
    \sb_1__1__7_chanx_right_out[3] ,
    \sb_1__1__7_chanx_right_out[4] ,
    \sb_1__1__7_chanx_right_out[5] ,
    \sb_1__1__7_chanx_right_out[6] ,
    \sb_1__1__7_chanx_right_out[7] ,
    \sb_1__1__7_chanx_right_out[8] ,
    \sb_1__1__7_chanx_right_out[9] ,
    \sb_1__1__7_chanx_right_out[10] ,
    \sb_1__1__7_chanx_right_out[11] ,
    \sb_1__1__7_chanx_right_out[12] ,
    \sb_1__1__7_chanx_right_out[13] ,
    \sb_1__1__7_chanx_right_out[14] ,
    \sb_1__1__7_chanx_right_out[15] ,
    \sb_1__1__7_chanx_right_out[16] ,
    \sb_1__1__7_chanx_right_out[17] ,
    \sb_1__1__7_chanx_right_out[18] ,
    \sb_1__1__7_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__14_chanx_left_out[0] ,
    \cbx_1__1__14_chanx_left_out[1] ,
    \cbx_1__1__14_chanx_left_out[2] ,
    \cbx_1__1__14_chanx_left_out[3] ,
    \cbx_1__1__14_chanx_left_out[4] ,
    \cbx_1__1__14_chanx_left_out[5] ,
    \cbx_1__1__14_chanx_left_out[6] ,
    \cbx_1__1__14_chanx_left_out[7] ,
    \cbx_1__1__14_chanx_left_out[8] ,
    \cbx_1__1__14_chanx_left_out[9] ,
    \cbx_1__1__14_chanx_left_out[10] ,
    \cbx_1__1__14_chanx_left_out[11] ,
    \cbx_1__1__14_chanx_left_out[12] ,
    \cbx_1__1__14_chanx_left_out[13] ,
    \cbx_1__1__14_chanx_left_out[14] ,
    \cbx_1__1__14_chanx_left_out[15] ,
    \cbx_1__1__14_chanx_left_out[16] ,
    \cbx_1__1__14_chanx_left_out[17] ,
    \cbx_1__1__14_chanx_left_out[18] ,
    \cbx_1__1__14_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__14_chanx_left_out[0] ,
    \sb_1__1__14_chanx_left_out[1] ,
    \sb_1__1__14_chanx_left_out[2] ,
    \sb_1__1__14_chanx_left_out[3] ,
    \sb_1__1__14_chanx_left_out[4] ,
    \sb_1__1__14_chanx_left_out[5] ,
    \sb_1__1__14_chanx_left_out[6] ,
    \sb_1__1__14_chanx_left_out[7] ,
    \sb_1__1__14_chanx_left_out[8] ,
    \sb_1__1__14_chanx_left_out[9] ,
    \sb_1__1__14_chanx_left_out[10] ,
    \sb_1__1__14_chanx_left_out[11] ,
    \sb_1__1__14_chanx_left_out[12] ,
    \sb_1__1__14_chanx_left_out[13] ,
    \sb_1__1__14_chanx_left_out[14] ,
    \sb_1__1__14_chanx_left_out[15] ,
    \sb_1__1__14_chanx_left_out[16] ,
    \sb_1__1__14_chanx_left_out[17] ,
    \sb_1__1__14_chanx_left_out[18] ,
    \sb_1__1__14_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__14_chanx_right_out[0] ,
    \cbx_1__1__14_chanx_right_out[1] ,
    \cbx_1__1__14_chanx_right_out[2] ,
    \cbx_1__1__14_chanx_right_out[3] ,
    \cbx_1__1__14_chanx_right_out[4] ,
    \cbx_1__1__14_chanx_right_out[5] ,
    \cbx_1__1__14_chanx_right_out[6] ,
    \cbx_1__1__14_chanx_right_out[7] ,
    \cbx_1__1__14_chanx_right_out[8] ,
    \cbx_1__1__14_chanx_right_out[9] ,
    \cbx_1__1__14_chanx_right_out[10] ,
    \cbx_1__1__14_chanx_right_out[11] ,
    \cbx_1__1__14_chanx_right_out[12] ,
    \cbx_1__1__14_chanx_right_out[13] ,
    \cbx_1__1__14_chanx_right_out[14] ,
    \cbx_1__1__14_chanx_right_out[15] ,
    \cbx_1__1__14_chanx_right_out[16] ,
    \cbx_1__1__14_chanx_right_out[17] ,
    \cbx_1__1__14_chanx_right_out[18] ,
    \cbx_1__1__14_chanx_right_out[19] }));
 cbx_1__1_ cbx_3__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[15] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[15] ),
    .SC_IN_TOP(\scff_Wires[49] ),
    .SC_OUT_BOT(\scff_Wires[50] ),
    .bottom_grid_pin_0_(cbx_1__1__15_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__15_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__15_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__15_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__15_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__15_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__15_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__15_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__15_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__15_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__15_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__15_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__15_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__15_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__15_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__15_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__15_ccff_tail),
    .ccff_tail(cbx_1__1__15_ccff_tail),
    .clk_2_E_out(\clk_2_wires[2] ),
    .clk_2_W_in(\clk_2_wires[1] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[75] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[2] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[1] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__8_chanx_right_out[0] ,
    \sb_1__1__8_chanx_right_out[1] ,
    \sb_1__1__8_chanx_right_out[2] ,
    \sb_1__1__8_chanx_right_out[3] ,
    \sb_1__1__8_chanx_right_out[4] ,
    \sb_1__1__8_chanx_right_out[5] ,
    \sb_1__1__8_chanx_right_out[6] ,
    \sb_1__1__8_chanx_right_out[7] ,
    \sb_1__1__8_chanx_right_out[8] ,
    \sb_1__1__8_chanx_right_out[9] ,
    \sb_1__1__8_chanx_right_out[10] ,
    \sb_1__1__8_chanx_right_out[11] ,
    \sb_1__1__8_chanx_right_out[12] ,
    \sb_1__1__8_chanx_right_out[13] ,
    \sb_1__1__8_chanx_right_out[14] ,
    \sb_1__1__8_chanx_right_out[15] ,
    \sb_1__1__8_chanx_right_out[16] ,
    \sb_1__1__8_chanx_right_out[17] ,
    \sb_1__1__8_chanx_right_out[18] ,
    \sb_1__1__8_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__15_chanx_left_out[0] ,
    \cbx_1__1__15_chanx_left_out[1] ,
    \cbx_1__1__15_chanx_left_out[2] ,
    \cbx_1__1__15_chanx_left_out[3] ,
    \cbx_1__1__15_chanx_left_out[4] ,
    \cbx_1__1__15_chanx_left_out[5] ,
    \cbx_1__1__15_chanx_left_out[6] ,
    \cbx_1__1__15_chanx_left_out[7] ,
    \cbx_1__1__15_chanx_left_out[8] ,
    \cbx_1__1__15_chanx_left_out[9] ,
    \cbx_1__1__15_chanx_left_out[10] ,
    \cbx_1__1__15_chanx_left_out[11] ,
    \cbx_1__1__15_chanx_left_out[12] ,
    \cbx_1__1__15_chanx_left_out[13] ,
    \cbx_1__1__15_chanx_left_out[14] ,
    \cbx_1__1__15_chanx_left_out[15] ,
    \cbx_1__1__15_chanx_left_out[16] ,
    \cbx_1__1__15_chanx_left_out[17] ,
    \cbx_1__1__15_chanx_left_out[18] ,
    \cbx_1__1__15_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__15_chanx_left_out[0] ,
    \sb_1__1__15_chanx_left_out[1] ,
    \sb_1__1__15_chanx_left_out[2] ,
    \sb_1__1__15_chanx_left_out[3] ,
    \sb_1__1__15_chanx_left_out[4] ,
    \sb_1__1__15_chanx_left_out[5] ,
    \sb_1__1__15_chanx_left_out[6] ,
    \sb_1__1__15_chanx_left_out[7] ,
    \sb_1__1__15_chanx_left_out[8] ,
    \sb_1__1__15_chanx_left_out[9] ,
    \sb_1__1__15_chanx_left_out[10] ,
    \sb_1__1__15_chanx_left_out[11] ,
    \sb_1__1__15_chanx_left_out[12] ,
    \sb_1__1__15_chanx_left_out[13] ,
    \sb_1__1__15_chanx_left_out[14] ,
    \sb_1__1__15_chanx_left_out[15] ,
    \sb_1__1__15_chanx_left_out[16] ,
    \sb_1__1__15_chanx_left_out[17] ,
    \sb_1__1__15_chanx_left_out[18] ,
    \sb_1__1__15_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__15_chanx_right_out[0] ,
    \cbx_1__1__15_chanx_right_out[1] ,
    \cbx_1__1__15_chanx_right_out[2] ,
    \cbx_1__1__15_chanx_right_out[3] ,
    \cbx_1__1__15_chanx_right_out[4] ,
    \cbx_1__1__15_chanx_right_out[5] ,
    \cbx_1__1__15_chanx_right_out[6] ,
    \cbx_1__1__15_chanx_right_out[7] ,
    \cbx_1__1__15_chanx_right_out[8] ,
    \cbx_1__1__15_chanx_right_out[9] ,
    \cbx_1__1__15_chanx_right_out[10] ,
    \cbx_1__1__15_chanx_right_out[11] ,
    \cbx_1__1__15_chanx_right_out[12] ,
    \cbx_1__1__15_chanx_right_out[13] ,
    \cbx_1__1__15_chanx_right_out[14] ,
    \cbx_1__1__15_chanx_right_out[15] ,
    \cbx_1__1__15_chanx_right_out[16] ,
    \cbx_1__1__15_chanx_right_out[17] ,
    \cbx_1__1__15_chanx_right_out[18] ,
    \cbx_1__1__15_chanx_right_out[19] }));
 cbx_1__1_ cbx_3__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[16] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[16] ),
    .SC_IN_TOP(\scff_Wires[47] ),
    .SC_OUT_BOT(\scff_Wires[48] ),
    .bottom_grid_pin_0_(cbx_1__1__16_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__16_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__16_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__16_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__16_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__16_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__16_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__16_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__16_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__16_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__16_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__16_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__16_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__16_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__16_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__16_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__16_ccff_tail),
    .ccff_tail(cbx_1__1__16_ccff_tail),
    .clk_1_N_out(\clk_1_wires[38] ),
    .clk_1_S_out(\clk_1_wires[39] ),
    .clk_1_W_in(\clk_1_wires[37] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[78] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[38] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[39] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[37] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__9_chanx_right_out[0] ,
    \sb_1__1__9_chanx_right_out[1] ,
    \sb_1__1__9_chanx_right_out[2] ,
    \sb_1__1__9_chanx_right_out[3] ,
    \sb_1__1__9_chanx_right_out[4] ,
    \sb_1__1__9_chanx_right_out[5] ,
    \sb_1__1__9_chanx_right_out[6] ,
    \sb_1__1__9_chanx_right_out[7] ,
    \sb_1__1__9_chanx_right_out[8] ,
    \sb_1__1__9_chanx_right_out[9] ,
    \sb_1__1__9_chanx_right_out[10] ,
    \sb_1__1__9_chanx_right_out[11] ,
    \sb_1__1__9_chanx_right_out[12] ,
    \sb_1__1__9_chanx_right_out[13] ,
    \sb_1__1__9_chanx_right_out[14] ,
    \sb_1__1__9_chanx_right_out[15] ,
    \sb_1__1__9_chanx_right_out[16] ,
    \sb_1__1__9_chanx_right_out[17] ,
    \sb_1__1__9_chanx_right_out[18] ,
    \sb_1__1__9_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__16_chanx_left_out[0] ,
    \cbx_1__1__16_chanx_left_out[1] ,
    \cbx_1__1__16_chanx_left_out[2] ,
    \cbx_1__1__16_chanx_left_out[3] ,
    \cbx_1__1__16_chanx_left_out[4] ,
    \cbx_1__1__16_chanx_left_out[5] ,
    \cbx_1__1__16_chanx_left_out[6] ,
    \cbx_1__1__16_chanx_left_out[7] ,
    \cbx_1__1__16_chanx_left_out[8] ,
    \cbx_1__1__16_chanx_left_out[9] ,
    \cbx_1__1__16_chanx_left_out[10] ,
    \cbx_1__1__16_chanx_left_out[11] ,
    \cbx_1__1__16_chanx_left_out[12] ,
    \cbx_1__1__16_chanx_left_out[13] ,
    \cbx_1__1__16_chanx_left_out[14] ,
    \cbx_1__1__16_chanx_left_out[15] ,
    \cbx_1__1__16_chanx_left_out[16] ,
    \cbx_1__1__16_chanx_left_out[17] ,
    \cbx_1__1__16_chanx_left_out[18] ,
    \cbx_1__1__16_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__16_chanx_left_out[0] ,
    \sb_1__1__16_chanx_left_out[1] ,
    \sb_1__1__16_chanx_left_out[2] ,
    \sb_1__1__16_chanx_left_out[3] ,
    \sb_1__1__16_chanx_left_out[4] ,
    \sb_1__1__16_chanx_left_out[5] ,
    \sb_1__1__16_chanx_left_out[6] ,
    \sb_1__1__16_chanx_left_out[7] ,
    \sb_1__1__16_chanx_left_out[8] ,
    \sb_1__1__16_chanx_left_out[9] ,
    \sb_1__1__16_chanx_left_out[10] ,
    \sb_1__1__16_chanx_left_out[11] ,
    \sb_1__1__16_chanx_left_out[12] ,
    \sb_1__1__16_chanx_left_out[13] ,
    \sb_1__1__16_chanx_left_out[14] ,
    \sb_1__1__16_chanx_left_out[15] ,
    \sb_1__1__16_chanx_left_out[16] ,
    \sb_1__1__16_chanx_left_out[17] ,
    \sb_1__1__16_chanx_left_out[18] ,
    \sb_1__1__16_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__16_chanx_right_out[0] ,
    \cbx_1__1__16_chanx_right_out[1] ,
    \cbx_1__1__16_chanx_right_out[2] ,
    \cbx_1__1__16_chanx_right_out[3] ,
    \cbx_1__1__16_chanx_right_out[4] ,
    \cbx_1__1__16_chanx_right_out[5] ,
    \cbx_1__1__16_chanx_right_out[6] ,
    \cbx_1__1__16_chanx_right_out[7] ,
    \cbx_1__1__16_chanx_right_out[8] ,
    \cbx_1__1__16_chanx_right_out[9] ,
    \cbx_1__1__16_chanx_right_out[10] ,
    \cbx_1__1__16_chanx_right_out[11] ,
    \cbx_1__1__16_chanx_right_out[12] ,
    \cbx_1__1__16_chanx_right_out[13] ,
    \cbx_1__1__16_chanx_right_out[14] ,
    \cbx_1__1__16_chanx_right_out[15] ,
    \cbx_1__1__16_chanx_right_out[16] ,
    \cbx_1__1__16_chanx_right_out[17] ,
    \cbx_1__1__16_chanx_right_out[18] ,
    \cbx_1__1__16_chanx_right_out[19] }));
 cbx_1__1_ cbx_3__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[17] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[17] ),
    .SC_IN_TOP(\scff_Wires[45] ),
    .SC_OUT_BOT(\scff_Wires[46] ),
    .bottom_grid_pin_0_(cbx_1__1__17_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__17_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__17_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__17_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__17_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__17_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__17_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__17_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__17_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__17_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__17_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__17_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__17_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__17_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__17_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__17_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__17_ccff_tail),
    .ccff_tail(cbx_1__1__17_ccff_tail),
    .clk_3_W_in(\clk_3_wires[8] ),
    .clk_3_W_out(\clk_3_wires[9] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[81] ),
    .prog_clk_3_W_in(\prog_clk_3_wires[8] ),
    .prog_clk_3_W_out(\prog_clk_3_wires[9] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__10_chanx_right_out[0] ,
    \sb_1__1__10_chanx_right_out[1] ,
    \sb_1__1__10_chanx_right_out[2] ,
    \sb_1__1__10_chanx_right_out[3] ,
    \sb_1__1__10_chanx_right_out[4] ,
    \sb_1__1__10_chanx_right_out[5] ,
    \sb_1__1__10_chanx_right_out[6] ,
    \sb_1__1__10_chanx_right_out[7] ,
    \sb_1__1__10_chanx_right_out[8] ,
    \sb_1__1__10_chanx_right_out[9] ,
    \sb_1__1__10_chanx_right_out[10] ,
    \sb_1__1__10_chanx_right_out[11] ,
    \sb_1__1__10_chanx_right_out[12] ,
    \sb_1__1__10_chanx_right_out[13] ,
    \sb_1__1__10_chanx_right_out[14] ,
    \sb_1__1__10_chanx_right_out[15] ,
    \sb_1__1__10_chanx_right_out[16] ,
    \sb_1__1__10_chanx_right_out[17] ,
    \sb_1__1__10_chanx_right_out[18] ,
    \sb_1__1__10_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__17_chanx_left_out[0] ,
    \cbx_1__1__17_chanx_left_out[1] ,
    \cbx_1__1__17_chanx_left_out[2] ,
    \cbx_1__1__17_chanx_left_out[3] ,
    \cbx_1__1__17_chanx_left_out[4] ,
    \cbx_1__1__17_chanx_left_out[5] ,
    \cbx_1__1__17_chanx_left_out[6] ,
    \cbx_1__1__17_chanx_left_out[7] ,
    \cbx_1__1__17_chanx_left_out[8] ,
    \cbx_1__1__17_chanx_left_out[9] ,
    \cbx_1__1__17_chanx_left_out[10] ,
    \cbx_1__1__17_chanx_left_out[11] ,
    \cbx_1__1__17_chanx_left_out[12] ,
    \cbx_1__1__17_chanx_left_out[13] ,
    \cbx_1__1__17_chanx_left_out[14] ,
    \cbx_1__1__17_chanx_left_out[15] ,
    \cbx_1__1__17_chanx_left_out[16] ,
    \cbx_1__1__17_chanx_left_out[17] ,
    \cbx_1__1__17_chanx_left_out[18] ,
    \cbx_1__1__17_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__17_chanx_left_out[0] ,
    \sb_1__1__17_chanx_left_out[1] ,
    \sb_1__1__17_chanx_left_out[2] ,
    \sb_1__1__17_chanx_left_out[3] ,
    \sb_1__1__17_chanx_left_out[4] ,
    \sb_1__1__17_chanx_left_out[5] ,
    \sb_1__1__17_chanx_left_out[6] ,
    \sb_1__1__17_chanx_left_out[7] ,
    \sb_1__1__17_chanx_left_out[8] ,
    \sb_1__1__17_chanx_left_out[9] ,
    \sb_1__1__17_chanx_left_out[10] ,
    \sb_1__1__17_chanx_left_out[11] ,
    \sb_1__1__17_chanx_left_out[12] ,
    \sb_1__1__17_chanx_left_out[13] ,
    \sb_1__1__17_chanx_left_out[14] ,
    \sb_1__1__17_chanx_left_out[15] ,
    \sb_1__1__17_chanx_left_out[16] ,
    \sb_1__1__17_chanx_left_out[17] ,
    \sb_1__1__17_chanx_left_out[18] ,
    \sb_1__1__17_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__17_chanx_right_out[0] ,
    \cbx_1__1__17_chanx_right_out[1] ,
    \cbx_1__1__17_chanx_right_out[2] ,
    \cbx_1__1__17_chanx_right_out[3] ,
    \cbx_1__1__17_chanx_right_out[4] ,
    \cbx_1__1__17_chanx_right_out[5] ,
    \cbx_1__1__17_chanx_right_out[6] ,
    \cbx_1__1__17_chanx_right_out[7] ,
    \cbx_1__1__17_chanx_right_out[8] ,
    \cbx_1__1__17_chanx_right_out[9] ,
    \cbx_1__1__17_chanx_right_out[10] ,
    \cbx_1__1__17_chanx_right_out[11] ,
    \cbx_1__1__17_chanx_right_out[12] ,
    \cbx_1__1__17_chanx_right_out[13] ,
    \cbx_1__1__17_chanx_right_out[14] ,
    \cbx_1__1__17_chanx_right_out[15] ,
    \cbx_1__1__17_chanx_right_out[16] ,
    \cbx_1__1__17_chanx_right_out[17] ,
    \cbx_1__1__17_chanx_right_out[18] ,
    \cbx_1__1__17_chanx_right_out[19] }));
 cbx_1__1_ cbx_3__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[18] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[18] ),
    .SC_IN_TOP(\scff_Wires[43] ),
    .SC_OUT_BOT(\scff_Wires[44] ),
    .bottom_grid_pin_0_(cbx_1__1__18_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__18_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__18_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__18_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__18_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__18_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__18_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__18_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__18_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__18_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__18_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__18_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__18_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__18_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__18_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__18_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__18_ccff_tail),
    .ccff_tail(cbx_1__1__18_ccff_tail),
    .clk_1_N_out(\clk_1_wires[45] ),
    .clk_1_S_out(\clk_1_wires[46] ),
    .clk_1_W_in(\clk_1_wires[44] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[84] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[45] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[46] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[44] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__11_chanx_right_out[0] ,
    \sb_1__1__11_chanx_right_out[1] ,
    \sb_1__1__11_chanx_right_out[2] ,
    \sb_1__1__11_chanx_right_out[3] ,
    \sb_1__1__11_chanx_right_out[4] ,
    \sb_1__1__11_chanx_right_out[5] ,
    \sb_1__1__11_chanx_right_out[6] ,
    \sb_1__1__11_chanx_right_out[7] ,
    \sb_1__1__11_chanx_right_out[8] ,
    \sb_1__1__11_chanx_right_out[9] ,
    \sb_1__1__11_chanx_right_out[10] ,
    \sb_1__1__11_chanx_right_out[11] ,
    \sb_1__1__11_chanx_right_out[12] ,
    \sb_1__1__11_chanx_right_out[13] ,
    \sb_1__1__11_chanx_right_out[14] ,
    \sb_1__1__11_chanx_right_out[15] ,
    \sb_1__1__11_chanx_right_out[16] ,
    \sb_1__1__11_chanx_right_out[17] ,
    \sb_1__1__11_chanx_right_out[18] ,
    \sb_1__1__11_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__18_chanx_left_out[0] ,
    \cbx_1__1__18_chanx_left_out[1] ,
    \cbx_1__1__18_chanx_left_out[2] ,
    \cbx_1__1__18_chanx_left_out[3] ,
    \cbx_1__1__18_chanx_left_out[4] ,
    \cbx_1__1__18_chanx_left_out[5] ,
    \cbx_1__1__18_chanx_left_out[6] ,
    \cbx_1__1__18_chanx_left_out[7] ,
    \cbx_1__1__18_chanx_left_out[8] ,
    \cbx_1__1__18_chanx_left_out[9] ,
    \cbx_1__1__18_chanx_left_out[10] ,
    \cbx_1__1__18_chanx_left_out[11] ,
    \cbx_1__1__18_chanx_left_out[12] ,
    \cbx_1__1__18_chanx_left_out[13] ,
    \cbx_1__1__18_chanx_left_out[14] ,
    \cbx_1__1__18_chanx_left_out[15] ,
    \cbx_1__1__18_chanx_left_out[16] ,
    \cbx_1__1__18_chanx_left_out[17] ,
    \cbx_1__1__18_chanx_left_out[18] ,
    \cbx_1__1__18_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__18_chanx_left_out[0] ,
    \sb_1__1__18_chanx_left_out[1] ,
    \sb_1__1__18_chanx_left_out[2] ,
    \sb_1__1__18_chanx_left_out[3] ,
    \sb_1__1__18_chanx_left_out[4] ,
    \sb_1__1__18_chanx_left_out[5] ,
    \sb_1__1__18_chanx_left_out[6] ,
    \sb_1__1__18_chanx_left_out[7] ,
    \sb_1__1__18_chanx_left_out[8] ,
    \sb_1__1__18_chanx_left_out[9] ,
    \sb_1__1__18_chanx_left_out[10] ,
    \sb_1__1__18_chanx_left_out[11] ,
    \sb_1__1__18_chanx_left_out[12] ,
    \sb_1__1__18_chanx_left_out[13] ,
    \sb_1__1__18_chanx_left_out[14] ,
    \sb_1__1__18_chanx_left_out[15] ,
    \sb_1__1__18_chanx_left_out[16] ,
    \sb_1__1__18_chanx_left_out[17] ,
    \sb_1__1__18_chanx_left_out[18] ,
    \sb_1__1__18_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__18_chanx_right_out[0] ,
    \cbx_1__1__18_chanx_right_out[1] ,
    \cbx_1__1__18_chanx_right_out[2] ,
    \cbx_1__1__18_chanx_right_out[3] ,
    \cbx_1__1__18_chanx_right_out[4] ,
    \cbx_1__1__18_chanx_right_out[5] ,
    \cbx_1__1__18_chanx_right_out[6] ,
    \cbx_1__1__18_chanx_right_out[7] ,
    \cbx_1__1__18_chanx_right_out[8] ,
    \cbx_1__1__18_chanx_right_out[9] ,
    \cbx_1__1__18_chanx_right_out[10] ,
    \cbx_1__1__18_chanx_right_out[11] ,
    \cbx_1__1__18_chanx_right_out[12] ,
    \cbx_1__1__18_chanx_right_out[13] ,
    \cbx_1__1__18_chanx_right_out[14] ,
    \cbx_1__1__18_chanx_right_out[15] ,
    \cbx_1__1__18_chanx_right_out[16] ,
    \cbx_1__1__18_chanx_right_out[17] ,
    \cbx_1__1__18_chanx_right_out[18] ,
    \cbx_1__1__18_chanx_right_out[19] }));
 cbx_1__1_ cbx_3__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[19] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[19] ),
    .SC_IN_TOP(\scff_Wires[41] ),
    .SC_OUT_BOT(\scff_Wires[42] ),
    .bottom_grid_pin_0_(cbx_1__1__19_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__19_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__19_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__19_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__19_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__19_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__19_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__19_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__19_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__19_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__19_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__19_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__19_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__19_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__19_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__19_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__19_ccff_tail),
    .ccff_tail(cbx_1__1__19_ccff_tail),
    .clk_2_E_out(\clk_2_wires[15] ),
    .clk_2_W_in(\clk_2_wires[14] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[87] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[15] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[14] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__12_chanx_right_out[0] ,
    \sb_1__1__12_chanx_right_out[1] ,
    \sb_1__1__12_chanx_right_out[2] ,
    \sb_1__1__12_chanx_right_out[3] ,
    \sb_1__1__12_chanx_right_out[4] ,
    \sb_1__1__12_chanx_right_out[5] ,
    \sb_1__1__12_chanx_right_out[6] ,
    \sb_1__1__12_chanx_right_out[7] ,
    \sb_1__1__12_chanx_right_out[8] ,
    \sb_1__1__12_chanx_right_out[9] ,
    \sb_1__1__12_chanx_right_out[10] ,
    \sb_1__1__12_chanx_right_out[11] ,
    \sb_1__1__12_chanx_right_out[12] ,
    \sb_1__1__12_chanx_right_out[13] ,
    \sb_1__1__12_chanx_right_out[14] ,
    \sb_1__1__12_chanx_right_out[15] ,
    \sb_1__1__12_chanx_right_out[16] ,
    \sb_1__1__12_chanx_right_out[17] ,
    \sb_1__1__12_chanx_right_out[18] ,
    \sb_1__1__12_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__19_chanx_left_out[0] ,
    \cbx_1__1__19_chanx_left_out[1] ,
    \cbx_1__1__19_chanx_left_out[2] ,
    \cbx_1__1__19_chanx_left_out[3] ,
    \cbx_1__1__19_chanx_left_out[4] ,
    \cbx_1__1__19_chanx_left_out[5] ,
    \cbx_1__1__19_chanx_left_out[6] ,
    \cbx_1__1__19_chanx_left_out[7] ,
    \cbx_1__1__19_chanx_left_out[8] ,
    \cbx_1__1__19_chanx_left_out[9] ,
    \cbx_1__1__19_chanx_left_out[10] ,
    \cbx_1__1__19_chanx_left_out[11] ,
    \cbx_1__1__19_chanx_left_out[12] ,
    \cbx_1__1__19_chanx_left_out[13] ,
    \cbx_1__1__19_chanx_left_out[14] ,
    \cbx_1__1__19_chanx_left_out[15] ,
    \cbx_1__1__19_chanx_left_out[16] ,
    \cbx_1__1__19_chanx_left_out[17] ,
    \cbx_1__1__19_chanx_left_out[18] ,
    \cbx_1__1__19_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__19_chanx_left_out[0] ,
    \sb_1__1__19_chanx_left_out[1] ,
    \sb_1__1__19_chanx_left_out[2] ,
    \sb_1__1__19_chanx_left_out[3] ,
    \sb_1__1__19_chanx_left_out[4] ,
    \sb_1__1__19_chanx_left_out[5] ,
    \sb_1__1__19_chanx_left_out[6] ,
    \sb_1__1__19_chanx_left_out[7] ,
    \sb_1__1__19_chanx_left_out[8] ,
    \sb_1__1__19_chanx_left_out[9] ,
    \sb_1__1__19_chanx_left_out[10] ,
    \sb_1__1__19_chanx_left_out[11] ,
    \sb_1__1__19_chanx_left_out[12] ,
    \sb_1__1__19_chanx_left_out[13] ,
    \sb_1__1__19_chanx_left_out[14] ,
    \sb_1__1__19_chanx_left_out[15] ,
    \sb_1__1__19_chanx_left_out[16] ,
    \sb_1__1__19_chanx_left_out[17] ,
    \sb_1__1__19_chanx_left_out[18] ,
    \sb_1__1__19_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__19_chanx_right_out[0] ,
    \cbx_1__1__19_chanx_right_out[1] ,
    \cbx_1__1__19_chanx_right_out[2] ,
    \cbx_1__1__19_chanx_right_out[3] ,
    \cbx_1__1__19_chanx_right_out[4] ,
    \cbx_1__1__19_chanx_right_out[5] ,
    \cbx_1__1__19_chanx_right_out[6] ,
    \cbx_1__1__19_chanx_right_out[7] ,
    \cbx_1__1__19_chanx_right_out[8] ,
    \cbx_1__1__19_chanx_right_out[9] ,
    \cbx_1__1__19_chanx_right_out[10] ,
    \cbx_1__1__19_chanx_right_out[11] ,
    \cbx_1__1__19_chanx_right_out[12] ,
    \cbx_1__1__19_chanx_right_out[13] ,
    \cbx_1__1__19_chanx_right_out[14] ,
    \cbx_1__1__19_chanx_right_out[15] ,
    \cbx_1__1__19_chanx_right_out[16] ,
    \cbx_1__1__19_chanx_right_out[17] ,
    \cbx_1__1__19_chanx_right_out[18] ,
    \cbx_1__1__19_chanx_right_out[19] }));
 cbx_1__1_ cbx_3__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[20] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[20] ),
    .SC_IN_TOP(\scff_Wires[39] ),
    .SC_OUT_BOT(\scff_Wires[40] ),
    .bottom_grid_pin_0_(cbx_1__1__20_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__20_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__20_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__20_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__20_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__20_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__20_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__20_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__20_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__20_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__20_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__20_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__20_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__20_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__20_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__20_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__20_ccff_tail),
    .ccff_tail(cbx_1__1__20_ccff_tail),
    .clk_1_N_out(\clk_1_wires[52] ),
    .clk_1_S_out(\clk_1_wires[53] ),
    .clk_1_W_in(\clk_1_wires[51] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[90] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[52] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[53] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[51] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__13_chanx_right_out[0] ,
    \sb_1__1__13_chanx_right_out[1] ,
    \sb_1__1__13_chanx_right_out[2] ,
    \sb_1__1__13_chanx_right_out[3] ,
    \sb_1__1__13_chanx_right_out[4] ,
    \sb_1__1__13_chanx_right_out[5] ,
    \sb_1__1__13_chanx_right_out[6] ,
    \sb_1__1__13_chanx_right_out[7] ,
    \sb_1__1__13_chanx_right_out[8] ,
    \sb_1__1__13_chanx_right_out[9] ,
    \sb_1__1__13_chanx_right_out[10] ,
    \sb_1__1__13_chanx_right_out[11] ,
    \sb_1__1__13_chanx_right_out[12] ,
    \sb_1__1__13_chanx_right_out[13] ,
    \sb_1__1__13_chanx_right_out[14] ,
    \sb_1__1__13_chanx_right_out[15] ,
    \sb_1__1__13_chanx_right_out[16] ,
    \sb_1__1__13_chanx_right_out[17] ,
    \sb_1__1__13_chanx_right_out[18] ,
    \sb_1__1__13_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__20_chanx_left_out[0] ,
    \cbx_1__1__20_chanx_left_out[1] ,
    \cbx_1__1__20_chanx_left_out[2] ,
    \cbx_1__1__20_chanx_left_out[3] ,
    \cbx_1__1__20_chanx_left_out[4] ,
    \cbx_1__1__20_chanx_left_out[5] ,
    \cbx_1__1__20_chanx_left_out[6] ,
    \cbx_1__1__20_chanx_left_out[7] ,
    \cbx_1__1__20_chanx_left_out[8] ,
    \cbx_1__1__20_chanx_left_out[9] ,
    \cbx_1__1__20_chanx_left_out[10] ,
    \cbx_1__1__20_chanx_left_out[11] ,
    \cbx_1__1__20_chanx_left_out[12] ,
    \cbx_1__1__20_chanx_left_out[13] ,
    \cbx_1__1__20_chanx_left_out[14] ,
    \cbx_1__1__20_chanx_left_out[15] ,
    \cbx_1__1__20_chanx_left_out[16] ,
    \cbx_1__1__20_chanx_left_out[17] ,
    \cbx_1__1__20_chanx_left_out[18] ,
    \cbx_1__1__20_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__20_chanx_left_out[0] ,
    \sb_1__1__20_chanx_left_out[1] ,
    \sb_1__1__20_chanx_left_out[2] ,
    \sb_1__1__20_chanx_left_out[3] ,
    \sb_1__1__20_chanx_left_out[4] ,
    \sb_1__1__20_chanx_left_out[5] ,
    \sb_1__1__20_chanx_left_out[6] ,
    \sb_1__1__20_chanx_left_out[7] ,
    \sb_1__1__20_chanx_left_out[8] ,
    \sb_1__1__20_chanx_left_out[9] ,
    \sb_1__1__20_chanx_left_out[10] ,
    \sb_1__1__20_chanx_left_out[11] ,
    \sb_1__1__20_chanx_left_out[12] ,
    \sb_1__1__20_chanx_left_out[13] ,
    \sb_1__1__20_chanx_left_out[14] ,
    \sb_1__1__20_chanx_left_out[15] ,
    \sb_1__1__20_chanx_left_out[16] ,
    \sb_1__1__20_chanx_left_out[17] ,
    \sb_1__1__20_chanx_left_out[18] ,
    \sb_1__1__20_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__20_chanx_right_out[0] ,
    \cbx_1__1__20_chanx_right_out[1] ,
    \cbx_1__1__20_chanx_right_out[2] ,
    \cbx_1__1__20_chanx_right_out[3] ,
    \cbx_1__1__20_chanx_right_out[4] ,
    \cbx_1__1__20_chanx_right_out[5] ,
    \cbx_1__1__20_chanx_right_out[6] ,
    \cbx_1__1__20_chanx_right_out[7] ,
    \cbx_1__1__20_chanx_right_out[8] ,
    \cbx_1__1__20_chanx_right_out[9] ,
    \cbx_1__1__20_chanx_right_out[10] ,
    \cbx_1__1__20_chanx_right_out[11] ,
    \cbx_1__1__20_chanx_right_out[12] ,
    \cbx_1__1__20_chanx_right_out[13] ,
    \cbx_1__1__20_chanx_right_out[14] ,
    \cbx_1__1__20_chanx_right_out[15] ,
    \cbx_1__1__20_chanx_right_out[16] ,
    \cbx_1__1__20_chanx_right_out[17] ,
    \cbx_1__1__20_chanx_right_out[18] ,
    \cbx_1__1__20_chanx_right_out[19] }));
 cbx_1__2_ cbx_3__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[37] ),
    .SC_OUT_BOT(\scff_Wires[38] ),
    .bottom_grid_pin_0_(cbx_1__8__2_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__2_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__2_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__2_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__2_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__2_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__2_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__2_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__2_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__2_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__2_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__2_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__2_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__2_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__2_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__2_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__2_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_2_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_2_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_1__8__2_ccff_tail),
    .ccff_tail(grid_io_top_2_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]),
    .prog_clk_0_S_in(\prog_clk_0_wires[93] ),
    .top_grid_pin_0_(cbx_1__8__2_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__8__1_chanx_right_out[0] ,
    \sb_1__8__1_chanx_right_out[1] ,
    \sb_1__8__1_chanx_right_out[2] ,
    \sb_1__8__1_chanx_right_out[3] ,
    \sb_1__8__1_chanx_right_out[4] ,
    \sb_1__8__1_chanx_right_out[5] ,
    \sb_1__8__1_chanx_right_out[6] ,
    \sb_1__8__1_chanx_right_out[7] ,
    \sb_1__8__1_chanx_right_out[8] ,
    \sb_1__8__1_chanx_right_out[9] ,
    \sb_1__8__1_chanx_right_out[10] ,
    \sb_1__8__1_chanx_right_out[11] ,
    \sb_1__8__1_chanx_right_out[12] ,
    \sb_1__8__1_chanx_right_out[13] ,
    \sb_1__8__1_chanx_right_out[14] ,
    \sb_1__8__1_chanx_right_out[15] ,
    \sb_1__8__1_chanx_right_out[16] ,
    \sb_1__8__1_chanx_right_out[17] ,
    \sb_1__8__1_chanx_right_out[18] ,
    \sb_1__8__1_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__2_chanx_left_out[0] ,
    \cbx_1__8__2_chanx_left_out[1] ,
    \cbx_1__8__2_chanx_left_out[2] ,
    \cbx_1__8__2_chanx_left_out[3] ,
    \cbx_1__8__2_chanx_left_out[4] ,
    \cbx_1__8__2_chanx_left_out[5] ,
    \cbx_1__8__2_chanx_left_out[6] ,
    \cbx_1__8__2_chanx_left_out[7] ,
    \cbx_1__8__2_chanx_left_out[8] ,
    \cbx_1__8__2_chanx_left_out[9] ,
    \cbx_1__8__2_chanx_left_out[10] ,
    \cbx_1__8__2_chanx_left_out[11] ,
    \cbx_1__8__2_chanx_left_out[12] ,
    \cbx_1__8__2_chanx_left_out[13] ,
    \cbx_1__8__2_chanx_left_out[14] ,
    \cbx_1__8__2_chanx_left_out[15] ,
    \cbx_1__8__2_chanx_left_out[16] ,
    \cbx_1__8__2_chanx_left_out[17] ,
    \cbx_1__8__2_chanx_left_out[18] ,
    \cbx_1__8__2_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__8__2_chanx_left_out[0] ,
    \sb_1__8__2_chanx_left_out[1] ,
    \sb_1__8__2_chanx_left_out[2] ,
    \sb_1__8__2_chanx_left_out[3] ,
    \sb_1__8__2_chanx_left_out[4] ,
    \sb_1__8__2_chanx_left_out[5] ,
    \sb_1__8__2_chanx_left_out[6] ,
    \sb_1__8__2_chanx_left_out[7] ,
    \sb_1__8__2_chanx_left_out[8] ,
    \sb_1__8__2_chanx_left_out[9] ,
    \sb_1__8__2_chanx_left_out[10] ,
    \sb_1__8__2_chanx_left_out[11] ,
    \sb_1__8__2_chanx_left_out[12] ,
    \sb_1__8__2_chanx_left_out[13] ,
    \sb_1__8__2_chanx_left_out[14] ,
    \sb_1__8__2_chanx_left_out[15] ,
    \sb_1__8__2_chanx_left_out[16] ,
    \sb_1__8__2_chanx_left_out[17] ,
    \sb_1__8__2_chanx_left_out[18] ,
    \sb_1__8__2_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__2_chanx_right_out[0] ,
    \cbx_1__8__2_chanx_right_out[1] ,
    \cbx_1__8__2_chanx_right_out[2] ,
    \cbx_1__8__2_chanx_right_out[3] ,
    \cbx_1__8__2_chanx_right_out[4] ,
    \cbx_1__8__2_chanx_right_out[5] ,
    \cbx_1__8__2_chanx_right_out[6] ,
    \cbx_1__8__2_chanx_right_out[7] ,
    \cbx_1__8__2_chanx_right_out[8] ,
    \cbx_1__8__2_chanx_right_out[9] ,
    \cbx_1__8__2_chanx_right_out[10] ,
    \cbx_1__8__2_chanx_right_out[11] ,
    \cbx_1__8__2_chanx_right_out[12] ,
    \cbx_1__8__2_chanx_right_out[13] ,
    \cbx_1__8__2_chanx_right_out[14] ,
    \cbx_1__8__2_chanx_right_out[15] ,
    \cbx_1__8__2_chanx_right_out[16] ,
    \cbx_1__8__2_chanx_right_out[17] ,
    \cbx_1__8__2_chanx_right_out[18] ,
    \cbx_1__8__2_chanx_right_out[19] }));
 cbx_1__0_ cbx_4__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[56] ),
    .SC_OUT_TOP(\scff_Wires[57] ),
    .bottom_grid_pin_0_(cbx_1__0__3_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__3_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__3_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__3_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__3_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__3_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__3_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__3_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__3_bottom_grid_pin_8_),
    .ccff_head(sb_1__0__3_ccff_tail),
    .ccff_tail(grid_io_bottom_4_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[95] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__3_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__3_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_4_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_4_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__3_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_4_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_4_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__3_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_4_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_4_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__3_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_4_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_4_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_4_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_4_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__3_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_4_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_4_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__3_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_4_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_4_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__3_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_4_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_4_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__3_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_4_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_4_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__0__2_chanx_right_out[0] ,
    \sb_1__0__2_chanx_right_out[1] ,
    \sb_1__0__2_chanx_right_out[2] ,
    \sb_1__0__2_chanx_right_out[3] ,
    \sb_1__0__2_chanx_right_out[4] ,
    \sb_1__0__2_chanx_right_out[5] ,
    \sb_1__0__2_chanx_right_out[6] ,
    \sb_1__0__2_chanx_right_out[7] ,
    \sb_1__0__2_chanx_right_out[8] ,
    \sb_1__0__2_chanx_right_out[9] ,
    \sb_1__0__2_chanx_right_out[10] ,
    \sb_1__0__2_chanx_right_out[11] ,
    \sb_1__0__2_chanx_right_out[12] ,
    \sb_1__0__2_chanx_right_out[13] ,
    \sb_1__0__2_chanx_right_out[14] ,
    \sb_1__0__2_chanx_right_out[15] ,
    \sb_1__0__2_chanx_right_out[16] ,
    \sb_1__0__2_chanx_right_out[17] ,
    \sb_1__0__2_chanx_right_out[18] ,
    \sb_1__0__2_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__3_chanx_left_out[0] ,
    \cbx_1__0__3_chanx_left_out[1] ,
    \cbx_1__0__3_chanx_left_out[2] ,
    \cbx_1__0__3_chanx_left_out[3] ,
    \cbx_1__0__3_chanx_left_out[4] ,
    \cbx_1__0__3_chanx_left_out[5] ,
    \cbx_1__0__3_chanx_left_out[6] ,
    \cbx_1__0__3_chanx_left_out[7] ,
    \cbx_1__0__3_chanx_left_out[8] ,
    \cbx_1__0__3_chanx_left_out[9] ,
    \cbx_1__0__3_chanx_left_out[10] ,
    \cbx_1__0__3_chanx_left_out[11] ,
    \cbx_1__0__3_chanx_left_out[12] ,
    \cbx_1__0__3_chanx_left_out[13] ,
    \cbx_1__0__3_chanx_left_out[14] ,
    \cbx_1__0__3_chanx_left_out[15] ,
    \cbx_1__0__3_chanx_left_out[16] ,
    \cbx_1__0__3_chanx_left_out[17] ,
    \cbx_1__0__3_chanx_left_out[18] ,
    \cbx_1__0__3_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__0__3_chanx_left_out[0] ,
    \sb_1__0__3_chanx_left_out[1] ,
    \sb_1__0__3_chanx_left_out[2] ,
    \sb_1__0__3_chanx_left_out[3] ,
    \sb_1__0__3_chanx_left_out[4] ,
    \sb_1__0__3_chanx_left_out[5] ,
    \sb_1__0__3_chanx_left_out[6] ,
    \sb_1__0__3_chanx_left_out[7] ,
    \sb_1__0__3_chanx_left_out[8] ,
    \sb_1__0__3_chanx_left_out[9] ,
    \sb_1__0__3_chanx_left_out[10] ,
    \sb_1__0__3_chanx_left_out[11] ,
    \sb_1__0__3_chanx_left_out[12] ,
    \sb_1__0__3_chanx_left_out[13] ,
    \sb_1__0__3_chanx_left_out[14] ,
    \sb_1__0__3_chanx_left_out[15] ,
    \sb_1__0__3_chanx_left_out[16] ,
    \sb_1__0__3_chanx_left_out[17] ,
    \sb_1__0__3_chanx_left_out[18] ,
    \sb_1__0__3_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__3_chanx_right_out[0] ,
    \cbx_1__0__3_chanx_right_out[1] ,
    \cbx_1__0__3_chanx_right_out[2] ,
    \cbx_1__0__3_chanx_right_out[3] ,
    \cbx_1__0__3_chanx_right_out[4] ,
    \cbx_1__0__3_chanx_right_out[5] ,
    \cbx_1__0__3_chanx_right_out[6] ,
    \cbx_1__0__3_chanx_right_out[7] ,
    \cbx_1__0__3_chanx_right_out[8] ,
    \cbx_1__0__3_chanx_right_out[9] ,
    \cbx_1__0__3_chanx_right_out[10] ,
    \cbx_1__0__3_chanx_right_out[11] ,
    \cbx_1__0__3_chanx_right_out[12] ,
    \cbx_1__0__3_chanx_right_out[13] ,
    \cbx_1__0__3_chanx_right_out[14] ,
    \cbx_1__0__3_chanx_right_out[15] ,
    \cbx_1__0__3_chanx_right_out[16] ,
    \cbx_1__0__3_chanx_right_out[17] ,
    \cbx_1__0__3_chanx_right_out[18] ,
    \cbx_1__0__3_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]}));
 cbx_1__1_ cbx_4__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[21] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[21] ),
    .SC_IN_BOT(\scff_Wires[58] ),
    .SC_OUT_TOP(\scff_Wires[59] ),
    .bottom_grid_pin_0_(cbx_1__1__21_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__21_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__21_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__21_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__21_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__21_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__21_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__21_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__21_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__21_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__21_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__21_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__21_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__21_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__21_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__21_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__21_ccff_tail),
    .ccff_tail(cbx_1__1__21_ccff_tail),
    .clk_1_N_out(\clk_1_wires[33] ),
    .clk_1_S_out(\clk_1_wires[34] ),
    .clk_1_W_in(\clk_1_wires[29] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[98] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[33] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[34] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[29] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__14_chanx_right_out[0] ,
    \sb_1__1__14_chanx_right_out[1] ,
    \sb_1__1__14_chanx_right_out[2] ,
    \sb_1__1__14_chanx_right_out[3] ,
    \sb_1__1__14_chanx_right_out[4] ,
    \sb_1__1__14_chanx_right_out[5] ,
    \sb_1__1__14_chanx_right_out[6] ,
    \sb_1__1__14_chanx_right_out[7] ,
    \sb_1__1__14_chanx_right_out[8] ,
    \sb_1__1__14_chanx_right_out[9] ,
    \sb_1__1__14_chanx_right_out[10] ,
    \sb_1__1__14_chanx_right_out[11] ,
    \sb_1__1__14_chanx_right_out[12] ,
    \sb_1__1__14_chanx_right_out[13] ,
    \sb_1__1__14_chanx_right_out[14] ,
    \sb_1__1__14_chanx_right_out[15] ,
    \sb_1__1__14_chanx_right_out[16] ,
    \sb_1__1__14_chanx_right_out[17] ,
    \sb_1__1__14_chanx_right_out[18] ,
    \sb_1__1__14_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__21_chanx_left_out[0] ,
    \cbx_1__1__21_chanx_left_out[1] ,
    \cbx_1__1__21_chanx_left_out[2] ,
    \cbx_1__1__21_chanx_left_out[3] ,
    \cbx_1__1__21_chanx_left_out[4] ,
    \cbx_1__1__21_chanx_left_out[5] ,
    \cbx_1__1__21_chanx_left_out[6] ,
    \cbx_1__1__21_chanx_left_out[7] ,
    \cbx_1__1__21_chanx_left_out[8] ,
    \cbx_1__1__21_chanx_left_out[9] ,
    \cbx_1__1__21_chanx_left_out[10] ,
    \cbx_1__1__21_chanx_left_out[11] ,
    \cbx_1__1__21_chanx_left_out[12] ,
    \cbx_1__1__21_chanx_left_out[13] ,
    \cbx_1__1__21_chanx_left_out[14] ,
    \cbx_1__1__21_chanx_left_out[15] ,
    \cbx_1__1__21_chanx_left_out[16] ,
    \cbx_1__1__21_chanx_left_out[17] ,
    \cbx_1__1__21_chanx_left_out[18] ,
    \cbx_1__1__21_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__21_chanx_left_out[0] ,
    \sb_1__1__21_chanx_left_out[1] ,
    \sb_1__1__21_chanx_left_out[2] ,
    \sb_1__1__21_chanx_left_out[3] ,
    \sb_1__1__21_chanx_left_out[4] ,
    \sb_1__1__21_chanx_left_out[5] ,
    \sb_1__1__21_chanx_left_out[6] ,
    \sb_1__1__21_chanx_left_out[7] ,
    \sb_1__1__21_chanx_left_out[8] ,
    \sb_1__1__21_chanx_left_out[9] ,
    \sb_1__1__21_chanx_left_out[10] ,
    \sb_1__1__21_chanx_left_out[11] ,
    \sb_1__1__21_chanx_left_out[12] ,
    \sb_1__1__21_chanx_left_out[13] ,
    \sb_1__1__21_chanx_left_out[14] ,
    \sb_1__1__21_chanx_left_out[15] ,
    \sb_1__1__21_chanx_left_out[16] ,
    \sb_1__1__21_chanx_left_out[17] ,
    \sb_1__1__21_chanx_left_out[18] ,
    \sb_1__1__21_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__21_chanx_right_out[0] ,
    \cbx_1__1__21_chanx_right_out[1] ,
    \cbx_1__1__21_chanx_right_out[2] ,
    \cbx_1__1__21_chanx_right_out[3] ,
    \cbx_1__1__21_chanx_right_out[4] ,
    \cbx_1__1__21_chanx_right_out[5] ,
    \cbx_1__1__21_chanx_right_out[6] ,
    \cbx_1__1__21_chanx_right_out[7] ,
    \cbx_1__1__21_chanx_right_out[8] ,
    \cbx_1__1__21_chanx_right_out[9] ,
    \cbx_1__1__21_chanx_right_out[10] ,
    \cbx_1__1__21_chanx_right_out[11] ,
    \cbx_1__1__21_chanx_right_out[12] ,
    \cbx_1__1__21_chanx_right_out[13] ,
    \cbx_1__1__21_chanx_right_out[14] ,
    \cbx_1__1__21_chanx_right_out[15] ,
    \cbx_1__1__21_chanx_right_out[16] ,
    \cbx_1__1__21_chanx_right_out[17] ,
    \cbx_1__1__21_chanx_right_out[18] ,
    \cbx_1__1__21_chanx_right_out[19] }));
 cbx_1__1_ cbx_4__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[22] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[22] ),
    .SC_IN_BOT(\scff_Wires[60] ),
    .SC_OUT_TOP(\scff_Wires[61] ),
    .bottom_grid_pin_0_(cbx_1__1__22_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__22_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__22_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__22_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__22_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__22_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__22_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__22_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__22_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__22_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__22_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__22_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__22_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__22_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__22_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__22_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__22_ccff_tail),
    .ccff_tail(cbx_1__1__22_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[101] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__15_chanx_right_out[0] ,
    \sb_1__1__15_chanx_right_out[1] ,
    \sb_1__1__15_chanx_right_out[2] ,
    \sb_1__1__15_chanx_right_out[3] ,
    \sb_1__1__15_chanx_right_out[4] ,
    \sb_1__1__15_chanx_right_out[5] ,
    \sb_1__1__15_chanx_right_out[6] ,
    \sb_1__1__15_chanx_right_out[7] ,
    \sb_1__1__15_chanx_right_out[8] ,
    \sb_1__1__15_chanx_right_out[9] ,
    \sb_1__1__15_chanx_right_out[10] ,
    \sb_1__1__15_chanx_right_out[11] ,
    \sb_1__1__15_chanx_right_out[12] ,
    \sb_1__1__15_chanx_right_out[13] ,
    \sb_1__1__15_chanx_right_out[14] ,
    \sb_1__1__15_chanx_right_out[15] ,
    \sb_1__1__15_chanx_right_out[16] ,
    \sb_1__1__15_chanx_right_out[17] ,
    \sb_1__1__15_chanx_right_out[18] ,
    \sb_1__1__15_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__22_chanx_left_out[0] ,
    \cbx_1__1__22_chanx_left_out[1] ,
    \cbx_1__1__22_chanx_left_out[2] ,
    \cbx_1__1__22_chanx_left_out[3] ,
    \cbx_1__1__22_chanx_left_out[4] ,
    \cbx_1__1__22_chanx_left_out[5] ,
    \cbx_1__1__22_chanx_left_out[6] ,
    \cbx_1__1__22_chanx_left_out[7] ,
    \cbx_1__1__22_chanx_left_out[8] ,
    \cbx_1__1__22_chanx_left_out[9] ,
    \cbx_1__1__22_chanx_left_out[10] ,
    \cbx_1__1__22_chanx_left_out[11] ,
    \cbx_1__1__22_chanx_left_out[12] ,
    \cbx_1__1__22_chanx_left_out[13] ,
    \cbx_1__1__22_chanx_left_out[14] ,
    \cbx_1__1__22_chanx_left_out[15] ,
    \cbx_1__1__22_chanx_left_out[16] ,
    \cbx_1__1__22_chanx_left_out[17] ,
    \cbx_1__1__22_chanx_left_out[18] ,
    \cbx_1__1__22_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__22_chanx_left_out[0] ,
    \sb_1__1__22_chanx_left_out[1] ,
    \sb_1__1__22_chanx_left_out[2] ,
    \sb_1__1__22_chanx_left_out[3] ,
    \sb_1__1__22_chanx_left_out[4] ,
    \sb_1__1__22_chanx_left_out[5] ,
    \sb_1__1__22_chanx_left_out[6] ,
    \sb_1__1__22_chanx_left_out[7] ,
    \sb_1__1__22_chanx_left_out[8] ,
    \sb_1__1__22_chanx_left_out[9] ,
    \sb_1__1__22_chanx_left_out[10] ,
    \sb_1__1__22_chanx_left_out[11] ,
    \sb_1__1__22_chanx_left_out[12] ,
    \sb_1__1__22_chanx_left_out[13] ,
    \sb_1__1__22_chanx_left_out[14] ,
    \sb_1__1__22_chanx_left_out[15] ,
    \sb_1__1__22_chanx_left_out[16] ,
    \sb_1__1__22_chanx_left_out[17] ,
    \sb_1__1__22_chanx_left_out[18] ,
    \sb_1__1__22_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__22_chanx_right_out[0] ,
    \cbx_1__1__22_chanx_right_out[1] ,
    \cbx_1__1__22_chanx_right_out[2] ,
    \cbx_1__1__22_chanx_right_out[3] ,
    \cbx_1__1__22_chanx_right_out[4] ,
    \cbx_1__1__22_chanx_right_out[5] ,
    \cbx_1__1__22_chanx_right_out[6] ,
    \cbx_1__1__22_chanx_right_out[7] ,
    \cbx_1__1__22_chanx_right_out[8] ,
    \cbx_1__1__22_chanx_right_out[9] ,
    \cbx_1__1__22_chanx_right_out[10] ,
    \cbx_1__1__22_chanx_right_out[11] ,
    \cbx_1__1__22_chanx_right_out[12] ,
    \cbx_1__1__22_chanx_right_out[13] ,
    \cbx_1__1__22_chanx_right_out[14] ,
    \cbx_1__1__22_chanx_right_out[15] ,
    \cbx_1__1__22_chanx_right_out[16] ,
    \cbx_1__1__22_chanx_right_out[17] ,
    \cbx_1__1__22_chanx_right_out[18] ,
    \cbx_1__1__22_chanx_right_out[19] }));
 cbx_1__1_ cbx_4__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[23] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[23] ),
    .SC_IN_BOT(\scff_Wires[62] ),
    .SC_OUT_TOP(\scff_Wires[63] ),
    .bottom_grid_pin_0_(cbx_1__1__23_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__23_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__23_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__23_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__23_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__23_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__23_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__23_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__23_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__23_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__23_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__23_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__23_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__23_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__23_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__23_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__23_ccff_tail),
    .ccff_tail(cbx_1__1__23_ccff_tail),
    .clk_1_N_out(\clk_1_wires[40] ),
    .clk_1_S_out(\clk_1_wires[41] ),
    .clk_1_W_in(\clk_1_wires[36] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[104] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[40] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[41] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[36] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__16_chanx_right_out[0] ,
    \sb_1__1__16_chanx_right_out[1] ,
    \sb_1__1__16_chanx_right_out[2] ,
    \sb_1__1__16_chanx_right_out[3] ,
    \sb_1__1__16_chanx_right_out[4] ,
    \sb_1__1__16_chanx_right_out[5] ,
    \sb_1__1__16_chanx_right_out[6] ,
    \sb_1__1__16_chanx_right_out[7] ,
    \sb_1__1__16_chanx_right_out[8] ,
    \sb_1__1__16_chanx_right_out[9] ,
    \sb_1__1__16_chanx_right_out[10] ,
    \sb_1__1__16_chanx_right_out[11] ,
    \sb_1__1__16_chanx_right_out[12] ,
    \sb_1__1__16_chanx_right_out[13] ,
    \sb_1__1__16_chanx_right_out[14] ,
    \sb_1__1__16_chanx_right_out[15] ,
    \sb_1__1__16_chanx_right_out[16] ,
    \sb_1__1__16_chanx_right_out[17] ,
    \sb_1__1__16_chanx_right_out[18] ,
    \sb_1__1__16_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__23_chanx_left_out[0] ,
    \cbx_1__1__23_chanx_left_out[1] ,
    \cbx_1__1__23_chanx_left_out[2] ,
    \cbx_1__1__23_chanx_left_out[3] ,
    \cbx_1__1__23_chanx_left_out[4] ,
    \cbx_1__1__23_chanx_left_out[5] ,
    \cbx_1__1__23_chanx_left_out[6] ,
    \cbx_1__1__23_chanx_left_out[7] ,
    \cbx_1__1__23_chanx_left_out[8] ,
    \cbx_1__1__23_chanx_left_out[9] ,
    \cbx_1__1__23_chanx_left_out[10] ,
    \cbx_1__1__23_chanx_left_out[11] ,
    \cbx_1__1__23_chanx_left_out[12] ,
    \cbx_1__1__23_chanx_left_out[13] ,
    \cbx_1__1__23_chanx_left_out[14] ,
    \cbx_1__1__23_chanx_left_out[15] ,
    \cbx_1__1__23_chanx_left_out[16] ,
    \cbx_1__1__23_chanx_left_out[17] ,
    \cbx_1__1__23_chanx_left_out[18] ,
    \cbx_1__1__23_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__23_chanx_left_out[0] ,
    \sb_1__1__23_chanx_left_out[1] ,
    \sb_1__1__23_chanx_left_out[2] ,
    \sb_1__1__23_chanx_left_out[3] ,
    \sb_1__1__23_chanx_left_out[4] ,
    \sb_1__1__23_chanx_left_out[5] ,
    \sb_1__1__23_chanx_left_out[6] ,
    \sb_1__1__23_chanx_left_out[7] ,
    \sb_1__1__23_chanx_left_out[8] ,
    \sb_1__1__23_chanx_left_out[9] ,
    \sb_1__1__23_chanx_left_out[10] ,
    \sb_1__1__23_chanx_left_out[11] ,
    \sb_1__1__23_chanx_left_out[12] ,
    \sb_1__1__23_chanx_left_out[13] ,
    \sb_1__1__23_chanx_left_out[14] ,
    \sb_1__1__23_chanx_left_out[15] ,
    \sb_1__1__23_chanx_left_out[16] ,
    \sb_1__1__23_chanx_left_out[17] ,
    \sb_1__1__23_chanx_left_out[18] ,
    \sb_1__1__23_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__23_chanx_right_out[0] ,
    \cbx_1__1__23_chanx_right_out[1] ,
    \cbx_1__1__23_chanx_right_out[2] ,
    \cbx_1__1__23_chanx_right_out[3] ,
    \cbx_1__1__23_chanx_right_out[4] ,
    \cbx_1__1__23_chanx_right_out[5] ,
    \cbx_1__1__23_chanx_right_out[6] ,
    \cbx_1__1__23_chanx_right_out[7] ,
    \cbx_1__1__23_chanx_right_out[8] ,
    \cbx_1__1__23_chanx_right_out[9] ,
    \cbx_1__1__23_chanx_right_out[10] ,
    \cbx_1__1__23_chanx_right_out[11] ,
    \cbx_1__1__23_chanx_right_out[12] ,
    \cbx_1__1__23_chanx_right_out[13] ,
    \cbx_1__1__23_chanx_right_out[14] ,
    \cbx_1__1__23_chanx_right_out[15] ,
    \cbx_1__1__23_chanx_right_out[16] ,
    \cbx_1__1__23_chanx_right_out[17] ,
    \cbx_1__1__23_chanx_right_out[18] ,
    \cbx_1__1__23_chanx_right_out[19] }));
 cbx_1__1_ cbx_4__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[24] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[24] ),
    .SC_IN_BOT(\scff_Wires[64] ),
    .SC_OUT_TOP(\scff_Wires[65] ),
    .bottom_grid_pin_0_(cbx_1__1__24_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__24_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__24_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__24_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__24_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__24_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__24_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__24_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__24_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__24_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__24_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__24_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__24_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__24_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__24_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__24_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__24_ccff_tail),
    .ccff_tail(cbx_1__1__24_ccff_tail),
    .clk_3_W_in(\clk_3_wires[3] ),
    .clk_3_W_out(\clk_3_wires[4] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[107] ),
    .prog_clk_3_W_in(\prog_clk_3_wires[3] ),
    .prog_clk_3_W_out(\prog_clk_3_wires[4] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__17_chanx_right_out[0] ,
    \sb_1__1__17_chanx_right_out[1] ,
    \sb_1__1__17_chanx_right_out[2] ,
    \sb_1__1__17_chanx_right_out[3] ,
    \sb_1__1__17_chanx_right_out[4] ,
    \sb_1__1__17_chanx_right_out[5] ,
    \sb_1__1__17_chanx_right_out[6] ,
    \sb_1__1__17_chanx_right_out[7] ,
    \sb_1__1__17_chanx_right_out[8] ,
    \sb_1__1__17_chanx_right_out[9] ,
    \sb_1__1__17_chanx_right_out[10] ,
    \sb_1__1__17_chanx_right_out[11] ,
    \sb_1__1__17_chanx_right_out[12] ,
    \sb_1__1__17_chanx_right_out[13] ,
    \sb_1__1__17_chanx_right_out[14] ,
    \sb_1__1__17_chanx_right_out[15] ,
    \sb_1__1__17_chanx_right_out[16] ,
    \sb_1__1__17_chanx_right_out[17] ,
    \sb_1__1__17_chanx_right_out[18] ,
    \sb_1__1__17_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__24_chanx_left_out[0] ,
    \cbx_1__1__24_chanx_left_out[1] ,
    \cbx_1__1__24_chanx_left_out[2] ,
    \cbx_1__1__24_chanx_left_out[3] ,
    \cbx_1__1__24_chanx_left_out[4] ,
    \cbx_1__1__24_chanx_left_out[5] ,
    \cbx_1__1__24_chanx_left_out[6] ,
    \cbx_1__1__24_chanx_left_out[7] ,
    \cbx_1__1__24_chanx_left_out[8] ,
    \cbx_1__1__24_chanx_left_out[9] ,
    \cbx_1__1__24_chanx_left_out[10] ,
    \cbx_1__1__24_chanx_left_out[11] ,
    \cbx_1__1__24_chanx_left_out[12] ,
    \cbx_1__1__24_chanx_left_out[13] ,
    \cbx_1__1__24_chanx_left_out[14] ,
    \cbx_1__1__24_chanx_left_out[15] ,
    \cbx_1__1__24_chanx_left_out[16] ,
    \cbx_1__1__24_chanx_left_out[17] ,
    \cbx_1__1__24_chanx_left_out[18] ,
    \cbx_1__1__24_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__24_chanx_left_out[0] ,
    \sb_1__1__24_chanx_left_out[1] ,
    \sb_1__1__24_chanx_left_out[2] ,
    \sb_1__1__24_chanx_left_out[3] ,
    \sb_1__1__24_chanx_left_out[4] ,
    \sb_1__1__24_chanx_left_out[5] ,
    \sb_1__1__24_chanx_left_out[6] ,
    \sb_1__1__24_chanx_left_out[7] ,
    \sb_1__1__24_chanx_left_out[8] ,
    \sb_1__1__24_chanx_left_out[9] ,
    \sb_1__1__24_chanx_left_out[10] ,
    \sb_1__1__24_chanx_left_out[11] ,
    \sb_1__1__24_chanx_left_out[12] ,
    \sb_1__1__24_chanx_left_out[13] ,
    \sb_1__1__24_chanx_left_out[14] ,
    \sb_1__1__24_chanx_left_out[15] ,
    \sb_1__1__24_chanx_left_out[16] ,
    \sb_1__1__24_chanx_left_out[17] ,
    \sb_1__1__24_chanx_left_out[18] ,
    \sb_1__1__24_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__24_chanx_right_out[0] ,
    \cbx_1__1__24_chanx_right_out[1] ,
    \cbx_1__1__24_chanx_right_out[2] ,
    \cbx_1__1__24_chanx_right_out[3] ,
    \cbx_1__1__24_chanx_right_out[4] ,
    \cbx_1__1__24_chanx_right_out[5] ,
    \cbx_1__1__24_chanx_right_out[6] ,
    \cbx_1__1__24_chanx_right_out[7] ,
    \cbx_1__1__24_chanx_right_out[8] ,
    \cbx_1__1__24_chanx_right_out[9] ,
    \cbx_1__1__24_chanx_right_out[10] ,
    \cbx_1__1__24_chanx_right_out[11] ,
    \cbx_1__1__24_chanx_right_out[12] ,
    \cbx_1__1__24_chanx_right_out[13] ,
    \cbx_1__1__24_chanx_right_out[14] ,
    \cbx_1__1__24_chanx_right_out[15] ,
    \cbx_1__1__24_chanx_right_out[16] ,
    \cbx_1__1__24_chanx_right_out[17] ,
    \cbx_1__1__24_chanx_right_out[18] ,
    \cbx_1__1__24_chanx_right_out[19] }));
 cbx_1__1_ cbx_4__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[25] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[25] ),
    .SC_IN_BOT(\scff_Wires[66] ),
    .SC_OUT_TOP(\scff_Wires[67] ),
    .bottom_grid_pin_0_(cbx_1__1__25_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__25_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__25_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__25_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__25_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__25_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__25_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__25_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__25_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__25_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__25_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__25_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__25_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__25_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__25_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__25_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__25_ccff_tail),
    .ccff_tail(cbx_1__1__25_ccff_tail),
    .clk_1_N_out(\clk_1_wires[47] ),
    .clk_1_S_out(\clk_1_wires[48] ),
    .clk_1_W_in(\clk_1_wires[43] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[110] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[47] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[48] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[43] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__18_chanx_right_out[0] ,
    \sb_1__1__18_chanx_right_out[1] ,
    \sb_1__1__18_chanx_right_out[2] ,
    \sb_1__1__18_chanx_right_out[3] ,
    \sb_1__1__18_chanx_right_out[4] ,
    \sb_1__1__18_chanx_right_out[5] ,
    \sb_1__1__18_chanx_right_out[6] ,
    \sb_1__1__18_chanx_right_out[7] ,
    \sb_1__1__18_chanx_right_out[8] ,
    \sb_1__1__18_chanx_right_out[9] ,
    \sb_1__1__18_chanx_right_out[10] ,
    \sb_1__1__18_chanx_right_out[11] ,
    \sb_1__1__18_chanx_right_out[12] ,
    \sb_1__1__18_chanx_right_out[13] ,
    \sb_1__1__18_chanx_right_out[14] ,
    \sb_1__1__18_chanx_right_out[15] ,
    \sb_1__1__18_chanx_right_out[16] ,
    \sb_1__1__18_chanx_right_out[17] ,
    \sb_1__1__18_chanx_right_out[18] ,
    \sb_1__1__18_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__25_chanx_left_out[0] ,
    \cbx_1__1__25_chanx_left_out[1] ,
    \cbx_1__1__25_chanx_left_out[2] ,
    \cbx_1__1__25_chanx_left_out[3] ,
    \cbx_1__1__25_chanx_left_out[4] ,
    \cbx_1__1__25_chanx_left_out[5] ,
    \cbx_1__1__25_chanx_left_out[6] ,
    \cbx_1__1__25_chanx_left_out[7] ,
    \cbx_1__1__25_chanx_left_out[8] ,
    \cbx_1__1__25_chanx_left_out[9] ,
    \cbx_1__1__25_chanx_left_out[10] ,
    \cbx_1__1__25_chanx_left_out[11] ,
    \cbx_1__1__25_chanx_left_out[12] ,
    \cbx_1__1__25_chanx_left_out[13] ,
    \cbx_1__1__25_chanx_left_out[14] ,
    \cbx_1__1__25_chanx_left_out[15] ,
    \cbx_1__1__25_chanx_left_out[16] ,
    \cbx_1__1__25_chanx_left_out[17] ,
    \cbx_1__1__25_chanx_left_out[18] ,
    \cbx_1__1__25_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__25_chanx_left_out[0] ,
    \sb_1__1__25_chanx_left_out[1] ,
    \sb_1__1__25_chanx_left_out[2] ,
    \sb_1__1__25_chanx_left_out[3] ,
    \sb_1__1__25_chanx_left_out[4] ,
    \sb_1__1__25_chanx_left_out[5] ,
    \sb_1__1__25_chanx_left_out[6] ,
    \sb_1__1__25_chanx_left_out[7] ,
    \sb_1__1__25_chanx_left_out[8] ,
    \sb_1__1__25_chanx_left_out[9] ,
    \sb_1__1__25_chanx_left_out[10] ,
    \sb_1__1__25_chanx_left_out[11] ,
    \sb_1__1__25_chanx_left_out[12] ,
    \sb_1__1__25_chanx_left_out[13] ,
    \sb_1__1__25_chanx_left_out[14] ,
    \sb_1__1__25_chanx_left_out[15] ,
    \sb_1__1__25_chanx_left_out[16] ,
    \sb_1__1__25_chanx_left_out[17] ,
    \sb_1__1__25_chanx_left_out[18] ,
    \sb_1__1__25_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__25_chanx_right_out[0] ,
    \cbx_1__1__25_chanx_right_out[1] ,
    \cbx_1__1__25_chanx_right_out[2] ,
    \cbx_1__1__25_chanx_right_out[3] ,
    \cbx_1__1__25_chanx_right_out[4] ,
    \cbx_1__1__25_chanx_right_out[5] ,
    \cbx_1__1__25_chanx_right_out[6] ,
    \cbx_1__1__25_chanx_right_out[7] ,
    \cbx_1__1__25_chanx_right_out[8] ,
    \cbx_1__1__25_chanx_right_out[9] ,
    \cbx_1__1__25_chanx_right_out[10] ,
    \cbx_1__1__25_chanx_right_out[11] ,
    \cbx_1__1__25_chanx_right_out[12] ,
    \cbx_1__1__25_chanx_right_out[13] ,
    \cbx_1__1__25_chanx_right_out[14] ,
    \cbx_1__1__25_chanx_right_out[15] ,
    \cbx_1__1__25_chanx_right_out[16] ,
    \cbx_1__1__25_chanx_right_out[17] ,
    \cbx_1__1__25_chanx_right_out[18] ,
    \cbx_1__1__25_chanx_right_out[19] }));
 cbx_1__1_ cbx_4__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[26] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[26] ),
    .SC_IN_BOT(\scff_Wires[68] ),
    .SC_OUT_TOP(\scff_Wires[69] ),
    .bottom_grid_pin_0_(cbx_1__1__26_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__26_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__26_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__26_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__26_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__26_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__26_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__26_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__26_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__26_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__26_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__26_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__26_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__26_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__26_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__26_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__26_ccff_tail),
    .ccff_tail(cbx_1__1__26_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[113] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__19_chanx_right_out[0] ,
    \sb_1__1__19_chanx_right_out[1] ,
    \sb_1__1__19_chanx_right_out[2] ,
    \sb_1__1__19_chanx_right_out[3] ,
    \sb_1__1__19_chanx_right_out[4] ,
    \sb_1__1__19_chanx_right_out[5] ,
    \sb_1__1__19_chanx_right_out[6] ,
    \sb_1__1__19_chanx_right_out[7] ,
    \sb_1__1__19_chanx_right_out[8] ,
    \sb_1__1__19_chanx_right_out[9] ,
    \sb_1__1__19_chanx_right_out[10] ,
    \sb_1__1__19_chanx_right_out[11] ,
    \sb_1__1__19_chanx_right_out[12] ,
    \sb_1__1__19_chanx_right_out[13] ,
    \sb_1__1__19_chanx_right_out[14] ,
    \sb_1__1__19_chanx_right_out[15] ,
    \sb_1__1__19_chanx_right_out[16] ,
    \sb_1__1__19_chanx_right_out[17] ,
    \sb_1__1__19_chanx_right_out[18] ,
    \sb_1__1__19_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__26_chanx_left_out[0] ,
    \cbx_1__1__26_chanx_left_out[1] ,
    \cbx_1__1__26_chanx_left_out[2] ,
    \cbx_1__1__26_chanx_left_out[3] ,
    \cbx_1__1__26_chanx_left_out[4] ,
    \cbx_1__1__26_chanx_left_out[5] ,
    \cbx_1__1__26_chanx_left_out[6] ,
    \cbx_1__1__26_chanx_left_out[7] ,
    \cbx_1__1__26_chanx_left_out[8] ,
    \cbx_1__1__26_chanx_left_out[9] ,
    \cbx_1__1__26_chanx_left_out[10] ,
    \cbx_1__1__26_chanx_left_out[11] ,
    \cbx_1__1__26_chanx_left_out[12] ,
    \cbx_1__1__26_chanx_left_out[13] ,
    \cbx_1__1__26_chanx_left_out[14] ,
    \cbx_1__1__26_chanx_left_out[15] ,
    \cbx_1__1__26_chanx_left_out[16] ,
    \cbx_1__1__26_chanx_left_out[17] ,
    \cbx_1__1__26_chanx_left_out[18] ,
    \cbx_1__1__26_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__26_chanx_left_out[0] ,
    \sb_1__1__26_chanx_left_out[1] ,
    \sb_1__1__26_chanx_left_out[2] ,
    \sb_1__1__26_chanx_left_out[3] ,
    \sb_1__1__26_chanx_left_out[4] ,
    \sb_1__1__26_chanx_left_out[5] ,
    \sb_1__1__26_chanx_left_out[6] ,
    \sb_1__1__26_chanx_left_out[7] ,
    \sb_1__1__26_chanx_left_out[8] ,
    \sb_1__1__26_chanx_left_out[9] ,
    \sb_1__1__26_chanx_left_out[10] ,
    \sb_1__1__26_chanx_left_out[11] ,
    \sb_1__1__26_chanx_left_out[12] ,
    \sb_1__1__26_chanx_left_out[13] ,
    \sb_1__1__26_chanx_left_out[14] ,
    \sb_1__1__26_chanx_left_out[15] ,
    \sb_1__1__26_chanx_left_out[16] ,
    \sb_1__1__26_chanx_left_out[17] ,
    \sb_1__1__26_chanx_left_out[18] ,
    \sb_1__1__26_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__26_chanx_right_out[0] ,
    \cbx_1__1__26_chanx_right_out[1] ,
    \cbx_1__1__26_chanx_right_out[2] ,
    \cbx_1__1__26_chanx_right_out[3] ,
    \cbx_1__1__26_chanx_right_out[4] ,
    \cbx_1__1__26_chanx_right_out[5] ,
    \cbx_1__1__26_chanx_right_out[6] ,
    \cbx_1__1__26_chanx_right_out[7] ,
    \cbx_1__1__26_chanx_right_out[8] ,
    \cbx_1__1__26_chanx_right_out[9] ,
    \cbx_1__1__26_chanx_right_out[10] ,
    \cbx_1__1__26_chanx_right_out[11] ,
    \cbx_1__1__26_chanx_right_out[12] ,
    \cbx_1__1__26_chanx_right_out[13] ,
    \cbx_1__1__26_chanx_right_out[14] ,
    \cbx_1__1__26_chanx_right_out[15] ,
    \cbx_1__1__26_chanx_right_out[16] ,
    \cbx_1__1__26_chanx_right_out[17] ,
    \cbx_1__1__26_chanx_right_out[18] ,
    \cbx_1__1__26_chanx_right_out[19] }));
 cbx_1__1_ cbx_4__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[27] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[27] ),
    .SC_IN_BOT(\scff_Wires[70] ),
    .SC_OUT_TOP(\scff_Wires[71] ),
    .bottom_grid_pin_0_(cbx_1__1__27_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__27_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__27_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__27_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__27_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__27_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__27_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__27_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__27_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__27_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__27_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__27_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__27_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__27_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__27_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__27_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__27_ccff_tail),
    .ccff_tail(cbx_1__1__27_ccff_tail),
    .clk_1_N_out(\clk_1_wires[54] ),
    .clk_1_S_out(\clk_1_wires[55] ),
    .clk_1_W_in(\clk_1_wires[50] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[116] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[54] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[55] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[50] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__20_chanx_right_out[0] ,
    \sb_1__1__20_chanx_right_out[1] ,
    \sb_1__1__20_chanx_right_out[2] ,
    \sb_1__1__20_chanx_right_out[3] ,
    \sb_1__1__20_chanx_right_out[4] ,
    \sb_1__1__20_chanx_right_out[5] ,
    \sb_1__1__20_chanx_right_out[6] ,
    \sb_1__1__20_chanx_right_out[7] ,
    \sb_1__1__20_chanx_right_out[8] ,
    \sb_1__1__20_chanx_right_out[9] ,
    \sb_1__1__20_chanx_right_out[10] ,
    \sb_1__1__20_chanx_right_out[11] ,
    \sb_1__1__20_chanx_right_out[12] ,
    \sb_1__1__20_chanx_right_out[13] ,
    \sb_1__1__20_chanx_right_out[14] ,
    \sb_1__1__20_chanx_right_out[15] ,
    \sb_1__1__20_chanx_right_out[16] ,
    \sb_1__1__20_chanx_right_out[17] ,
    \sb_1__1__20_chanx_right_out[18] ,
    \sb_1__1__20_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__27_chanx_left_out[0] ,
    \cbx_1__1__27_chanx_left_out[1] ,
    \cbx_1__1__27_chanx_left_out[2] ,
    \cbx_1__1__27_chanx_left_out[3] ,
    \cbx_1__1__27_chanx_left_out[4] ,
    \cbx_1__1__27_chanx_left_out[5] ,
    \cbx_1__1__27_chanx_left_out[6] ,
    \cbx_1__1__27_chanx_left_out[7] ,
    \cbx_1__1__27_chanx_left_out[8] ,
    \cbx_1__1__27_chanx_left_out[9] ,
    \cbx_1__1__27_chanx_left_out[10] ,
    \cbx_1__1__27_chanx_left_out[11] ,
    \cbx_1__1__27_chanx_left_out[12] ,
    \cbx_1__1__27_chanx_left_out[13] ,
    \cbx_1__1__27_chanx_left_out[14] ,
    \cbx_1__1__27_chanx_left_out[15] ,
    \cbx_1__1__27_chanx_left_out[16] ,
    \cbx_1__1__27_chanx_left_out[17] ,
    \cbx_1__1__27_chanx_left_out[18] ,
    \cbx_1__1__27_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__27_chanx_left_out[0] ,
    \sb_1__1__27_chanx_left_out[1] ,
    \sb_1__1__27_chanx_left_out[2] ,
    \sb_1__1__27_chanx_left_out[3] ,
    \sb_1__1__27_chanx_left_out[4] ,
    \sb_1__1__27_chanx_left_out[5] ,
    \sb_1__1__27_chanx_left_out[6] ,
    \sb_1__1__27_chanx_left_out[7] ,
    \sb_1__1__27_chanx_left_out[8] ,
    \sb_1__1__27_chanx_left_out[9] ,
    \sb_1__1__27_chanx_left_out[10] ,
    \sb_1__1__27_chanx_left_out[11] ,
    \sb_1__1__27_chanx_left_out[12] ,
    \sb_1__1__27_chanx_left_out[13] ,
    \sb_1__1__27_chanx_left_out[14] ,
    \sb_1__1__27_chanx_left_out[15] ,
    \sb_1__1__27_chanx_left_out[16] ,
    \sb_1__1__27_chanx_left_out[17] ,
    \sb_1__1__27_chanx_left_out[18] ,
    \sb_1__1__27_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__27_chanx_right_out[0] ,
    \cbx_1__1__27_chanx_right_out[1] ,
    \cbx_1__1__27_chanx_right_out[2] ,
    \cbx_1__1__27_chanx_right_out[3] ,
    \cbx_1__1__27_chanx_right_out[4] ,
    \cbx_1__1__27_chanx_right_out[5] ,
    \cbx_1__1__27_chanx_right_out[6] ,
    \cbx_1__1__27_chanx_right_out[7] ,
    \cbx_1__1__27_chanx_right_out[8] ,
    \cbx_1__1__27_chanx_right_out[9] ,
    \cbx_1__1__27_chanx_right_out[10] ,
    \cbx_1__1__27_chanx_right_out[11] ,
    \cbx_1__1__27_chanx_right_out[12] ,
    \cbx_1__1__27_chanx_right_out[13] ,
    \cbx_1__1__27_chanx_right_out[14] ,
    \cbx_1__1__27_chanx_right_out[15] ,
    \cbx_1__1__27_chanx_right_out[16] ,
    \cbx_1__1__27_chanx_right_out[17] ,
    \cbx_1__1__27_chanx_right_out[18] ,
    \cbx_1__1__27_chanx_right_out[19] }));
 cbx_1__2_ cbx_4__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[72] ),
    .SC_OUT_TOP(\scff_Wires[73] ),
    .bottom_grid_pin_0_(cbx_1__8__3_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__3_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__3_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__3_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__3_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__3_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__3_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__3_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__3_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__3_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__3_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__3_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__3_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__3_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__3_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__3_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__3_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_3_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_3_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_1__8__3_ccff_tail),
    .ccff_tail(grid_io_top_3_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]),
    .prog_clk_0_S_in(\prog_clk_0_wires[119] ),
    .top_grid_pin_0_(cbx_1__8__3_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__8__2_chanx_right_out[0] ,
    \sb_1__8__2_chanx_right_out[1] ,
    \sb_1__8__2_chanx_right_out[2] ,
    \sb_1__8__2_chanx_right_out[3] ,
    \sb_1__8__2_chanx_right_out[4] ,
    \sb_1__8__2_chanx_right_out[5] ,
    \sb_1__8__2_chanx_right_out[6] ,
    \sb_1__8__2_chanx_right_out[7] ,
    \sb_1__8__2_chanx_right_out[8] ,
    \sb_1__8__2_chanx_right_out[9] ,
    \sb_1__8__2_chanx_right_out[10] ,
    \sb_1__8__2_chanx_right_out[11] ,
    \sb_1__8__2_chanx_right_out[12] ,
    \sb_1__8__2_chanx_right_out[13] ,
    \sb_1__8__2_chanx_right_out[14] ,
    \sb_1__8__2_chanx_right_out[15] ,
    \sb_1__8__2_chanx_right_out[16] ,
    \sb_1__8__2_chanx_right_out[17] ,
    \sb_1__8__2_chanx_right_out[18] ,
    \sb_1__8__2_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__3_chanx_left_out[0] ,
    \cbx_1__8__3_chanx_left_out[1] ,
    \cbx_1__8__3_chanx_left_out[2] ,
    \cbx_1__8__3_chanx_left_out[3] ,
    \cbx_1__8__3_chanx_left_out[4] ,
    \cbx_1__8__3_chanx_left_out[5] ,
    \cbx_1__8__3_chanx_left_out[6] ,
    \cbx_1__8__3_chanx_left_out[7] ,
    \cbx_1__8__3_chanx_left_out[8] ,
    \cbx_1__8__3_chanx_left_out[9] ,
    \cbx_1__8__3_chanx_left_out[10] ,
    \cbx_1__8__3_chanx_left_out[11] ,
    \cbx_1__8__3_chanx_left_out[12] ,
    \cbx_1__8__3_chanx_left_out[13] ,
    \cbx_1__8__3_chanx_left_out[14] ,
    \cbx_1__8__3_chanx_left_out[15] ,
    \cbx_1__8__3_chanx_left_out[16] ,
    \cbx_1__8__3_chanx_left_out[17] ,
    \cbx_1__8__3_chanx_left_out[18] ,
    \cbx_1__8__3_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__8__3_chanx_left_out[0] ,
    \sb_1__8__3_chanx_left_out[1] ,
    \sb_1__8__3_chanx_left_out[2] ,
    \sb_1__8__3_chanx_left_out[3] ,
    \sb_1__8__3_chanx_left_out[4] ,
    \sb_1__8__3_chanx_left_out[5] ,
    \sb_1__8__3_chanx_left_out[6] ,
    \sb_1__8__3_chanx_left_out[7] ,
    \sb_1__8__3_chanx_left_out[8] ,
    \sb_1__8__3_chanx_left_out[9] ,
    \sb_1__8__3_chanx_left_out[10] ,
    \sb_1__8__3_chanx_left_out[11] ,
    \sb_1__8__3_chanx_left_out[12] ,
    \sb_1__8__3_chanx_left_out[13] ,
    \sb_1__8__3_chanx_left_out[14] ,
    \sb_1__8__3_chanx_left_out[15] ,
    \sb_1__8__3_chanx_left_out[16] ,
    \sb_1__8__3_chanx_left_out[17] ,
    \sb_1__8__3_chanx_left_out[18] ,
    \sb_1__8__3_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__3_chanx_right_out[0] ,
    \cbx_1__8__3_chanx_right_out[1] ,
    \cbx_1__8__3_chanx_right_out[2] ,
    \cbx_1__8__3_chanx_right_out[3] ,
    \cbx_1__8__3_chanx_right_out[4] ,
    \cbx_1__8__3_chanx_right_out[5] ,
    \cbx_1__8__3_chanx_right_out[6] ,
    \cbx_1__8__3_chanx_right_out[7] ,
    \cbx_1__8__3_chanx_right_out[8] ,
    \cbx_1__8__3_chanx_right_out[9] ,
    \cbx_1__8__3_chanx_right_out[10] ,
    \cbx_1__8__3_chanx_right_out[11] ,
    \cbx_1__8__3_chanx_right_out[12] ,
    \cbx_1__8__3_chanx_right_out[13] ,
    \cbx_1__8__3_chanx_right_out[14] ,
    \cbx_1__8__3_chanx_right_out[15] ,
    \cbx_1__8__3_chanx_right_out[16] ,
    \cbx_1__8__3_chanx_right_out[17] ,
    \cbx_1__8__3_chanx_right_out[18] ,
    \cbx_1__8__3_chanx_right_out[19] }));
 cbx_1__0_ cbx_5__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[91] ),
    .SC_OUT_BOT(\scff_Wires[92] ),
    .bottom_grid_pin_0_(cbx_1__0__4_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__4_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__4_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__4_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__4_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__4_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__4_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__4_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__4_bottom_grid_pin_8_),
    .ccff_head(sb_1__0__4_ccff_tail),
    .ccff_tail(grid_io_bottom_3_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[121] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__4_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__4_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_3_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_3_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__4_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_3_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_3_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__4_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_3_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_3_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__4_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_3_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_3_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_3_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_3_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__4_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_3_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_3_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__4_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_3_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_3_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__4_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_3_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_3_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__4_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_3_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_3_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__0__3_chanx_right_out[0] ,
    \sb_1__0__3_chanx_right_out[1] ,
    \sb_1__0__3_chanx_right_out[2] ,
    \sb_1__0__3_chanx_right_out[3] ,
    \sb_1__0__3_chanx_right_out[4] ,
    \sb_1__0__3_chanx_right_out[5] ,
    \sb_1__0__3_chanx_right_out[6] ,
    \sb_1__0__3_chanx_right_out[7] ,
    \sb_1__0__3_chanx_right_out[8] ,
    \sb_1__0__3_chanx_right_out[9] ,
    \sb_1__0__3_chanx_right_out[10] ,
    \sb_1__0__3_chanx_right_out[11] ,
    \sb_1__0__3_chanx_right_out[12] ,
    \sb_1__0__3_chanx_right_out[13] ,
    \sb_1__0__3_chanx_right_out[14] ,
    \sb_1__0__3_chanx_right_out[15] ,
    \sb_1__0__3_chanx_right_out[16] ,
    \sb_1__0__3_chanx_right_out[17] ,
    \sb_1__0__3_chanx_right_out[18] ,
    \sb_1__0__3_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__4_chanx_left_out[0] ,
    \cbx_1__0__4_chanx_left_out[1] ,
    \cbx_1__0__4_chanx_left_out[2] ,
    \cbx_1__0__4_chanx_left_out[3] ,
    \cbx_1__0__4_chanx_left_out[4] ,
    \cbx_1__0__4_chanx_left_out[5] ,
    \cbx_1__0__4_chanx_left_out[6] ,
    \cbx_1__0__4_chanx_left_out[7] ,
    \cbx_1__0__4_chanx_left_out[8] ,
    \cbx_1__0__4_chanx_left_out[9] ,
    \cbx_1__0__4_chanx_left_out[10] ,
    \cbx_1__0__4_chanx_left_out[11] ,
    \cbx_1__0__4_chanx_left_out[12] ,
    \cbx_1__0__4_chanx_left_out[13] ,
    \cbx_1__0__4_chanx_left_out[14] ,
    \cbx_1__0__4_chanx_left_out[15] ,
    \cbx_1__0__4_chanx_left_out[16] ,
    \cbx_1__0__4_chanx_left_out[17] ,
    \cbx_1__0__4_chanx_left_out[18] ,
    \cbx_1__0__4_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__0__4_chanx_left_out[0] ,
    \sb_1__0__4_chanx_left_out[1] ,
    \sb_1__0__4_chanx_left_out[2] ,
    \sb_1__0__4_chanx_left_out[3] ,
    \sb_1__0__4_chanx_left_out[4] ,
    \sb_1__0__4_chanx_left_out[5] ,
    \sb_1__0__4_chanx_left_out[6] ,
    \sb_1__0__4_chanx_left_out[7] ,
    \sb_1__0__4_chanx_left_out[8] ,
    \sb_1__0__4_chanx_left_out[9] ,
    \sb_1__0__4_chanx_left_out[10] ,
    \sb_1__0__4_chanx_left_out[11] ,
    \sb_1__0__4_chanx_left_out[12] ,
    \sb_1__0__4_chanx_left_out[13] ,
    \sb_1__0__4_chanx_left_out[14] ,
    \sb_1__0__4_chanx_left_out[15] ,
    \sb_1__0__4_chanx_left_out[16] ,
    \sb_1__0__4_chanx_left_out[17] ,
    \sb_1__0__4_chanx_left_out[18] ,
    \sb_1__0__4_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__4_chanx_right_out[0] ,
    \cbx_1__0__4_chanx_right_out[1] ,
    \cbx_1__0__4_chanx_right_out[2] ,
    \cbx_1__0__4_chanx_right_out[3] ,
    \cbx_1__0__4_chanx_right_out[4] ,
    \cbx_1__0__4_chanx_right_out[5] ,
    \cbx_1__0__4_chanx_right_out[6] ,
    \cbx_1__0__4_chanx_right_out[7] ,
    \cbx_1__0__4_chanx_right_out[8] ,
    \cbx_1__0__4_chanx_right_out[9] ,
    \cbx_1__0__4_chanx_right_out[10] ,
    \cbx_1__0__4_chanx_right_out[11] ,
    \cbx_1__0__4_chanx_right_out[12] ,
    \cbx_1__0__4_chanx_right_out[13] ,
    \cbx_1__0__4_chanx_right_out[14] ,
    \cbx_1__0__4_chanx_right_out[15] ,
    \cbx_1__0__4_chanx_right_out[16] ,
    \cbx_1__0__4_chanx_right_out[17] ,
    \cbx_1__0__4_chanx_right_out[18] ,
    \cbx_1__0__4_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]}));
 cbx_1__1_ cbx_5__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[28] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[28] ),
    .SC_IN_TOP(\scff_Wires[88] ),
    .SC_OUT_BOT(\scff_Wires[89] ),
    .bottom_grid_pin_0_(cbx_1__1__28_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__28_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__28_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__28_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__28_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__28_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__28_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__28_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__28_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__28_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__28_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__28_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__28_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__28_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__28_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__28_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__28_ccff_tail),
    .ccff_tail(cbx_1__1__28_ccff_tail),
    .clk_1_N_out(\clk_1_wires[59] ),
    .clk_1_S_out(\clk_1_wires[60] ),
    .clk_1_W_in(\clk_1_wires[58] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[124] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[59] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[60] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[58] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__21_chanx_right_out[0] ,
    \sb_1__1__21_chanx_right_out[1] ,
    \sb_1__1__21_chanx_right_out[2] ,
    \sb_1__1__21_chanx_right_out[3] ,
    \sb_1__1__21_chanx_right_out[4] ,
    \sb_1__1__21_chanx_right_out[5] ,
    \sb_1__1__21_chanx_right_out[6] ,
    \sb_1__1__21_chanx_right_out[7] ,
    \sb_1__1__21_chanx_right_out[8] ,
    \sb_1__1__21_chanx_right_out[9] ,
    \sb_1__1__21_chanx_right_out[10] ,
    \sb_1__1__21_chanx_right_out[11] ,
    \sb_1__1__21_chanx_right_out[12] ,
    \sb_1__1__21_chanx_right_out[13] ,
    \sb_1__1__21_chanx_right_out[14] ,
    \sb_1__1__21_chanx_right_out[15] ,
    \sb_1__1__21_chanx_right_out[16] ,
    \sb_1__1__21_chanx_right_out[17] ,
    \sb_1__1__21_chanx_right_out[18] ,
    \sb_1__1__21_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__28_chanx_left_out[0] ,
    \cbx_1__1__28_chanx_left_out[1] ,
    \cbx_1__1__28_chanx_left_out[2] ,
    \cbx_1__1__28_chanx_left_out[3] ,
    \cbx_1__1__28_chanx_left_out[4] ,
    \cbx_1__1__28_chanx_left_out[5] ,
    \cbx_1__1__28_chanx_left_out[6] ,
    \cbx_1__1__28_chanx_left_out[7] ,
    \cbx_1__1__28_chanx_left_out[8] ,
    \cbx_1__1__28_chanx_left_out[9] ,
    \cbx_1__1__28_chanx_left_out[10] ,
    \cbx_1__1__28_chanx_left_out[11] ,
    \cbx_1__1__28_chanx_left_out[12] ,
    \cbx_1__1__28_chanx_left_out[13] ,
    \cbx_1__1__28_chanx_left_out[14] ,
    \cbx_1__1__28_chanx_left_out[15] ,
    \cbx_1__1__28_chanx_left_out[16] ,
    \cbx_1__1__28_chanx_left_out[17] ,
    \cbx_1__1__28_chanx_left_out[18] ,
    \cbx_1__1__28_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__28_chanx_left_out[0] ,
    \sb_1__1__28_chanx_left_out[1] ,
    \sb_1__1__28_chanx_left_out[2] ,
    \sb_1__1__28_chanx_left_out[3] ,
    \sb_1__1__28_chanx_left_out[4] ,
    \sb_1__1__28_chanx_left_out[5] ,
    \sb_1__1__28_chanx_left_out[6] ,
    \sb_1__1__28_chanx_left_out[7] ,
    \sb_1__1__28_chanx_left_out[8] ,
    \sb_1__1__28_chanx_left_out[9] ,
    \sb_1__1__28_chanx_left_out[10] ,
    \sb_1__1__28_chanx_left_out[11] ,
    \sb_1__1__28_chanx_left_out[12] ,
    \sb_1__1__28_chanx_left_out[13] ,
    \sb_1__1__28_chanx_left_out[14] ,
    \sb_1__1__28_chanx_left_out[15] ,
    \sb_1__1__28_chanx_left_out[16] ,
    \sb_1__1__28_chanx_left_out[17] ,
    \sb_1__1__28_chanx_left_out[18] ,
    \sb_1__1__28_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__28_chanx_right_out[0] ,
    \cbx_1__1__28_chanx_right_out[1] ,
    \cbx_1__1__28_chanx_right_out[2] ,
    \cbx_1__1__28_chanx_right_out[3] ,
    \cbx_1__1__28_chanx_right_out[4] ,
    \cbx_1__1__28_chanx_right_out[5] ,
    \cbx_1__1__28_chanx_right_out[6] ,
    \cbx_1__1__28_chanx_right_out[7] ,
    \cbx_1__1__28_chanx_right_out[8] ,
    \cbx_1__1__28_chanx_right_out[9] ,
    \cbx_1__1__28_chanx_right_out[10] ,
    \cbx_1__1__28_chanx_right_out[11] ,
    \cbx_1__1__28_chanx_right_out[12] ,
    \cbx_1__1__28_chanx_right_out[13] ,
    \cbx_1__1__28_chanx_right_out[14] ,
    \cbx_1__1__28_chanx_right_out[15] ,
    \cbx_1__1__28_chanx_right_out[16] ,
    \cbx_1__1__28_chanx_right_out[17] ,
    \cbx_1__1__28_chanx_right_out[18] ,
    \cbx_1__1__28_chanx_right_out[19] }));
 cbx_1__1_ cbx_5__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[29] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[29] ),
    .SC_IN_TOP(\scff_Wires[86] ),
    .SC_OUT_BOT(\scff_Wires[87] ),
    .bottom_grid_pin_0_(cbx_1__1__29_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__29_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__29_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__29_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__29_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__29_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__29_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__29_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__29_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__29_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__29_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__29_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__29_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__29_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__29_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__29_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__29_ccff_tail),
    .ccff_tail(cbx_1__1__29_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[127] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__22_chanx_right_out[0] ,
    \sb_1__1__22_chanx_right_out[1] ,
    \sb_1__1__22_chanx_right_out[2] ,
    \sb_1__1__22_chanx_right_out[3] ,
    \sb_1__1__22_chanx_right_out[4] ,
    \sb_1__1__22_chanx_right_out[5] ,
    \sb_1__1__22_chanx_right_out[6] ,
    \sb_1__1__22_chanx_right_out[7] ,
    \sb_1__1__22_chanx_right_out[8] ,
    \sb_1__1__22_chanx_right_out[9] ,
    \sb_1__1__22_chanx_right_out[10] ,
    \sb_1__1__22_chanx_right_out[11] ,
    \sb_1__1__22_chanx_right_out[12] ,
    \sb_1__1__22_chanx_right_out[13] ,
    \sb_1__1__22_chanx_right_out[14] ,
    \sb_1__1__22_chanx_right_out[15] ,
    \sb_1__1__22_chanx_right_out[16] ,
    \sb_1__1__22_chanx_right_out[17] ,
    \sb_1__1__22_chanx_right_out[18] ,
    \sb_1__1__22_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__29_chanx_left_out[0] ,
    \cbx_1__1__29_chanx_left_out[1] ,
    \cbx_1__1__29_chanx_left_out[2] ,
    \cbx_1__1__29_chanx_left_out[3] ,
    \cbx_1__1__29_chanx_left_out[4] ,
    \cbx_1__1__29_chanx_left_out[5] ,
    \cbx_1__1__29_chanx_left_out[6] ,
    \cbx_1__1__29_chanx_left_out[7] ,
    \cbx_1__1__29_chanx_left_out[8] ,
    \cbx_1__1__29_chanx_left_out[9] ,
    \cbx_1__1__29_chanx_left_out[10] ,
    \cbx_1__1__29_chanx_left_out[11] ,
    \cbx_1__1__29_chanx_left_out[12] ,
    \cbx_1__1__29_chanx_left_out[13] ,
    \cbx_1__1__29_chanx_left_out[14] ,
    \cbx_1__1__29_chanx_left_out[15] ,
    \cbx_1__1__29_chanx_left_out[16] ,
    \cbx_1__1__29_chanx_left_out[17] ,
    \cbx_1__1__29_chanx_left_out[18] ,
    \cbx_1__1__29_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__29_chanx_left_out[0] ,
    \sb_1__1__29_chanx_left_out[1] ,
    \sb_1__1__29_chanx_left_out[2] ,
    \sb_1__1__29_chanx_left_out[3] ,
    \sb_1__1__29_chanx_left_out[4] ,
    \sb_1__1__29_chanx_left_out[5] ,
    \sb_1__1__29_chanx_left_out[6] ,
    \sb_1__1__29_chanx_left_out[7] ,
    \sb_1__1__29_chanx_left_out[8] ,
    \sb_1__1__29_chanx_left_out[9] ,
    \sb_1__1__29_chanx_left_out[10] ,
    \sb_1__1__29_chanx_left_out[11] ,
    \sb_1__1__29_chanx_left_out[12] ,
    \sb_1__1__29_chanx_left_out[13] ,
    \sb_1__1__29_chanx_left_out[14] ,
    \sb_1__1__29_chanx_left_out[15] ,
    \sb_1__1__29_chanx_left_out[16] ,
    \sb_1__1__29_chanx_left_out[17] ,
    \sb_1__1__29_chanx_left_out[18] ,
    \sb_1__1__29_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__29_chanx_right_out[0] ,
    \cbx_1__1__29_chanx_right_out[1] ,
    \cbx_1__1__29_chanx_right_out[2] ,
    \cbx_1__1__29_chanx_right_out[3] ,
    \cbx_1__1__29_chanx_right_out[4] ,
    \cbx_1__1__29_chanx_right_out[5] ,
    \cbx_1__1__29_chanx_right_out[6] ,
    \cbx_1__1__29_chanx_right_out[7] ,
    \cbx_1__1__29_chanx_right_out[8] ,
    \cbx_1__1__29_chanx_right_out[9] ,
    \cbx_1__1__29_chanx_right_out[10] ,
    \cbx_1__1__29_chanx_right_out[11] ,
    \cbx_1__1__29_chanx_right_out[12] ,
    \cbx_1__1__29_chanx_right_out[13] ,
    \cbx_1__1__29_chanx_right_out[14] ,
    \cbx_1__1__29_chanx_right_out[15] ,
    \cbx_1__1__29_chanx_right_out[16] ,
    \cbx_1__1__29_chanx_right_out[17] ,
    \cbx_1__1__29_chanx_right_out[18] ,
    \cbx_1__1__29_chanx_right_out[19] }));
 cbx_1__1_ cbx_5__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[30] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[30] ),
    .SC_IN_TOP(\scff_Wires[84] ),
    .SC_OUT_BOT(\scff_Wires[85] ),
    .bottom_grid_pin_0_(cbx_1__1__30_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__30_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__30_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__30_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__30_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__30_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__30_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__30_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__30_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__30_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__30_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__30_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__30_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__30_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__30_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__30_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__30_ccff_tail),
    .ccff_tail(cbx_1__1__30_ccff_tail),
    .clk_1_N_out(\clk_1_wires[66] ),
    .clk_1_S_out(\clk_1_wires[67] ),
    .clk_1_W_in(\clk_1_wires[65] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[130] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[66] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[67] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[65] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__23_chanx_right_out[0] ,
    \sb_1__1__23_chanx_right_out[1] ,
    \sb_1__1__23_chanx_right_out[2] ,
    \sb_1__1__23_chanx_right_out[3] ,
    \sb_1__1__23_chanx_right_out[4] ,
    \sb_1__1__23_chanx_right_out[5] ,
    \sb_1__1__23_chanx_right_out[6] ,
    \sb_1__1__23_chanx_right_out[7] ,
    \sb_1__1__23_chanx_right_out[8] ,
    \sb_1__1__23_chanx_right_out[9] ,
    \sb_1__1__23_chanx_right_out[10] ,
    \sb_1__1__23_chanx_right_out[11] ,
    \sb_1__1__23_chanx_right_out[12] ,
    \sb_1__1__23_chanx_right_out[13] ,
    \sb_1__1__23_chanx_right_out[14] ,
    \sb_1__1__23_chanx_right_out[15] ,
    \sb_1__1__23_chanx_right_out[16] ,
    \sb_1__1__23_chanx_right_out[17] ,
    \sb_1__1__23_chanx_right_out[18] ,
    \sb_1__1__23_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__30_chanx_left_out[0] ,
    \cbx_1__1__30_chanx_left_out[1] ,
    \cbx_1__1__30_chanx_left_out[2] ,
    \cbx_1__1__30_chanx_left_out[3] ,
    \cbx_1__1__30_chanx_left_out[4] ,
    \cbx_1__1__30_chanx_left_out[5] ,
    \cbx_1__1__30_chanx_left_out[6] ,
    \cbx_1__1__30_chanx_left_out[7] ,
    \cbx_1__1__30_chanx_left_out[8] ,
    \cbx_1__1__30_chanx_left_out[9] ,
    \cbx_1__1__30_chanx_left_out[10] ,
    \cbx_1__1__30_chanx_left_out[11] ,
    \cbx_1__1__30_chanx_left_out[12] ,
    \cbx_1__1__30_chanx_left_out[13] ,
    \cbx_1__1__30_chanx_left_out[14] ,
    \cbx_1__1__30_chanx_left_out[15] ,
    \cbx_1__1__30_chanx_left_out[16] ,
    \cbx_1__1__30_chanx_left_out[17] ,
    \cbx_1__1__30_chanx_left_out[18] ,
    \cbx_1__1__30_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__30_chanx_left_out[0] ,
    \sb_1__1__30_chanx_left_out[1] ,
    \sb_1__1__30_chanx_left_out[2] ,
    \sb_1__1__30_chanx_left_out[3] ,
    \sb_1__1__30_chanx_left_out[4] ,
    \sb_1__1__30_chanx_left_out[5] ,
    \sb_1__1__30_chanx_left_out[6] ,
    \sb_1__1__30_chanx_left_out[7] ,
    \sb_1__1__30_chanx_left_out[8] ,
    \sb_1__1__30_chanx_left_out[9] ,
    \sb_1__1__30_chanx_left_out[10] ,
    \sb_1__1__30_chanx_left_out[11] ,
    \sb_1__1__30_chanx_left_out[12] ,
    \sb_1__1__30_chanx_left_out[13] ,
    \sb_1__1__30_chanx_left_out[14] ,
    \sb_1__1__30_chanx_left_out[15] ,
    \sb_1__1__30_chanx_left_out[16] ,
    \sb_1__1__30_chanx_left_out[17] ,
    \sb_1__1__30_chanx_left_out[18] ,
    \sb_1__1__30_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__30_chanx_right_out[0] ,
    \cbx_1__1__30_chanx_right_out[1] ,
    \cbx_1__1__30_chanx_right_out[2] ,
    \cbx_1__1__30_chanx_right_out[3] ,
    \cbx_1__1__30_chanx_right_out[4] ,
    \cbx_1__1__30_chanx_right_out[5] ,
    \cbx_1__1__30_chanx_right_out[6] ,
    \cbx_1__1__30_chanx_right_out[7] ,
    \cbx_1__1__30_chanx_right_out[8] ,
    \cbx_1__1__30_chanx_right_out[9] ,
    \cbx_1__1__30_chanx_right_out[10] ,
    \cbx_1__1__30_chanx_right_out[11] ,
    \cbx_1__1__30_chanx_right_out[12] ,
    \cbx_1__1__30_chanx_right_out[13] ,
    \cbx_1__1__30_chanx_right_out[14] ,
    \cbx_1__1__30_chanx_right_out[15] ,
    \cbx_1__1__30_chanx_right_out[16] ,
    \cbx_1__1__30_chanx_right_out[17] ,
    \cbx_1__1__30_chanx_right_out[18] ,
    \cbx_1__1__30_chanx_right_out[19] }));
 cbx_1__1_ cbx_5__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[31] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[31] ),
    .SC_IN_TOP(\scff_Wires[82] ),
    .SC_OUT_BOT(\scff_Wires[83] ),
    .bottom_grid_pin_0_(cbx_1__1__31_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__31_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__31_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__31_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__31_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__31_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__31_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__31_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__31_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__31_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__31_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__31_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__31_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__31_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__31_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__31_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__31_ccff_tail),
    .ccff_tail(cbx_1__1__31_ccff_tail),
    .clk_3_E_out(\clk_3_wires[2] ),
    .clk_3_W_in(\clk_3_wires[1] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[133] ),
    .prog_clk_3_E_out(\prog_clk_3_wires[2] ),
    .prog_clk_3_W_in(\prog_clk_3_wires[1] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__24_chanx_right_out[0] ,
    \sb_1__1__24_chanx_right_out[1] ,
    \sb_1__1__24_chanx_right_out[2] ,
    \sb_1__1__24_chanx_right_out[3] ,
    \sb_1__1__24_chanx_right_out[4] ,
    \sb_1__1__24_chanx_right_out[5] ,
    \sb_1__1__24_chanx_right_out[6] ,
    \sb_1__1__24_chanx_right_out[7] ,
    \sb_1__1__24_chanx_right_out[8] ,
    \sb_1__1__24_chanx_right_out[9] ,
    \sb_1__1__24_chanx_right_out[10] ,
    \sb_1__1__24_chanx_right_out[11] ,
    \sb_1__1__24_chanx_right_out[12] ,
    \sb_1__1__24_chanx_right_out[13] ,
    \sb_1__1__24_chanx_right_out[14] ,
    \sb_1__1__24_chanx_right_out[15] ,
    \sb_1__1__24_chanx_right_out[16] ,
    \sb_1__1__24_chanx_right_out[17] ,
    \sb_1__1__24_chanx_right_out[18] ,
    \sb_1__1__24_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__31_chanx_left_out[0] ,
    \cbx_1__1__31_chanx_left_out[1] ,
    \cbx_1__1__31_chanx_left_out[2] ,
    \cbx_1__1__31_chanx_left_out[3] ,
    \cbx_1__1__31_chanx_left_out[4] ,
    \cbx_1__1__31_chanx_left_out[5] ,
    \cbx_1__1__31_chanx_left_out[6] ,
    \cbx_1__1__31_chanx_left_out[7] ,
    \cbx_1__1__31_chanx_left_out[8] ,
    \cbx_1__1__31_chanx_left_out[9] ,
    \cbx_1__1__31_chanx_left_out[10] ,
    \cbx_1__1__31_chanx_left_out[11] ,
    \cbx_1__1__31_chanx_left_out[12] ,
    \cbx_1__1__31_chanx_left_out[13] ,
    \cbx_1__1__31_chanx_left_out[14] ,
    \cbx_1__1__31_chanx_left_out[15] ,
    \cbx_1__1__31_chanx_left_out[16] ,
    \cbx_1__1__31_chanx_left_out[17] ,
    \cbx_1__1__31_chanx_left_out[18] ,
    \cbx_1__1__31_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__31_chanx_left_out[0] ,
    \sb_1__1__31_chanx_left_out[1] ,
    \sb_1__1__31_chanx_left_out[2] ,
    \sb_1__1__31_chanx_left_out[3] ,
    \sb_1__1__31_chanx_left_out[4] ,
    \sb_1__1__31_chanx_left_out[5] ,
    \sb_1__1__31_chanx_left_out[6] ,
    \sb_1__1__31_chanx_left_out[7] ,
    \sb_1__1__31_chanx_left_out[8] ,
    \sb_1__1__31_chanx_left_out[9] ,
    \sb_1__1__31_chanx_left_out[10] ,
    \sb_1__1__31_chanx_left_out[11] ,
    \sb_1__1__31_chanx_left_out[12] ,
    \sb_1__1__31_chanx_left_out[13] ,
    \sb_1__1__31_chanx_left_out[14] ,
    \sb_1__1__31_chanx_left_out[15] ,
    \sb_1__1__31_chanx_left_out[16] ,
    \sb_1__1__31_chanx_left_out[17] ,
    \sb_1__1__31_chanx_left_out[18] ,
    \sb_1__1__31_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__31_chanx_right_out[0] ,
    \cbx_1__1__31_chanx_right_out[1] ,
    \cbx_1__1__31_chanx_right_out[2] ,
    \cbx_1__1__31_chanx_right_out[3] ,
    \cbx_1__1__31_chanx_right_out[4] ,
    \cbx_1__1__31_chanx_right_out[5] ,
    \cbx_1__1__31_chanx_right_out[6] ,
    \cbx_1__1__31_chanx_right_out[7] ,
    \cbx_1__1__31_chanx_right_out[8] ,
    \cbx_1__1__31_chanx_right_out[9] ,
    \cbx_1__1__31_chanx_right_out[10] ,
    \cbx_1__1__31_chanx_right_out[11] ,
    \cbx_1__1__31_chanx_right_out[12] ,
    \cbx_1__1__31_chanx_right_out[13] ,
    \cbx_1__1__31_chanx_right_out[14] ,
    \cbx_1__1__31_chanx_right_out[15] ,
    \cbx_1__1__31_chanx_right_out[16] ,
    \cbx_1__1__31_chanx_right_out[17] ,
    \cbx_1__1__31_chanx_right_out[18] ,
    \cbx_1__1__31_chanx_right_out[19] }));
 cbx_1__1_ cbx_5__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[32] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[32] ),
    .SC_IN_TOP(\scff_Wires[80] ),
    .SC_OUT_BOT(\scff_Wires[81] ),
    .bottom_grid_pin_0_(cbx_1__1__32_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__32_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__32_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__32_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__32_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__32_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__32_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__32_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__32_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__32_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__32_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__32_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__32_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__32_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__32_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__32_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__32_ccff_tail),
    .ccff_tail(cbx_1__1__32_ccff_tail),
    .clk_1_N_out(\clk_1_wires[73] ),
    .clk_1_S_out(\clk_1_wires[74] ),
    .clk_1_W_in(\clk_1_wires[72] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[136] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[73] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[74] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[72] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__25_chanx_right_out[0] ,
    \sb_1__1__25_chanx_right_out[1] ,
    \sb_1__1__25_chanx_right_out[2] ,
    \sb_1__1__25_chanx_right_out[3] ,
    \sb_1__1__25_chanx_right_out[4] ,
    \sb_1__1__25_chanx_right_out[5] ,
    \sb_1__1__25_chanx_right_out[6] ,
    \sb_1__1__25_chanx_right_out[7] ,
    \sb_1__1__25_chanx_right_out[8] ,
    \sb_1__1__25_chanx_right_out[9] ,
    \sb_1__1__25_chanx_right_out[10] ,
    \sb_1__1__25_chanx_right_out[11] ,
    \sb_1__1__25_chanx_right_out[12] ,
    \sb_1__1__25_chanx_right_out[13] ,
    \sb_1__1__25_chanx_right_out[14] ,
    \sb_1__1__25_chanx_right_out[15] ,
    \sb_1__1__25_chanx_right_out[16] ,
    \sb_1__1__25_chanx_right_out[17] ,
    \sb_1__1__25_chanx_right_out[18] ,
    \sb_1__1__25_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__32_chanx_left_out[0] ,
    \cbx_1__1__32_chanx_left_out[1] ,
    \cbx_1__1__32_chanx_left_out[2] ,
    \cbx_1__1__32_chanx_left_out[3] ,
    \cbx_1__1__32_chanx_left_out[4] ,
    \cbx_1__1__32_chanx_left_out[5] ,
    \cbx_1__1__32_chanx_left_out[6] ,
    \cbx_1__1__32_chanx_left_out[7] ,
    \cbx_1__1__32_chanx_left_out[8] ,
    \cbx_1__1__32_chanx_left_out[9] ,
    \cbx_1__1__32_chanx_left_out[10] ,
    \cbx_1__1__32_chanx_left_out[11] ,
    \cbx_1__1__32_chanx_left_out[12] ,
    \cbx_1__1__32_chanx_left_out[13] ,
    \cbx_1__1__32_chanx_left_out[14] ,
    \cbx_1__1__32_chanx_left_out[15] ,
    \cbx_1__1__32_chanx_left_out[16] ,
    \cbx_1__1__32_chanx_left_out[17] ,
    \cbx_1__1__32_chanx_left_out[18] ,
    \cbx_1__1__32_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__32_chanx_left_out[0] ,
    \sb_1__1__32_chanx_left_out[1] ,
    \sb_1__1__32_chanx_left_out[2] ,
    \sb_1__1__32_chanx_left_out[3] ,
    \sb_1__1__32_chanx_left_out[4] ,
    \sb_1__1__32_chanx_left_out[5] ,
    \sb_1__1__32_chanx_left_out[6] ,
    \sb_1__1__32_chanx_left_out[7] ,
    \sb_1__1__32_chanx_left_out[8] ,
    \sb_1__1__32_chanx_left_out[9] ,
    \sb_1__1__32_chanx_left_out[10] ,
    \sb_1__1__32_chanx_left_out[11] ,
    \sb_1__1__32_chanx_left_out[12] ,
    \sb_1__1__32_chanx_left_out[13] ,
    \sb_1__1__32_chanx_left_out[14] ,
    \sb_1__1__32_chanx_left_out[15] ,
    \sb_1__1__32_chanx_left_out[16] ,
    \sb_1__1__32_chanx_left_out[17] ,
    \sb_1__1__32_chanx_left_out[18] ,
    \sb_1__1__32_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__32_chanx_right_out[0] ,
    \cbx_1__1__32_chanx_right_out[1] ,
    \cbx_1__1__32_chanx_right_out[2] ,
    \cbx_1__1__32_chanx_right_out[3] ,
    \cbx_1__1__32_chanx_right_out[4] ,
    \cbx_1__1__32_chanx_right_out[5] ,
    \cbx_1__1__32_chanx_right_out[6] ,
    \cbx_1__1__32_chanx_right_out[7] ,
    \cbx_1__1__32_chanx_right_out[8] ,
    \cbx_1__1__32_chanx_right_out[9] ,
    \cbx_1__1__32_chanx_right_out[10] ,
    \cbx_1__1__32_chanx_right_out[11] ,
    \cbx_1__1__32_chanx_right_out[12] ,
    \cbx_1__1__32_chanx_right_out[13] ,
    \cbx_1__1__32_chanx_right_out[14] ,
    \cbx_1__1__32_chanx_right_out[15] ,
    \cbx_1__1__32_chanx_right_out[16] ,
    \cbx_1__1__32_chanx_right_out[17] ,
    \cbx_1__1__32_chanx_right_out[18] ,
    \cbx_1__1__32_chanx_right_out[19] }));
 cbx_1__1_ cbx_5__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[33] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[33] ),
    .SC_IN_TOP(\scff_Wires[78] ),
    .SC_OUT_BOT(\scff_Wires[79] ),
    .bottom_grid_pin_0_(cbx_1__1__33_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__33_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__33_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__33_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__33_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__33_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__33_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__33_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__33_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__33_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__33_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__33_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__33_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__33_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__33_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__33_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__33_ccff_tail),
    .ccff_tail(cbx_1__1__33_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[139] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__26_chanx_right_out[0] ,
    \sb_1__1__26_chanx_right_out[1] ,
    \sb_1__1__26_chanx_right_out[2] ,
    \sb_1__1__26_chanx_right_out[3] ,
    \sb_1__1__26_chanx_right_out[4] ,
    \sb_1__1__26_chanx_right_out[5] ,
    \sb_1__1__26_chanx_right_out[6] ,
    \sb_1__1__26_chanx_right_out[7] ,
    \sb_1__1__26_chanx_right_out[8] ,
    \sb_1__1__26_chanx_right_out[9] ,
    \sb_1__1__26_chanx_right_out[10] ,
    \sb_1__1__26_chanx_right_out[11] ,
    \sb_1__1__26_chanx_right_out[12] ,
    \sb_1__1__26_chanx_right_out[13] ,
    \sb_1__1__26_chanx_right_out[14] ,
    \sb_1__1__26_chanx_right_out[15] ,
    \sb_1__1__26_chanx_right_out[16] ,
    \sb_1__1__26_chanx_right_out[17] ,
    \sb_1__1__26_chanx_right_out[18] ,
    \sb_1__1__26_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__33_chanx_left_out[0] ,
    \cbx_1__1__33_chanx_left_out[1] ,
    \cbx_1__1__33_chanx_left_out[2] ,
    \cbx_1__1__33_chanx_left_out[3] ,
    \cbx_1__1__33_chanx_left_out[4] ,
    \cbx_1__1__33_chanx_left_out[5] ,
    \cbx_1__1__33_chanx_left_out[6] ,
    \cbx_1__1__33_chanx_left_out[7] ,
    \cbx_1__1__33_chanx_left_out[8] ,
    \cbx_1__1__33_chanx_left_out[9] ,
    \cbx_1__1__33_chanx_left_out[10] ,
    \cbx_1__1__33_chanx_left_out[11] ,
    \cbx_1__1__33_chanx_left_out[12] ,
    \cbx_1__1__33_chanx_left_out[13] ,
    \cbx_1__1__33_chanx_left_out[14] ,
    \cbx_1__1__33_chanx_left_out[15] ,
    \cbx_1__1__33_chanx_left_out[16] ,
    \cbx_1__1__33_chanx_left_out[17] ,
    \cbx_1__1__33_chanx_left_out[18] ,
    \cbx_1__1__33_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__33_chanx_left_out[0] ,
    \sb_1__1__33_chanx_left_out[1] ,
    \sb_1__1__33_chanx_left_out[2] ,
    \sb_1__1__33_chanx_left_out[3] ,
    \sb_1__1__33_chanx_left_out[4] ,
    \sb_1__1__33_chanx_left_out[5] ,
    \sb_1__1__33_chanx_left_out[6] ,
    \sb_1__1__33_chanx_left_out[7] ,
    \sb_1__1__33_chanx_left_out[8] ,
    \sb_1__1__33_chanx_left_out[9] ,
    \sb_1__1__33_chanx_left_out[10] ,
    \sb_1__1__33_chanx_left_out[11] ,
    \sb_1__1__33_chanx_left_out[12] ,
    \sb_1__1__33_chanx_left_out[13] ,
    \sb_1__1__33_chanx_left_out[14] ,
    \sb_1__1__33_chanx_left_out[15] ,
    \sb_1__1__33_chanx_left_out[16] ,
    \sb_1__1__33_chanx_left_out[17] ,
    \sb_1__1__33_chanx_left_out[18] ,
    \sb_1__1__33_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__33_chanx_right_out[0] ,
    \cbx_1__1__33_chanx_right_out[1] ,
    \cbx_1__1__33_chanx_right_out[2] ,
    \cbx_1__1__33_chanx_right_out[3] ,
    \cbx_1__1__33_chanx_right_out[4] ,
    \cbx_1__1__33_chanx_right_out[5] ,
    \cbx_1__1__33_chanx_right_out[6] ,
    \cbx_1__1__33_chanx_right_out[7] ,
    \cbx_1__1__33_chanx_right_out[8] ,
    \cbx_1__1__33_chanx_right_out[9] ,
    \cbx_1__1__33_chanx_right_out[10] ,
    \cbx_1__1__33_chanx_right_out[11] ,
    \cbx_1__1__33_chanx_right_out[12] ,
    \cbx_1__1__33_chanx_right_out[13] ,
    \cbx_1__1__33_chanx_right_out[14] ,
    \cbx_1__1__33_chanx_right_out[15] ,
    \cbx_1__1__33_chanx_right_out[16] ,
    \cbx_1__1__33_chanx_right_out[17] ,
    \cbx_1__1__33_chanx_right_out[18] ,
    \cbx_1__1__33_chanx_right_out[19] }));
 cbx_1__1_ cbx_5__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[34] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[34] ),
    .SC_IN_TOP(\scff_Wires[76] ),
    .SC_OUT_BOT(\scff_Wires[77] ),
    .bottom_grid_pin_0_(cbx_1__1__34_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__34_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__34_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__34_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__34_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__34_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__34_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__34_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__34_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__34_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__34_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__34_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__34_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__34_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__34_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__34_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__34_ccff_tail),
    .ccff_tail(cbx_1__1__34_ccff_tail),
    .clk_1_N_out(\clk_1_wires[80] ),
    .clk_1_S_out(\clk_1_wires[81] ),
    .clk_1_W_in(\clk_1_wires[79] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[142] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[80] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[81] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[79] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__27_chanx_right_out[0] ,
    \sb_1__1__27_chanx_right_out[1] ,
    \sb_1__1__27_chanx_right_out[2] ,
    \sb_1__1__27_chanx_right_out[3] ,
    \sb_1__1__27_chanx_right_out[4] ,
    \sb_1__1__27_chanx_right_out[5] ,
    \sb_1__1__27_chanx_right_out[6] ,
    \sb_1__1__27_chanx_right_out[7] ,
    \sb_1__1__27_chanx_right_out[8] ,
    \sb_1__1__27_chanx_right_out[9] ,
    \sb_1__1__27_chanx_right_out[10] ,
    \sb_1__1__27_chanx_right_out[11] ,
    \sb_1__1__27_chanx_right_out[12] ,
    \sb_1__1__27_chanx_right_out[13] ,
    \sb_1__1__27_chanx_right_out[14] ,
    \sb_1__1__27_chanx_right_out[15] ,
    \sb_1__1__27_chanx_right_out[16] ,
    \sb_1__1__27_chanx_right_out[17] ,
    \sb_1__1__27_chanx_right_out[18] ,
    \sb_1__1__27_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__34_chanx_left_out[0] ,
    \cbx_1__1__34_chanx_left_out[1] ,
    \cbx_1__1__34_chanx_left_out[2] ,
    \cbx_1__1__34_chanx_left_out[3] ,
    \cbx_1__1__34_chanx_left_out[4] ,
    \cbx_1__1__34_chanx_left_out[5] ,
    \cbx_1__1__34_chanx_left_out[6] ,
    \cbx_1__1__34_chanx_left_out[7] ,
    \cbx_1__1__34_chanx_left_out[8] ,
    \cbx_1__1__34_chanx_left_out[9] ,
    \cbx_1__1__34_chanx_left_out[10] ,
    \cbx_1__1__34_chanx_left_out[11] ,
    \cbx_1__1__34_chanx_left_out[12] ,
    \cbx_1__1__34_chanx_left_out[13] ,
    \cbx_1__1__34_chanx_left_out[14] ,
    \cbx_1__1__34_chanx_left_out[15] ,
    \cbx_1__1__34_chanx_left_out[16] ,
    \cbx_1__1__34_chanx_left_out[17] ,
    \cbx_1__1__34_chanx_left_out[18] ,
    \cbx_1__1__34_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__34_chanx_left_out[0] ,
    \sb_1__1__34_chanx_left_out[1] ,
    \sb_1__1__34_chanx_left_out[2] ,
    \sb_1__1__34_chanx_left_out[3] ,
    \sb_1__1__34_chanx_left_out[4] ,
    \sb_1__1__34_chanx_left_out[5] ,
    \sb_1__1__34_chanx_left_out[6] ,
    \sb_1__1__34_chanx_left_out[7] ,
    \sb_1__1__34_chanx_left_out[8] ,
    \sb_1__1__34_chanx_left_out[9] ,
    \sb_1__1__34_chanx_left_out[10] ,
    \sb_1__1__34_chanx_left_out[11] ,
    \sb_1__1__34_chanx_left_out[12] ,
    \sb_1__1__34_chanx_left_out[13] ,
    \sb_1__1__34_chanx_left_out[14] ,
    \sb_1__1__34_chanx_left_out[15] ,
    \sb_1__1__34_chanx_left_out[16] ,
    \sb_1__1__34_chanx_left_out[17] ,
    \sb_1__1__34_chanx_left_out[18] ,
    \sb_1__1__34_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__34_chanx_right_out[0] ,
    \cbx_1__1__34_chanx_right_out[1] ,
    \cbx_1__1__34_chanx_right_out[2] ,
    \cbx_1__1__34_chanx_right_out[3] ,
    \cbx_1__1__34_chanx_right_out[4] ,
    \cbx_1__1__34_chanx_right_out[5] ,
    \cbx_1__1__34_chanx_right_out[6] ,
    \cbx_1__1__34_chanx_right_out[7] ,
    \cbx_1__1__34_chanx_right_out[8] ,
    \cbx_1__1__34_chanx_right_out[9] ,
    \cbx_1__1__34_chanx_right_out[10] ,
    \cbx_1__1__34_chanx_right_out[11] ,
    \cbx_1__1__34_chanx_right_out[12] ,
    \cbx_1__1__34_chanx_right_out[13] ,
    \cbx_1__1__34_chanx_right_out[14] ,
    \cbx_1__1__34_chanx_right_out[15] ,
    \cbx_1__1__34_chanx_right_out[16] ,
    \cbx_1__1__34_chanx_right_out[17] ,
    \cbx_1__1__34_chanx_right_out[18] ,
    \cbx_1__1__34_chanx_right_out[19] }));
 cbx_1__2_ cbx_5__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[74] ),
    .SC_OUT_BOT(\scff_Wires[75] ),
    .bottom_grid_pin_0_(cbx_1__8__4_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__4_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__4_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__4_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__4_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__4_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__4_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__4_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__4_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__4_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__4_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__4_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__4_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__4_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__4_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__4_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__4_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_4_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_4_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_1__8__4_ccff_tail),
    .ccff_tail(grid_io_top_4_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]),
    .prog_clk_0_S_in(\prog_clk_0_wires[145] ),
    .top_grid_pin_0_(cbx_1__8__4_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__8__3_chanx_right_out[0] ,
    \sb_1__8__3_chanx_right_out[1] ,
    \sb_1__8__3_chanx_right_out[2] ,
    \sb_1__8__3_chanx_right_out[3] ,
    \sb_1__8__3_chanx_right_out[4] ,
    \sb_1__8__3_chanx_right_out[5] ,
    \sb_1__8__3_chanx_right_out[6] ,
    \sb_1__8__3_chanx_right_out[7] ,
    \sb_1__8__3_chanx_right_out[8] ,
    \sb_1__8__3_chanx_right_out[9] ,
    \sb_1__8__3_chanx_right_out[10] ,
    \sb_1__8__3_chanx_right_out[11] ,
    \sb_1__8__3_chanx_right_out[12] ,
    \sb_1__8__3_chanx_right_out[13] ,
    \sb_1__8__3_chanx_right_out[14] ,
    \sb_1__8__3_chanx_right_out[15] ,
    \sb_1__8__3_chanx_right_out[16] ,
    \sb_1__8__3_chanx_right_out[17] ,
    \sb_1__8__3_chanx_right_out[18] ,
    \sb_1__8__3_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__4_chanx_left_out[0] ,
    \cbx_1__8__4_chanx_left_out[1] ,
    \cbx_1__8__4_chanx_left_out[2] ,
    \cbx_1__8__4_chanx_left_out[3] ,
    \cbx_1__8__4_chanx_left_out[4] ,
    \cbx_1__8__4_chanx_left_out[5] ,
    \cbx_1__8__4_chanx_left_out[6] ,
    \cbx_1__8__4_chanx_left_out[7] ,
    \cbx_1__8__4_chanx_left_out[8] ,
    \cbx_1__8__4_chanx_left_out[9] ,
    \cbx_1__8__4_chanx_left_out[10] ,
    \cbx_1__8__4_chanx_left_out[11] ,
    \cbx_1__8__4_chanx_left_out[12] ,
    \cbx_1__8__4_chanx_left_out[13] ,
    \cbx_1__8__4_chanx_left_out[14] ,
    \cbx_1__8__4_chanx_left_out[15] ,
    \cbx_1__8__4_chanx_left_out[16] ,
    \cbx_1__8__4_chanx_left_out[17] ,
    \cbx_1__8__4_chanx_left_out[18] ,
    \cbx_1__8__4_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__8__4_chanx_left_out[0] ,
    \sb_1__8__4_chanx_left_out[1] ,
    \sb_1__8__4_chanx_left_out[2] ,
    \sb_1__8__4_chanx_left_out[3] ,
    \sb_1__8__4_chanx_left_out[4] ,
    \sb_1__8__4_chanx_left_out[5] ,
    \sb_1__8__4_chanx_left_out[6] ,
    \sb_1__8__4_chanx_left_out[7] ,
    \sb_1__8__4_chanx_left_out[8] ,
    \sb_1__8__4_chanx_left_out[9] ,
    \sb_1__8__4_chanx_left_out[10] ,
    \sb_1__8__4_chanx_left_out[11] ,
    \sb_1__8__4_chanx_left_out[12] ,
    \sb_1__8__4_chanx_left_out[13] ,
    \sb_1__8__4_chanx_left_out[14] ,
    \sb_1__8__4_chanx_left_out[15] ,
    \sb_1__8__4_chanx_left_out[16] ,
    \sb_1__8__4_chanx_left_out[17] ,
    \sb_1__8__4_chanx_left_out[18] ,
    \sb_1__8__4_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__4_chanx_right_out[0] ,
    \cbx_1__8__4_chanx_right_out[1] ,
    \cbx_1__8__4_chanx_right_out[2] ,
    \cbx_1__8__4_chanx_right_out[3] ,
    \cbx_1__8__4_chanx_right_out[4] ,
    \cbx_1__8__4_chanx_right_out[5] ,
    \cbx_1__8__4_chanx_right_out[6] ,
    \cbx_1__8__4_chanx_right_out[7] ,
    \cbx_1__8__4_chanx_right_out[8] ,
    \cbx_1__8__4_chanx_right_out[9] ,
    \cbx_1__8__4_chanx_right_out[10] ,
    \cbx_1__8__4_chanx_right_out[11] ,
    \cbx_1__8__4_chanx_right_out[12] ,
    \cbx_1__8__4_chanx_right_out[13] ,
    \cbx_1__8__4_chanx_right_out[14] ,
    \cbx_1__8__4_chanx_right_out[15] ,
    \cbx_1__8__4_chanx_right_out[16] ,
    \cbx_1__8__4_chanx_right_out[17] ,
    \cbx_1__8__4_chanx_right_out[18] ,
    \cbx_1__8__4_chanx_right_out[19] }));
 cbx_1__0_ cbx_6__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[93] ),
    .SC_OUT_TOP(\scff_Wires[94] ),
    .bottom_grid_pin_0_(cbx_1__0__5_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__5_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__5_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__5_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__5_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__5_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__5_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__5_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__5_bottom_grid_pin_8_),
    .ccff_head(sb_1__0__5_ccff_tail),
    .ccff_tail(grid_io_bottom_2_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[147] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__5_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__5_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_2_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_2_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__5_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_2_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_2_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__5_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_2_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_2_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__5_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_2_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_2_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_2_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_2_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__5_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_2_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_2_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__5_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_2_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_2_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__5_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_2_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_2_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__5_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_2_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_2_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__0__4_chanx_right_out[0] ,
    \sb_1__0__4_chanx_right_out[1] ,
    \sb_1__0__4_chanx_right_out[2] ,
    \sb_1__0__4_chanx_right_out[3] ,
    \sb_1__0__4_chanx_right_out[4] ,
    \sb_1__0__4_chanx_right_out[5] ,
    \sb_1__0__4_chanx_right_out[6] ,
    \sb_1__0__4_chanx_right_out[7] ,
    \sb_1__0__4_chanx_right_out[8] ,
    \sb_1__0__4_chanx_right_out[9] ,
    \sb_1__0__4_chanx_right_out[10] ,
    \sb_1__0__4_chanx_right_out[11] ,
    \sb_1__0__4_chanx_right_out[12] ,
    \sb_1__0__4_chanx_right_out[13] ,
    \sb_1__0__4_chanx_right_out[14] ,
    \sb_1__0__4_chanx_right_out[15] ,
    \sb_1__0__4_chanx_right_out[16] ,
    \sb_1__0__4_chanx_right_out[17] ,
    \sb_1__0__4_chanx_right_out[18] ,
    \sb_1__0__4_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__5_chanx_left_out[0] ,
    \cbx_1__0__5_chanx_left_out[1] ,
    \cbx_1__0__5_chanx_left_out[2] ,
    \cbx_1__0__5_chanx_left_out[3] ,
    \cbx_1__0__5_chanx_left_out[4] ,
    \cbx_1__0__5_chanx_left_out[5] ,
    \cbx_1__0__5_chanx_left_out[6] ,
    \cbx_1__0__5_chanx_left_out[7] ,
    \cbx_1__0__5_chanx_left_out[8] ,
    \cbx_1__0__5_chanx_left_out[9] ,
    \cbx_1__0__5_chanx_left_out[10] ,
    \cbx_1__0__5_chanx_left_out[11] ,
    \cbx_1__0__5_chanx_left_out[12] ,
    \cbx_1__0__5_chanx_left_out[13] ,
    \cbx_1__0__5_chanx_left_out[14] ,
    \cbx_1__0__5_chanx_left_out[15] ,
    \cbx_1__0__5_chanx_left_out[16] ,
    \cbx_1__0__5_chanx_left_out[17] ,
    \cbx_1__0__5_chanx_left_out[18] ,
    \cbx_1__0__5_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__0__5_chanx_left_out[0] ,
    \sb_1__0__5_chanx_left_out[1] ,
    \sb_1__0__5_chanx_left_out[2] ,
    \sb_1__0__5_chanx_left_out[3] ,
    \sb_1__0__5_chanx_left_out[4] ,
    \sb_1__0__5_chanx_left_out[5] ,
    \sb_1__0__5_chanx_left_out[6] ,
    \sb_1__0__5_chanx_left_out[7] ,
    \sb_1__0__5_chanx_left_out[8] ,
    \sb_1__0__5_chanx_left_out[9] ,
    \sb_1__0__5_chanx_left_out[10] ,
    \sb_1__0__5_chanx_left_out[11] ,
    \sb_1__0__5_chanx_left_out[12] ,
    \sb_1__0__5_chanx_left_out[13] ,
    \sb_1__0__5_chanx_left_out[14] ,
    \sb_1__0__5_chanx_left_out[15] ,
    \sb_1__0__5_chanx_left_out[16] ,
    \sb_1__0__5_chanx_left_out[17] ,
    \sb_1__0__5_chanx_left_out[18] ,
    \sb_1__0__5_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__5_chanx_right_out[0] ,
    \cbx_1__0__5_chanx_right_out[1] ,
    \cbx_1__0__5_chanx_right_out[2] ,
    \cbx_1__0__5_chanx_right_out[3] ,
    \cbx_1__0__5_chanx_right_out[4] ,
    \cbx_1__0__5_chanx_right_out[5] ,
    \cbx_1__0__5_chanx_right_out[6] ,
    \cbx_1__0__5_chanx_right_out[7] ,
    \cbx_1__0__5_chanx_right_out[8] ,
    \cbx_1__0__5_chanx_right_out[9] ,
    \cbx_1__0__5_chanx_right_out[10] ,
    \cbx_1__0__5_chanx_right_out[11] ,
    \cbx_1__0__5_chanx_right_out[12] ,
    \cbx_1__0__5_chanx_right_out[13] ,
    \cbx_1__0__5_chanx_right_out[14] ,
    \cbx_1__0__5_chanx_right_out[15] ,
    \cbx_1__0__5_chanx_right_out[16] ,
    \cbx_1__0__5_chanx_right_out[17] ,
    \cbx_1__0__5_chanx_right_out[18] ,
    \cbx_1__0__5_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]}));
 cbx_1__1_ cbx_6__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[35] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[35] ),
    .SC_IN_BOT(\scff_Wires[95] ),
    .SC_OUT_TOP(\scff_Wires[96] ),
    .bottom_grid_pin_0_(cbx_1__1__35_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__35_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__35_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__35_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__35_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__35_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__35_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__35_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__35_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__35_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__35_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__35_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__35_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__35_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__35_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__35_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__35_ccff_tail),
    .ccff_tail(cbx_1__1__35_ccff_tail),
    .clk_1_N_out(\clk_1_wires[61] ),
    .clk_1_S_out(\clk_1_wires[62] ),
    .clk_1_W_in(\clk_1_wires[57] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[150] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[61] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[62] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[57] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__28_chanx_right_out[0] ,
    \sb_1__1__28_chanx_right_out[1] ,
    \sb_1__1__28_chanx_right_out[2] ,
    \sb_1__1__28_chanx_right_out[3] ,
    \sb_1__1__28_chanx_right_out[4] ,
    \sb_1__1__28_chanx_right_out[5] ,
    \sb_1__1__28_chanx_right_out[6] ,
    \sb_1__1__28_chanx_right_out[7] ,
    \sb_1__1__28_chanx_right_out[8] ,
    \sb_1__1__28_chanx_right_out[9] ,
    \sb_1__1__28_chanx_right_out[10] ,
    \sb_1__1__28_chanx_right_out[11] ,
    \sb_1__1__28_chanx_right_out[12] ,
    \sb_1__1__28_chanx_right_out[13] ,
    \sb_1__1__28_chanx_right_out[14] ,
    \sb_1__1__28_chanx_right_out[15] ,
    \sb_1__1__28_chanx_right_out[16] ,
    \sb_1__1__28_chanx_right_out[17] ,
    \sb_1__1__28_chanx_right_out[18] ,
    \sb_1__1__28_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__35_chanx_left_out[0] ,
    \cbx_1__1__35_chanx_left_out[1] ,
    \cbx_1__1__35_chanx_left_out[2] ,
    \cbx_1__1__35_chanx_left_out[3] ,
    \cbx_1__1__35_chanx_left_out[4] ,
    \cbx_1__1__35_chanx_left_out[5] ,
    \cbx_1__1__35_chanx_left_out[6] ,
    \cbx_1__1__35_chanx_left_out[7] ,
    \cbx_1__1__35_chanx_left_out[8] ,
    \cbx_1__1__35_chanx_left_out[9] ,
    \cbx_1__1__35_chanx_left_out[10] ,
    \cbx_1__1__35_chanx_left_out[11] ,
    \cbx_1__1__35_chanx_left_out[12] ,
    \cbx_1__1__35_chanx_left_out[13] ,
    \cbx_1__1__35_chanx_left_out[14] ,
    \cbx_1__1__35_chanx_left_out[15] ,
    \cbx_1__1__35_chanx_left_out[16] ,
    \cbx_1__1__35_chanx_left_out[17] ,
    \cbx_1__1__35_chanx_left_out[18] ,
    \cbx_1__1__35_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__35_chanx_left_out[0] ,
    \sb_1__1__35_chanx_left_out[1] ,
    \sb_1__1__35_chanx_left_out[2] ,
    \sb_1__1__35_chanx_left_out[3] ,
    \sb_1__1__35_chanx_left_out[4] ,
    \sb_1__1__35_chanx_left_out[5] ,
    \sb_1__1__35_chanx_left_out[6] ,
    \sb_1__1__35_chanx_left_out[7] ,
    \sb_1__1__35_chanx_left_out[8] ,
    \sb_1__1__35_chanx_left_out[9] ,
    \sb_1__1__35_chanx_left_out[10] ,
    \sb_1__1__35_chanx_left_out[11] ,
    \sb_1__1__35_chanx_left_out[12] ,
    \sb_1__1__35_chanx_left_out[13] ,
    \sb_1__1__35_chanx_left_out[14] ,
    \sb_1__1__35_chanx_left_out[15] ,
    \sb_1__1__35_chanx_left_out[16] ,
    \sb_1__1__35_chanx_left_out[17] ,
    \sb_1__1__35_chanx_left_out[18] ,
    \sb_1__1__35_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__35_chanx_right_out[0] ,
    \cbx_1__1__35_chanx_right_out[1] ,
    \cbx_1__1__35_chanx_right_out[2] ,
    \cbx_1__1__35_chanx_right_out[3] ,
    \cbx_1__1__35_chanx_right_out[4] ,
    \cbx_1__1__35_chanx_right_out[5] ,
    \cbx_1__1__35_chanx_right_out[6] ,
    \cbx_1__1__35_chanx_right_out[7] ,
    \cbx_1__1__35_chanx_right_out[8] ,
    \cbx_1__1__35_chanx_right_out[9] ,
    \cbx_1__1__35_chanx_right_out[10] ,
    \cbx_1__1__35_chanx_right_out[11] ,
    \cbx_1__1__35_chanx_right_out[12] ,
    \cbx_1__1__35_chanx_right_out[13] ,
    \cbx_1__1__35_chanx_right_out[14] ,
    \cbx_1__1__35_chanx_right_out[15] ,
    \cbx_1__1__35_chanx_right_out[16] ,
    \cbx_1__1__35_chanx_right_out[17] ,
    \cbx_1__1__35_chanx_right_out[18] ,
    \cbx_1__1__35_chanx_right_out[19] }));
 cbx_1__1_ cbx_6__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[36] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[36] ),
    .SC_IN_BOT(\scff_Wires[97] ),
    .SC_OUT_TOP(\scff_Wires[98] ),
    .bottom_grid_pin_0_(cbx_1__1__36_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__36_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__36_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__36_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__36_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__36_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__36_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__36_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__36_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__36_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__36_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__36_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__36_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__36_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__36_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__36_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__36_ccff_tail),
    .ccff_tail(cbx_1__1__36_ccff_tail),
    .clk_2_W_in(\clk_2_wires[29] ),
    .clk_2_W_out(\clk_2_wires[30] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[153] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[29] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[30] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__29_chanx_right_out[0] ,
    \sb_1__1__29_chanx_right_out[1] ,
    \sb_1__1__29_chanx_right_out[2] ,
    \sb_1__1__29_chanx_right_out[3] ,
    \sb_1__1__29_chanx_right_out[4] ,
    \sb_1__1__29_chanx_right_out[5] ,
    \sb_1__1__29_chanx_right_out[6] ,
    \sb_1__1__29_chanx_right_out[7] ,
    \sb_1__1__29_chanx_right_out[8] ,
    \sb_1__1__29_chanx_right_out[9] ,
    \sb_1__1__29_chanx_right_out[10] ,
    \sb_1__1__29_chanx_right_out[11] ,
    \sb_1__1__29_chanx_right_out[12] ,
    \sb_1__1__29_chanx_right_out[13] ,
    \sb_1__1__29_chanx_right_out[14] ,
    \sb_1__1__29_chanx_right_out[15] ,
    \sb_1__1__29_chanx_right_out[16] ,
    \sb_1__1__29_chanx_right_out[17] ,
    \sb_1__1__29_chanx_right_out[18] ,
    \sb_1__1__29_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__36_chanx_left_out[0] ,
    \cbx_1__1__36_chanx_left_out[1] ,
    \cbx_1__1__36_chanx_left_out[2] ,
    \cbx_1__1__36_chanx_left_out[3] ,
    \cbx_1__1__36_chanx_left_out[4] ,
    \cbx_1__1__36_chanx_left_out[5] ,
    \cbx_1__1__36_chanx_left_out[6] ,
    \cbx_1__1__36_chanx_left_out[7] ,
    \cbx_1__1__36_chanx_left_out[8] ,
    \cbx_1__1__36_chanx_left_out[9] ,
    \cbx_1__1__36_chanx_left_out[10] ,
    \cbx_1__1__36_chanx_left_out[11] ,
    \cbx_1__1__36_chanx_left_out[12] ,
    \cbx_1__1__36_chanx_left_out[13] ,
    \cbx_1__1__36_chanx_left_out[14] ,
    \cbx_1__1__36_chanx_left_out[15] ,
    \cbx_1__1__36_chanx_left_out[16] ,
    \cbx_1__1__36_chanx_left_out[17] ,
    \cbx_1__1__36_chanx_left_out[18] ,
    \cbx_1__1__36_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__36_chanx_left_out[0] ,
    \sb_1__1__36_chanx_left_out[1] ,
    \sb_1__1__36_chanx_left_out[2] ,
    \sb_1__1__36_chanx_left_out[3] ,
    \sb_1__1__36_chanx_left_out[4] ,
    \sb_1__1__36_chanx_left_out[5] ,
    \sb_1__1__36_chanx_left_out[6] ,
    \sb_1__1__36_chanx_left_out[7] ,
    \sb_1__1__36_chanx_left_out[8] ,
    \sb_1__1__36_chanx_left_out[9] ,
    \sb_1__1__36_chanx_left_out[10] ,
    \sb_1__1__36_chanx_left_out[11] ,
    \sb_1__1__36_chanx_left_out[12] ,
    \sb_1__1__36_chanx_left_out[13] ,
    \sb_1__1__36_chanx_left_out[14] ,
    \sb_1__1__36_chanx_left_out[15] ,
    \sb_1__1__36_chanx_left_out[16] ,
    \sb_1__1__36_chanx_left_out[17] ,
    \sb_1__1__36_chanx_left_out[18] ,
    \sb_1__1__36_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__36_chanx_right_out[0] ,
    \cbx_1__1__36_chanx_right_out[1] ,
    \cbx_1__1__36_chanx_right_out[2] ,
    \cbx_1__1__36_chanx_right_out[3] ,
    \cbx_1__1__36_chanx_right_out[4] ,
    \cbx_1__1__36_chanx_right_out[5] ,
    \cbx_1__1__36_chanx_right_out[6] ,
    \cbx_1__1__36_chanx_right_out[7] ,
    \cbx_1__1__36_chanx_right_out[8] ,
    \cbx_1__1__36_chanx_right_out[9] ,
    \cbx_1__1__36_chanx_right_out[10] ,
    \cbx_1__1__36_chanx_right_out[11] ,
    \cbx_1__1__36_chanx_right_out[12] ,
    \cbx_1__1__36_chanx_right_out[13] ,
    \cbx_1__1__36_chanx_right_out[14] ,
    \cbx_1__1__36_chanx_right_out[15] ,
    \cbx_1__1__36_chanx_right_out[16] ,
    \cbx_1__1__36_chanx_right_out[17] ,
    \cbx_1__1__36_chanx_right_out[18] ,
    \cbx_1__1__36_chanx_right_out[19] }));
 cbx_1__1_ cbx_6__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[37] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[37] ),
    .SC_IN_BOT(\scff_Wires[99] ),
    .SC_OUT_TOP(\scff_Wires[100] ),
    .bottom_grid_pin_0_(cbx_1__1__37_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__37_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__37_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__37_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__37_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__37_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__37_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__37_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__37_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__37_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__37_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__37_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__37_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__37_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__37_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__37_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__37_ccff_tail),
    .ccff_tail(cbx_1__1__37_ccff_tail),
    .clk_1_N_out(\clk_1_wires[68] ),
    .clk_1_S_out(\clk_1_wires[69] ),
    .clk_1_W_in(\clk_1_wires[64] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[156] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[68] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[69] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[64] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__30_chanx_right_out[0] ,
    \sb_1__1__30_chanx_right_out[1] ,
    \sb_1__1__30_chanx_right_out[2] ,
    \sb_1__1__30_chanx_right_out[3] ,
    \sb_1__1__30_chanx_right_out[4] ,
    \sb_1__1__30_chanx_right_out[5] ,
    \sb_1__1__30_chanx_right_out[6] ,
    \sb_1__1__30_chanx_right_out[7] ,
    \sb_1__1__30_chanx_right_out[8] ,
    \sb_1__1__30_chanx_right_out[9] ,
    \sb_1__1__30_chanx_right_out[10] ,
    \sb_1__1__30_chanx_right_out[11] ,
    \sb_1__1__30_chanx_right_out[12] ,
    \sb_1__1__30_chanx_right_out[13] ,
    \sb_1__1__30_chanx_right_out[14] ,
    \sb_1__1__30_chanx_right_out[15] ,
    \sb_1__1__30_chanx_right_out[16] ,
    \sb_1__1__30_chanx_right_out[17] ,
    \sb_1__1__30_chanx_right_out[18] ,
    \sb_1__1__30_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__37_chanx_left_out[0] ,
    \cbx_1__1__37_chanx_left_out[1] ,
    \cbx_1__1__37_chanx_left_out[2] ,
    \cbx_1__1__37_chanx_left_out[3] ,
    \cbx_1__1__37_chanx_left_out[4] ,
    \cbx_1__1__37_chanx_left_out[5] ,
    \cbx_1__1__37_chanx_left_out[6] ,
    \cbx_1__1__37_chanx_left_out[7] ,
    \cbx_1__1__37_chanx_left_out[8] ,
    \cbx_1__1__37_chanx_left_out[9] ,
    \cbx_1__1__37_chanx_left_out[10] ,
    \cbx_1__1__37_chanx_left_out[11] ,
    \cbx_1__1__37_chanx_left_out[12] ,
    \cbx_1__1__37_chanx_left_out[13] ,
    \cbx_1__1__37_chanx_left_out[14] ,
    \cbx_1__1__37_chanx_left_out[15] ,
    \cbx_1__1__37_chanx_left_out[16] ,
    \cbx_1__1__37_chanx_left_out[17] ,
    \cbx_1__1__37_chanx_left_out[18] ,
    \cbx_1__1__37_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__37_chanx_left_out[0] ,
    \sb_1__1__37_chanx_left_out[1] ,
    \sb_1__1__37_chanx_left_out[2] ,
    \sb_1__1__37_chanx_left_out[3] ,
    \sb_1__1__37_chanx_left_out[4] ,
    \sb_1__1__37_chanx_left_out[5] ,
    \sb_1__1__37_chanx_left_out[6] ,
    \sb_1__1__37_chanx_left_out[7] ,
    \sb_1__1__37_chanx_left_out[8] ,
    \sb_1__1__37_chanx_left_out[9] ,
    \sb_1__1__37_chanx_left_out[10] ,
    \sb_1__1__37_chanx_left_out[11] ,
    \sb_1__1__37_chanx_left_out[12] ,
    \sb_1__1__37_chanx_left_out[13] ,
    \sb_1__1__37_chanx_left_out[14] ,
    \sb_1__1__37_chanx_left_out[15] ,
    \sb_1__1__37_chanx_left_out[16] ,
    \sb_1__1__37_chanx_left_out[17] ,
    \sb_1__1__37_chanx_left_out[18] ,
    \sb_1__1__37_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__37_chanx_right_out[0] ,
    \cbx_1__1__37_chanx_right_out[1] ,
    \cbx_1__1__37_chanx_right_out[2] ,
    \cbx_1__1__37_chanx_right_out[3] ,
    \cbx_1__1__37_chanx_right_out[4] ,
    \cbx_1__1__37_chanx_right_out[5] ,
    \cbx_1__1__37_chanx_right_out[6] ,
    \cbx_1__1__37_chanx_right_out[7] ,
    \cbx_1__1__37_chanx_right_out[8] ,
    \cbx_1__1__37_chanx_right_out[9] ,
    \cbx_1__1__37_chanx_right_out[10] ,
    \cbx_1__1__37_chanx_right_out[11] ,
    \cbx_1__1__37_chanx_right_out[12] ,
    \cbx_1__1__37_chanx_right_out[13] ,
    \cbx_1__1__37_chanx_right_out[14] ,
    \cbx_1__1__37_chanx_right_out[15] ,
    \cbx_1__1__37_chanx_right_out[16] ,
    \cbx_1__1__37_chanx_right_out[17] ,
    \cbx_1__1__37_chanx_right_out[18] ,
    \cbx_1__1__37_chanx_right_out[19] }));
 cbx_1__1_ cbx_6__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[38] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[38] ),
    .SC_IN_BOT(\scff_Wires[101] ),
    .SC_OUT_TOP(\scff_Wires[102] ),
    .bottom_grid_pin_0_(cbx_1__1__38_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__38_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__38_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__38_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__38_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__38_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__38_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__38_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__38_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__38_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__38_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__38_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__38_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__38_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__38_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__38_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__38_ccff_tail),
    .ccff_tail(cbx_1__1__38_ccff_tail),
    .clk_3_E_out(\clk_3_wires[7] ),
    .clk_3_W_in(\clk_3_wires[6] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[159] ),
    .prog_clk_3_E_out(\prog_clk_3_wires[7] ),
    .prog_clk_3_W_in(\prog_clk_3_wires[6] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__31_chanx_right_out[0] ,
    \sb_1__1__31_chanx_right_out[1] ,
    \sb_1__1__31_chanx_right_out[2] ,
    \sb_1__1__31_chanx_right_out[3] ,
    \sb_1__1__31_chanx_right_out[4] ,
    \sb_1__1__31_chanx_right_out[5] ,
    \sb_1__1__31_chanx_right_out[6] ,
    \sb_1__1__31_chanx_right_out[7] ,
    \sb_1__1__31_chanx_right_out[8] ,
    \sb_1__1__31_chanx_right_out[9] ,
    \sb_1__1__31_chanx_right_out[10] ,
    \sb_1__1__31_chanx_right_out[11] ,
    \sb_1__1__31_chanx_right_out[12] ,
    \sb_1__1__31_chanx_right_out[13] ,
    \sb_1__1__31_chanx_right_out[14] ,
    \sb_1__1__31_chanx_right_out[15] ,
    \sb_1__1__31_chanx_right_out[16] ,
    \sb_1__1__31_chanx_right_out[17] ,
    \sb_1__1__31_chanx_right_out[18] ,
    \sb_1__1__31_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__38_chanx_left_out[0] ,
    \cbx_1__1__38_chanx_left_out[1] ,
    \cbx_1__1__38_chanx_left_out[2] ,
    \cbx_1__1__38_chanx_left_out[3] ,
    \cbx_1__1__38_chanx_left_out[4] ,
    \cbx_1__1__38_chanx_left_out[5] ,
    \cbx_1__1__38_chanx_left_out[6] ,
    \cbx_1__1__38_chanx_left_out[7] ,
    \cbx_1__1__38_chanx_left_out[8] ,
    \cbx_1__1__38_chanx_left_out[9] ,
    \cbx_1__1__38_chanx_left_out[10] ,
    \cbx_1__1__38_chanx_left_out[11] ,
    \cbx_1__1__38_chanx_left_out[12] ,
    \cbx_1__1__38_chanx_left_out[13] ,
    \cbx_1__1__38_chanx_left_out[14] ,
    \cbx_1__1__38_chanx_left_out[15] ,
    \cbx_1__1__38_chanx_left_out[16] ,
    \cbx_1__1__38_chanx_left_out[17] ,
    \cbx_1__1__38_chanx_left_out[18] ,
    \cbx_1__1__38_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__38_chanx_left_out[0] ,
    \sb_1__1__38_chanx_left_out[1] ,
    \sb_1__1__38_chanx_left_out[2] ,
    \sb_1__1__38_chanx_left_out[3] ,
    \sb_1__1__38_chanx_left_out[4] ,
    \sb_1__1__38_chanx_left_out[5] ,
    \sb_1__1__38_chanx_left_out[6] ,
    \sb_1__1__38_chanx_left_out[7] ,
    \sb_1__1__38_chanx_left_out[8] ,
    \sb_1__1__38_chanx_left_out[9] ,
    \sb_1__1__38_chanx_left_out[10] ,
    \sb_1__1__38_chanx_left_out[11] ,
    \sb_1__1__38_chanx_left_out[12] ,
    \sb_1__1__38_chanx_left_out[13] ,
    \sb_1__1__38_chanx_left_out[14] ,
    \sb_1__1__38_chanx_left_out[15] ,
    \sb_1__1__38_chanx_left_out[16] ,
    \sb_1__1__38_chanx_left_out[17] ,
    \sb_1__1__38_chanx_left_out[18] ,
    \sb_1__1__38_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__38_chanx_right_out[0] ,
    \cbx_1__1__38_chanx_right_out[1] ,
    \cbx_1__1__38_chanx_right_out[2] ,
    \cbx_1__1__38_chanx_right_out[3] ,
    \cbx_1__1__38_chanx_right_out[4] ,
    \cbx_1__1__38_chanx_right_out[5] ,
    \cbx_1__1__38_chanx_right_out[6] ,
    \cbx_1__1__38_chanx_right_out[7] ,
    \cbx_1__1__38_chanx_right_out[8] ,
    \cbx_1__1__38_chanx_right_out[9] ,
    \cbx_1__1__38_chanx_right_out[10] ,
    \cbx_1__1__38_chanx_right_out[11] ,
    \cbx_1__1__38_chanx_right_out[12] ,
    \cbx_1__1__38_chanx_right_out[13] ,
    \cbx_1__1__38_chanx_right_out[14] ,
    \cbx_1__1__38_chanx_right_out[15] ,
    \cbx_1__1__38_chanx_right_out[16] ,
    \cbx_1__1__38_chanx_right_out[17] ,
    \cbx_1__1__38_chanx_right_out[18] ,
    \cbx_1__1__38_chanx_right_out[19] }));
 cbx_1__1_ cbx_6__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[39] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[39] ),
    .SC_IN_BOT(\scff_Wires[103] ),
    .SC_OUT_TOP(\scff_Wires[104] ),
    .bottom_grid_pin_0_(cbx_1__1__39_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__39_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__39_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__39_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__39_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__39_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__39_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__39_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__39_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__39_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__39_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__39_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__39_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__39_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__39_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__39_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__39_ccff_tail),
    .ccff_tail(cbx_1__1__39_ccff_tail),
    .clk_1_N_out(\clk_1_wires[75] ),
    .clk_1_S_out(\clk_1_wires[76] ),
    .clk_1_W_in(\clk_1_wires[71] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[162] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[75] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[76] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[71] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__32_chanx_right_out[0] ,
    \sb_1__1__32_chanx_right_out[1] ,
    \sb_1__1__32_chanx_right_out[2] ,
    \sb_1__1__32_chanx_right_out[3] ,
    \sb_1__1__32_chanx_right_out[4] ,
    \sb_1__1__32_chanx_right_out[5] ,
    \sb_1__1__32_chanx_right_out[6] ,
    \sb_1__1__32_chanx_right_out[7] ,
    \sb_1__1__32_chanx_right_out[8] ,
    \sb_1__1__32_chanx_right_out[9] ,
    \sb_1__1__32_chanx_right_out[10] ,
    \sb_1__1__32_chanx_right_out[11] ,
    \sb_1__1__32_chanx_right_out[12] ,
    \sb_1__1__32_chanx_right_out[13] ,
    \sb_1__1__32_chanx_right_out[14] ,
    \sb_1__1__32_chanx_right_out[15] ,
    \sb_1__1__32_chanx_right_out[16] ,
    \sb_1__1__32_chanx_right_out[17] ,
    \sb_1__1__32_chanx_right_out[18] ,
    \sb_1__1__32_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__39_chanx_left_out[0] ,
    \cbx_1__1__39_chanx_left_out[1] ,
    \cbx_1__1__39_chanx_left_out[2] ,
    \cbx_1__1__39_chanx_left_out[3] ,
    \cbx_1__1__39_chanx_left_out[4] ,
    \cbx_1__1__39_chanx_left_out[5] ,
    \cbx_1__1__39_chanx_left_out[6] ,
    \cbx_1__1__39_chanx_left_out[7] ,
    \cbx_1__1__39_chanx_left_out[8] ,
    \cbx_1__1__39_chanx_left_out[9] ,
    \cbx_1__1__39_chanx_left_out[10] ,
    \cbx_1__1__39_chanx_left_out[11] ,
    \cbx_1__1__39_chanx_left_out[12] ,
    \cbx_1__1__39_chanx_left_out[13] ,
    \cbx_1__1__39_chanx_left_out[14] ,
    \cbx_1__1__39_chanx_left_out[15] ,
    \cbx_1__1__39_chanx_left_out[16] ,
    \cbx_1__1__39_chanx_left_out[17] ,
    \cbx_1__1__39_chanx_left_out[18] ,
    \cbx_1__1__39_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__39_chanx_left_out[0] ,
    \sb_1__1__39_chanx_left_out[1] ,
    \sb_1__1__39_chanx_left_out[2] ,
    \sb_1__1__39_chanx_left_out[3] ,
    \sb_1__1__39_chanx_left_out[4] ,
    \sb_1__1__39_chanx_left_out[5] ,
    \sb_1__1__39_chanx_left_out[6] ,
    \sb_1__1__39_chanx_left_out[7] ,
    \sb_1__1__39_chanx_left_out[8] ,
    \sb_1__1__39_chanx_left_out[9] ,
    \sb_1__1__39_chanx_left_out[10] ,
    \sb_1__1__39_chanx_left_out[11] ,
    \sb_1__1__39_chanx_left_out[12] ,
    \sb_1__1__39_chanx_left_out[13] ,
    \sb_1__1__39_chanx_left_out[14] ,
    \sb_1__1__39_chanx_left_out[15] ,
    \sb_1__1__39_chanx_left_out[16] ,
    \sb_1__1__39_chanx_left_out[17] ,
    \sb_1__1__39_chanx_left_out[18] ,
    \sb_1__1__39_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__39_chanx_right_out[0] ,
    \cbx_1__1__39_chanx_right_out[1] ,
    \cbx_1__1__39_chanx_right_out[2] ,
    \cbx_1__1__39_chanx_right_out[3] ,
    \cbx_1__1__39_chanx_right_out[4] ,
    \cbx_1__1__39_chanx_right_out[5] ,
    \cbx_1__1__39_chanx_right_out[6] ,
    \cbx_1__1__39_chanx_right_out[7] ,
    \cbx_1__1__39_chanx_right_out[8] ,
    \cbx_1__1__39_chanx_right_out[9] ,
    \cbx_1__1__39_chanx_right_out[10] ,
    \cbx_1__1__39_chanx_right_out[11] ,
    \cbx_1__1__39_chanx_right_out[12] ,
    \cbx_1__1__39_chanx_right_out[13] ,
    \cbx_1__1__39_chanx_right_out[14] ,
    \cbx_1__1__39_chanx_right_out[15] ,
    \cbx_1__1__39_chanx_right_out[16] ,
    \cbx_1__1__39_chanx_right_out[17] ,
    \cbx_1__1__39_chanx_right_out[18] ,
    \cbx_1__1__39_chanx_right_out[19] }));
 cbx_1__1_ cbx_6__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[40] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[40] ),
    .SC_IN_BOT(\scff_Wires[105] ),
    .SC_OUT_TOP(\scff_Wires[106] ),
    .bottom_grid_pin_0_(cbx_1__1__40_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__40_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__40_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__40_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__40_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__40_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__40_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__40_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__40_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__40_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__40_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__40_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__40_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__40_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__40_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__40_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__40_ccff_tail),
    .ccff_tail(cbx_1__1__40_ccff_tail),
    .clk_2_W_in(\clk_2_wires[42] ),
    .clk_2_W_out(\clk_2_wires[43] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[165] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[42] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[43] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__33_chanx_right_out[0] ,
    \sb_1__1__33_chanx_right_out[1] ,
    \sb_1__1__33_chanx_right_out[2] ,
    \sb_1__1__33_chanx_right_out[3] ,
    \sb_1__1__33_chanx_right_out[4] ,
    \sb_1__1__33_chanx_right_out[5] ,
    \sb_1__1__33_chanx_right_out[6] ,
    \sb_1__1__33_chanx_right_out[7] ,
    \sb_1__1__33_chanx_right_out[8] ,
    \sb_1__1__33_chanx_right_out[9] ,
    \sb_1__1__33_chanx_right_out[10] ,
    \sb_1__1__33_chanx_right_out[11] ,
    \sb_1__1__33_chanx_right_out[12] ,
    \sb_1__1__33_chanx_right_out[13] ,
    \sb_1__1__33_chanx_right_out[14] ,
    \sb_1__1__33_chanx_right_out[15] ,
    \sb_1__1__33_chanx_right_out[16] ,
    \sb_1__1__33_chanx_right_out[17] ,
    \sb_1__1__33_chanx_right_out[18] ,
    \sb_1__1__33_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__40_chanx_left_out[0] ,
    \cbx_1__1__40_chanx_left_out[1] ,
    \cbx_1__1__40_chanx_left_out[2] ,
    \cbx_1__1__40_chanx_left_out[3] ,
    \cbx_1__1__40_chanx_left_out[4] ,
    \cbx_1__1__40_chanx_left_out[5] ,
    \cbx_1__1__40_chanx_left_out[6] ,
    \cbx_1__1__40_chanx_left_out[7] ,
    \cbx_1__1__40_chanx_left_out[8] ,
    \cbx_1__1__40_chanx_left_out[9] ,
    \cbx_1__1__40_chanx_left_out[10] ,
    \cbx_1__1__40_chanx_left_out[11] ,
    \cbx_1__1__40_chanx_left_out[12] ,
    \cbx_1__1__40_chanx_left_out[13] ,
    \cbx_1__1__40_chanx_left_out[14] ,
    \cbx_1__1__40_chanx_left_out[15] ,
    \cbx_1__1__40_chanx_left_out[16] ,
    \cbx_1__1__40_chanx_left_out[17] ,
    \cbx_1__1__40_chanx_left_out[18] ,
    \cbx_1__1__40_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__40_chanx_left_out[0] ,
    \sb_1__1__40_chanx_left_out[1] ,
    \sb_1__1__40_chanx_left_out[2] ,
    \sb_1__1__40_chanx_left_out[3] ,
    \sb_1__1__40_chanx_left_out[4] ,
    \sb_1__1__40_chanx_left_out[5] ,
    \sb_1__1__40_chanx_left_out[6] ,
    \sb_1__1__40_chanx_left_out[7] ,
    \sb_1__1__40_chanx_left_out[8] ,
    \sb_1__1__40_chanx_left_out[9] ,
    \sb_1__1__40_chanx_left_out[10] ,
    \sb_1__1__40_chanx_left_out[11] ,
    \sb_1__1__40_chanx_left_out[12] ,
    \sb_1__1__40_chanx_left_out[13] ,
    \sb_1__1__40_chanx_left_out[14] ,
    \sb_1__1__40_chanx_left_out[15] ,
    \sb_1__1__40_chanx_left_out[16] ,
    \sb_1__1__40_chanx_left_out[17] ,
    \sb_1__1__40_chanx_left_out[18] ,
    \sb_1__1__40_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__40_chanx_right_out[0] ,
    \cbx_1__1__40_chanx_right_out[1] ,
    \cbx_1__1__40_chanx_right_out[2] ,
    \cbx_1__1__40_chanx_right_out[3] ,
    \cbx_1__1__40_chanx_right_out[4] ,
    \cbx_1__1__40_chanx_right_out[5] ,
    \cbx_1__1__40_chanx_right_out[6] ,
    \cbx_1__1__40_chanx_right_out[7] ,
    \cbx_1__1__40_chanx_right_out[8] ,
    \cbx_1__1__40_chanx_right_out[9] ,
    \cbx_1__1__40_chanx_right_out[10] ,
    \cbx_1__1__40_chanx_right_out[11] ,
    \cbx_1__1__40_chanx_right_out[12] ,
    \cbx_1__1__40_chanx_right_out[13] ,
    \cbx_1__1__40_chanx_right_out[14] ,
    \cbx_1__1__40_chanx_right_out[15] ,
    \cbx_1__1__40_chanx_right_out[16] ,
    \cbx_1__1__40_chanx_right_out[17] ,
    \cbx_1__1__40_chanx_right_out[18] ,
    \cbx_1__1__40_chanx_right_out[19] }));
 cbx_1__1_ cbx_6__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[41] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[41] ),
    .SC_IN_BOT(\scff_Wires[107] ),
    .SC_OUT_TOP(\scff_Wires[108] ),
    .bottom_grid_pin_0_(cbx_1__1__41_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__41_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__41_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__41_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__41_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__41_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__41_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__41_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__41_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__41_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__41_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__41_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__41_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__41_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__41_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__41_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__41_ccff_tail),
    .ccff_tail(cbx_1__1__41_ccff_tail),
    .clk_1_N_out(\clk_1_wires[82] ),
    .clk_1_S_out(\clk_1_wires[83] ),
    .clk_1_W_in(\clk_1_wires[78] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[168] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[82] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[83] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[78] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__34_chanx_right_out[0] ,
    \sb_1__1__34_chanx_right_out[1] ,
    \sb_1__1__34_chanx_right_out[2] ,
    \sb_1__1__34_chanx_right_out[3] ,
    \sb_1__1__34_chanx_right_out[4] ,
    \sb_1__1__34_chanx_right_out[5] ,
    \sb_1__1__34_chanx_right_out[6] ,
    \sb_1__1__34_chanx_right_out[7] ,
    \sb_1__1__34_chanx_right_out[8] ,
    \sb_1__1__34_chanx_right_out[9] ,
    \sb_1__1__34_chanx_right_out[10] ,
    \sb_1__1__34_chanx_right_out[11] ,
    \sb_1__1__34_chanx_right_out[12] ,
    \sb_1__1__34_chanx_right_out[13] ,
    \sb_1__1__34_chanx_right_out[14] ,
    \sb_1__1__34_chanx_right_out[15] ,
    \sb_1__1__34_chanx_right_out[16] ,
    \sb_1__1__34_chanx_right_out[17] ,
    \sb_1__1__34_chanx_right_out[18] ,
    \sb_1__1__34_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__41_chanx_left_out[0] ,
    \cbx_1__1__41_chanx_left_out[1] ,
    \cbx_1__1__41_chanx_left_out[2] ,
    \cbx_1__1__41_chanx_left_out[3] ,
    \cbx_1__1__41_chanx_left_out[4] ,
    \cbx_1__1__41_chanx_left_out[5] ,
    \cbx_1__1__41_chanx_left_out[6] ,
    \cbx_1__1__41_chanx_left_out[7] ,
    \cbx_1__1__41_chanx_left_out[8] ,
    \cbx_1__1__41_chanx_left_out[9] ,
    \cbx_1__1__41_chanx_left_out[10] ,
    \cbx_1__1__41_chanx_left_out[11] ,
    \cbx_1__1__41_chanx_left_out[12] ,
    \cbx_1__1__41_chanx_left_out[13] ,
    \cbx_1__1__41_chanx_left_out[14] ,
    \cbx_1__1__41_chanx_left_out[15] ,
    \cbx_1__1__41_chanx_left_out[16] ,
    \cbx_1__1__41_chanx_left_out[17] ,
    \cbx_1__1__41_chanx_left_out[18] ,
    \cbx_1__1__41_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__41_chanx_left_out[0] ,
    \sb_1__1__41_chanx_left_out[1] ,
    \sb_1__1__41_chanx_left_out[2] ,
    \sb_1__1__41_chanx_left_out[3] ,
    \sb_1__1__41_chanx_left_out[4] ,
    \sb_1__1__41_chanx_left_out[5] ,
    \sb_1__1__41_chanx_left_out[6] ,
    \sb_1__1__41_chanx_left_out[7] ,
    \sb_1__1__41_chanx_left_out[8] ,
    \sb_1__1__41_chanx_left_out[9] ,
    \sb_1__1__41_chanx_left_out[10] ,
    \sb_1__1__41_chanx_left_out[11] ,
    \sb_1__1__41_chanx_left_out[12] ,
    \sb_1__1__41_chanx_left_out[13] ,
    \sb_1__1__41_chanx_left_out[14] ,
    \sb_1__1__41_chanx_left_out[15] ,
    \sb_1__1__41_chanx_left_out[16] ,
    \sb_1__1__41_chanx_left_out[17] ,
    \sb_1__1__41_chanx_left_out[18] ,
    \sb_1__1__41_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__41_chanx_right_out[0] ,
    \cbx_1__1__41_chanx_right_out[1] ,
    \cbx_1__1__41_chanx_right_out[2] ,
    \cbx_1__1__41_chanx_right_out[3] ,
    \cbx_1__1__41_chanx_right_out[4] ,
    \cbx_1__1__41_chanx_right_out[5] ,
    \cbx_1__1__41_chanx_right_out[6] ,
    \cbx_1__1__41_chanx_right_out[7] ,
    \cbx_1__1__41_chanx_right_out[8] ,
    \cbx_1__1__41_chanx_right_out[9] ,
    \cbx_1__1__41_chanx_right_out[10] ,
    \cbx_1__1__41_chanx_right_out[11] ,
    \cbx_1__1__41_chanx_right_out[12] ,
    \cbx_1__1__41_chanx_right_out[13] ,
    \cbx_1__1__41_chanx_right_out[14] ,
    \cbx_1__1__41_chanx_right_out[15] ,
    \cbx_1__1__41_chanx_right_out[16] ,
    \cbx_1__1__41_chanx_right_out[17] ,
    \cbx_1__1__41_chanx_right_out[18] ,
    \cbx_1__1__41_chanx_right_out[19] }));
 cbx_1__2_ cbx_6__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[109] ),
    .SC_OUT_TOP(\scff_Wires[110] ),
    .bottom_grid_pin_0_(cbx_1__8__5_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__5_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__5_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__5_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__5_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__5_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__5_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__5_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__5_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__5_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__5_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__5_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__5_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__5_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__5_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__5_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__5_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_5_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_5_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_1__8__5_ccff_tail),
    .ccff_tail(grid_io_top_5_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]),
    .prog_clk_0_S_in(\prog_clk_0_wires[171] ),
    .top_grid_pin_0_(cbx_1__8__5_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__8__4_chanx_right_out[0] ,
    \sb_1__8__4_chanx_right_out[1] ,
    \sb_1__8__4_chanx_right_out[2] ,
    \sb_1__8__4_chanx_right_out[3] ,
    \sb_1__8__4_chanx_right_out[4] ,
    \sb_1__8__4_chanx_right_out[5] ,
    \sb_1__8__4_chanx_right_out[6] ,
    \sb_1__8__4_chanx_right_out[7] ,
    \sb_1__8__4_chanx_right_out[8] ,
    \sb_1__8__4_chanx_right_out[9] ,
    \sb_1__8__4_chanx_right_out[10] ,
    \sb_1__8__4_chanx_right_out[11] ,
    \sb_1__8__4_chanx_right_out[12] ,
    \sb_1__8__4_chanx_right_out[13] ,
    \sb_1__8__4_chanx_right_out[14] ,
    \sb_1__8__4_chanx_right_out[15] ,
    \sb_1__8__4_chanx_right_out[16] ,
    \sb_1__8__4_chanx_right_out[17] ,
    \sb_1__8__4_chanx_right_out[18] ,
    \sb_1__8__4_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__5_chanx_left_out[0] ,
    \cbx_1__8__5_chanx_left_out[1] ,
    \cbx_1__8__5_chanx_left_out[2] ,
    \cbx_1__8__5_chanx_left_out[3] ,
    \cbx_1__8__5_chanx_left_out[4] ,
    \cbx_1__8__5_chanx_left_out[5] ,
    \cbx_1__8__5_chanx_left_out[6] ,
    \cbx_1__8__5_chanx_left_out[7] ,
    \cbx_1__8__5_chanx_left_out[8] ,
    \cbx_1__8__5_chanx_left_out[9] ,
    \cbx_1__8__5_chanx_left_out[10] ,
    \cbx_1__8__5_chanx_left_out[11] ,
    \cbx_1__8__5_chanx_left_out[12] ,
    \cbx_1__8__5_chanx_left_out[13] ,
    \cbx_1__8__5_chanx_left_out[14] ,
    \cbx_1__8__5_chanx_left_out[15] ,
    \cbx_1__8__5_chanx_left_out[16] ,
    \cbx_1__8__5_chanx_left_out[17] ,
    \cbx_1__8__5_chanx_left_out[18] ,
    \cbx_1__8__5_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__8__5_chanx_left_out[0] ,
    \sb_1__8__5_chanx_left_out[1] ,
    \sb_1__8__5_chanx_left_out[2] ,
    \sb_1__8__5_chanx_left_out[3] ,
    \sb_1__8__5_chanx_left_out[4] ,
    \sb_1__8__5_chanx_left_out[5] ,
    \sb_1__8__5_chanx_left_out[6] ,
    \sb_1__8__5_chanx_left_out[7] ,
    \sb_1__8__5_chanx_left_out[8] ,
    \sb_1__8__5_chanx_left_out[9] ,
    \sb_1__8__5_chanx_left_out[10] ,
    \sb_1__8__5_chanx_left_out[11] ,
    \sb_1__8__5_chanx_left_out[12] ,
    \sb_1__8__5_chanx_left_out[13] ,
    \sb_1__8__5_chanx_left_out[14] ,
    \sb_1__8__5_chanx_left_out[15] ,
    \sb_1__8__5_chanx_left_out[16] ,
    \sb_1__8__5_chanx_left_out[17] ,
    \sb_1__8__5_chanx_left_out[18] ,
    \sb_1__8__5_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__5_chanx_right_out[0] ,
    \cbx_1__8__5_chanx_right_out[1] ,
    \cbx_1__8__5_chanx_right_out[2] ,
    \cbx_1__8__5_chanx_right_out[3] ,
    \cbx_1__8__5_chanx_right_out[4] ,
    \cbx_1__8__5_chanx_right_out[5] ,
    \cbx_1__8__5_chanx_right_out[6] ,
    \cbx_1__8__5_chanx_right_out[7] ,
    \cbx_1__8__5_chanx_right_out[8] ,
    \cbx_1__8__5_chanx_right_out[9] ,
    \cbx_1__8__5_chanx_right_out[10] ,
    \cbx_1__8__5_chanx_right_out[11] ,
    \cbx_1__8__5_chanx_right_out[12] ,
    \cbx_1__8__5_chanx_right_out[13] ,
    \cbx_1__8__5_chanx_right_out[14] ,
    \cbx_1__8__5_chanx_right_out[15] ,
    \cbx_1__8__5_chanx_right_out[16] ,
    \cbx_1__8__5_chanx_right_out[17] ,
    \cbx_1__8__5_chanx_right_out[18] ,
    \cbx_1__8__5_chanx_right_out[19] }));
 cbx_1__0_ cbx_7__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[128] ),
    .SC_OUT_BOT(\scff_Wires[129] ),
    .bottom_grid_pin_0_(cbx_1__0__6_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__6_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__6_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__6_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__6_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__6_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__6_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__6_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__6_bottom_grid_pin_8_),
    .ccff_head(sb_1__0__6_ccff_tail),
    .ccff_tail(grid_io_bottom_1_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[173] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__6_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__6_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_1_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_1_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__6_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_1_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_1_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__6_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_1_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_1_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__6_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_1_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_1_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_1_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_1_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__6_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_1_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_1_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__6_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_1_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_1_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__6_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_1_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_1_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__6_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_1_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_1_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__0__5_chanx_right_out[0] ,
    \sb_1__0__5_chanx_right_out[1] ,
    \sb_1__0__5_chanx_right_out[2] ,
    \sb_1__0__5_chanx_right_out[3] ,
    \sb_1__0__5_chanx_right_out[4] ,
    \sb_1__0__5_chanx_right_out[5] ,
    \sb_1__0__5_chanx_right_out[6] ,
    \sb_1__0__5_chanx_right_out[7] ,
    \sb_1__0__5_chanx_right_out[8] ,
    \sb_1__0__5_chanx_right_out[9] ,
    \sb_1__0__5_chanx_right_out[10] ,
    \sb_1__0__5_chanx_right_out[11] ,
    \sb_1__0__5_chanx_right_out[12] ,
    \sb_1__0__5_chanx_right_out[13] ,
    \sb_1__0__5_chanx_right_out[14] ,
    \sb_1__0__5_chanx_right_out[15] ,
    \sb_1__0__5_chanx_right_out[16] ,
    \sb_1__0__5_chanx_right_out[17] ,
    \sb_1__0__5_chanx_right_out[18] ,
    \sb_1__0__5_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__6_chanx_left_out[0] ,
    \cbx_1__0__6_chanx_left_out[1] ,
    \cbx_1__0__6_chanx_left_out[2] ,
    \cbx_1__0__6_chanx_left_out[3] ,
    \cbx_1__0__6_chanx_left_out[4] ,
    \cbx_1__0__6_chanx_left_out[5] ,
    \cbx_1__0__6_chanx_left_out[6] ,
    \cbx_1__0__6_chanx_left_out[7] ,
    \cbx_1__0__6_chanx_left_out[8] ,
    \cbx_1__0__6_chanx_left_out[9] ,
    \cbx_1__0__6_chanx_left_out[10] ,
    \cbx_1__0__6_chanx_left_out[11] ,
    \cbx_1__0__6_chanx_left_out[12] ,
    \cbx_1__0__6_chanx_left_out[13] ,
    \cbx_1__0__6_chanx_left_out[14] ,
    \cbx_1__0__6_chanx_left_out[15] ,
    \cbx_1__0__6_chanx_left_out[16] ,
    \cbx_1__0__6_chanx_left_out[17] ,
    \cbx_1__0__6_chanx_left_out[18] ,
    \cbx_1__0__6_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__0__6_chanx_left_out[0] ,
    \sb_1__0__6_chanx_left_out[1] ,
    \sb_1__0__6_chanx_left_out[2] ,
    \sb_1__0__6_chanx_left_out[3] ,
    \sb_1__0__6_chanx_left_out[4] ,
    \sb_1__0__6_chanx_left_out[5] ,
    \sb_1__0__6_chanx_left_out[6] ,
    \sb_1__0__6_chanx_left_out[7] ,
    \sb_1__0__6_chanx_left_out[8] ,
    \sb_1__0__6_chanx_left_out[9] ,
    \sb_1__0__6_chanx_left_out[10] ,
    \sb_1__0__6_chanx_left_out[11] ,
    \sb_1__0__6_chanx_left_out[12] ,
    \sb_1__0__6_chanx_left_out[13] ,
    \sb_1__0__6_chanx_left_out[14] ,
    \sb_1__0__6_chanx_left_out[15] ,
    \sb_1__0__6_chanx_left_out[16] ,
    \sb_1__0__6_chanx_left_out[17] ,
    \sb_1__0__6_chanx_left_out[18] ,
    \sb_1__0__6_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__6_chanx_right_out[0] ,
    \cbx_1__0__6_chanx_right_out[1] ,
    \cbx_1__0__6_chanx_right_out[2] ,
    \cbx_1__0__6_chanx_right_out[3] ,
    \cbx_1__0__6_chanx_right_out[4] ,
    \cbx_1__0__6_chanx_right_out[5] ,
    \cbx_1__0__6_chanx_right_out[6] ,
    \cbx_1__0__6_chanx_right_out[7] ,
    \cbx_1__0__6_chanx_right_out[8] ,
    \cbx_1__0__6_chanx_right_out[9] ,
    \cbx_1__0__6_chanx_right_out[10] ,
    \cbx_1__0__6_chanx_right_out[11] ,
    \cbx_1__0__6_chanx_right_out[12] ,
    \cbx_1__0__6_chanx_right_out[13] ,
    \cbx_1__0__6_chanx_right_out[14] ,
    \cbx_1__0__6_chanx_right_out[15] ,
    \cbx_1__0__6_chanx_right_out[16] ,
    \cbx_1__0__6_chanx_right_out[17] ,
    \cbx_1__0__6_chanx_right_out[18] ,
    \cbx_1__0__6_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]}));
 cbx_1__1_ cbx_7__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[42] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[42] ),
    .SC_IN_TOP(\scff_Wires[125] ),
    .SC_OUT_BOT(\scff_Wires[126] ),
    .bottom_grid_pin_0_(cbx_1__1__42_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__42_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__42_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__42_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__42_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__42_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__42_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__42_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__42_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__42_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__42_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__42_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__42_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__42_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__42_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__42_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__42_ccff_tail),
    .ccff_tail(cbx_1__1__42_ccff_tail),
    .clk_1_N_out(\clk_1_wires[87] ),
    .clk_1_S_out(\clk_1_wires[88] ),
    .clk_1_W_in(\clk_1_wires[86] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[176] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[87] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[88] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[86] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__35_chanx_right_out[0] ,
    \sb_1__1__35_chanx_right_out[1] ,
    \sb_1__1__35_chanx_right_out[2] ,
    \sb_1__1__35_chanx_right_out[3] ,
    \sb_1__1__35_chanx_right_out[4] ,
    \sb_1__1__35_chanx_right_out[5] ,
    \sb_1__1__35_chanx_right_out[6] ,
    \sb_1__1__35_chanx_right_out[7] ,
    \sb_1__1__35_chanx_right_out[8] ,
    \sb_1__1__35_chanx_right_out[9] ,
    \sb_1__1__35_chanx_right_out[10] ,
    \sb_1__1__35_chanx_right_out[11] ,
    \sb_1__1__35_chanx_right_out[12] ,
    \sb_1__1__35_chanx_right_out[13] ,
    \sb_1__1__35_chanx_right_out[14] ,
    \sb_1__1__35_chanx_right_out[15] ,
    \sb_1__1__35_chanx_right_out[16] ,
    \sb_1__1__35_chanx_right_out[17] ,
    \sb_1__1__35_chanx_right_out[18] ,
    \sb_1__1__35_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__42_chanx_left_out[0] ,
    \cbx_1__1__42_chanx_left_out[1] ,
    \cbx_1__1__42_chanx_left_out[2] ,
    \cbx_1__1__42_chanx_left_out[3] ,
    \cbx_1__1__42_chanx_left_out[4] ,
    \cbx_1__1__42_chanx_left_out[5] ,
    \cbx_1__1__42_chanx_left_out[6] ,
    \cbx_1__1__42_chanx_left_out[7] ,
    \cbx_1__1__42_chanx_left_out[8] ,
    \cbx_1__1__42_chanx_left_out[9] ,
    \cbx_1__1__42_chanx_left_out[10] ,
    \cbx_1__1__42_chanx_left_out[11] ,
    \cbx_1__1__42_chanx_left_out[12] ,
    \cbx_1__1__42_chanx_left_out[13] ,
    \cbx_1__1__42_chanx_left_out[14] ,
    \cbx_1__1__42_chanx_left_out[15] ,
    \cbx_1__1__42_chanx_left_out[16] ,
    \cbx_1__1__42_chanx_left_out[17] ,
    \cbx_1__1__42_chanx_left_out[18] ,
    \cbx_1__1__42_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__42_chanx_left_out[0] ,
    \sb_1__1__42_chanx_left_out[1] ,
    \sb_1__1__42_chanx_left_out[2] ,
    \sb_1__1__42_chanx_left_out[3] ,
    \sb_1__1__42_chanx_left_out[4] ,
    \sb_1__1__42_chanx_left_out[5] ,
    \sb_1__1__42_chanx_left_out[6] ,
    \sb_1__1__42_chanx_left_out[7] ,
    \sb_1__1__42_chanx_left_out[8] ,
    \sb_1__1__42_chanx_left_out[9] ,
    \sb_1__1__42_chanx_left_out[10] ,
    \sb_1__1__42_chanx_left_out[11] ,
    \sb_1__1__42_chanx_left_out[12] ,
    \sb_1__1__42_chanx_left_out[13] ,
    \sb_1__1__42_chanx_left_out[14] ,
    \sb_1__1__42_chanx_left_out[15] ,
    \sb_1__1__42_chanx_left_out[16] ,
    \sb_1__1__42_chanx_left_out[17] ,
    \sb_1__1__42_chanx_left_out[18] ,
    \sb_1__1__42_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__42_chanx_right_out[0] ,
    \cbx_1__1__42_chanx_right_out[1] ,
    \cbx_1__1__42_chanx_right_out[2] ,
    \cbx_1__1__42_chanx_right_out[3] ,
    \cbx_1__1__42_chanx_right_out[4] ,
    \cbx_1__1__42_chanx_right_out[5] ,
    \cbx_1__1__42_chanx_right_out[6] ,
    \cbx_1__1__42_chanx_right_out[7] ,
    \cbx_1__1__42_chanx_right_out[8] ,
    \cbx_1__1__42_chanx_right_out[9] ,
    \cbx_1__1__42_chanx_right_out[10] ,
    \cbx_1__1__42_chanx_right_out[11] ,
    \cbx_1__1__42_chanx_right_out[12] ,
    \cbx_1__1__42_chanx_right_out[13] ,
    \cbx_1__1__42_chanx_right_out[14] ,
    \cbx_1__1__42_chanx_right_out[15] ,
    \cbx_1__1__42_chanx_right_out[16] ,
    \cbx_1__1__42_chanx_right_out[17] ,
    \cbx_1__1__42_chanx_right_out[18] ,
    \cbx_1__1__42_chanx_right_out[19] }));
 cbx_1__1_ cbx_7__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[43] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[43] ),
    .SC_IN_TOP(\scff_Wires[123] ),
    .SC_OUT_BOT(\scff_Wires[124] ),
    .bottom_grid_pin_0_(cbx_1__1__43_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__43_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__43_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__43_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__43_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__43_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__43_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__43_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__43_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__43_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__43_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__43_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__43_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__43_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__43_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__43_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__43_ccff_tail),
    .ccff_tail(cbx_1__1__43_ccff_tail),
    .clk_2_E_out(\clk_2_wires[28] ),
    .clk_2_W_in(\clk_2_wires[27] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[179] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[28] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[27] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__36_chanx_right_out[0] ,
    \sb_1__1__36_chanx_right_out[1] ,
    \sb_1__1__36_chanx_right_out[2] ,
    \sb_1__1__36_chanx_right_out[3] ,
    \sb_1__1__36_chanx_right_out[4] ,
    \sb_1__1__36_chanx_right_out[5] ,
    \sb_1__1__36_chanx_right_out[6] ,
    \sb_1__1__36_chanx_right_out[7] ,
    \sb_1__1__36_chanx_right_out[8] ,
    \sb_1__1__36_chanx_right_out[9] ,
    \sb_1__1__36_chanx_right_out[10] ,
    \sb_1__1__36_chanx_right_out[11] ,
    \sb_1__1__36_chanx_right_out[12] ,
    \sb_1__1__36_chanx_right_out[13] ,
    \sb_1__1__36_chanx_right_out[14] ,
    \sb_1__1__36_chanx_right_out[15] ,
    \sb_1__1__36_chanx_right_out[16] ,
    \sb_1__1__36_chanx_right_out[17] ,
    \sb_1__1__36_chanx_right_out[18] ,
    \sb_1__1__36_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__43_chanx_left_out[0] ,
    \cbx_1__1__43_chanx_left_out[1] ,
    \cbx_1__1__43_chanx_left_out[2] ,
    \cbx_1__1__43_chanx_left_out[3] ,
    \cbx_1__1__43_chanx_left_out[4] ,
    \cbx_1__1__43_chanx_left_out[5] ,
    \cbx_1__1__43_chanx_left_out[6] ,
    \cbx_1__1__43_chanx_left_out[7] ,
    \cbx_1__1__43_chanx_left_out[8] ,
    \cbx_1__1__43_chanx_left_out[9] ,
    \cbx_1__1__43_chanx_left_out[10] ,
    \cbx_1__1__43_chanx_left_out[11] ,
    \cbx_1__1__43_chanx_left_out[12] ,
    \cbx_1__1__43_chanx_left_out[13] ,
    \cbx_1__1__43_chanx_left_out[14] ,
    \cbx_1__1__43_chanx_left_out[15] ,
    \cbx_1__1__43_chanx_left_out[16] ,
    \cbx_1__1__43_chanx_left_out[17] ,
    \cbx_1__1__43_chanx_left_out[18] ,
    \cbx_1__1__43_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__43_chanx_left_out[0] ,
    \sb_1__1__43_chanx_left_out[1] ,
    \sb_1__1__43_chanx_left_out[2] ,
    \sb_1__1__43_chanx_left_out[3] ,
    \sb_1__1__43_chanx_left_out[4] ,
    \sb_1__1__43_chanx_left_out[5] ,
    \sb_1__1__43_chanx_left_out[6] ,
    \sb_1__1__43_chanx_left_out[7] ,
    \sb_1__1__43_chanx_left_out[8] ,
    \sb_1__1__43_chanx_left_out[9] ,
    \sb_1__1__43_chanx_left_out[10] ,
    \sb_1__1__43_chanx_left_out[11] ,
    \sb_1__1__43_chanx_left_out[12] ,
    \sb_1__1__43_chanx_left_out[13] ,
    \sb_1__1__43_chanx_left_out[14] ,
    \sb_1__1__43_chanx_left_out[15] ,
    \sb_1__1__43_chanx_left_out[16] ,
    \sb_1__1__43_chanx_left_out[17] ,
    \sb_1__1__43_chanx_left_out[18] ,
    \sb_1__1__43_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__43_chanx_right_out[0] ,
    \cbx_1__1__43_chanx_right_out[1] ,
    \cbx_1__1__43_chanx_right_out[2] ,
    \cbx_1__1__43_chanx_right_out[3] ,
    \cbx_1__1__43_chanx_right_out[4] ,
    \cbx_1__1__43_chanx_right_out[5] ,
    \cbx_1__1__43_chanx_right_out[6] ,
    \cbx_1__1__43_chanx_right_out[7] ,
    \cbx_1__1__43_chanx_right_out[8] ,
    \cbx_1__1__43_chanx_right_out[9] ,
    \cbx_1__1__43_chanx_right_out[10] ,
    \cbx_1__1__43_chanx_right_out[11] ,
    \cbx_1__1__43_chanx_right_out[12] ,
    \cbx_1__1__43_chanx_right_out[13] ,
    \cbx_1__1__43_chanx_right_out[14] ,
    \cbx_1__1__43_chanx_right_out[15] ,
    \cbx_1__1__43_chanx_right_out[16] ,
    \cbx_1__1__43_chanx_right_out[17] ,
    \cbx_1__1__43_chanx_right_out[18] ,
    \cbx_1__1__43_chanx_right_out[19] }));
 cbx_1__1_ cbx_7__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[44] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[44] ),
    .SC_IN_TOP(\scff_Wires[121] ),
    .SC_OUT_BOT(\scff_Wires[122] ),
    .bottom_grid_pin_0_(cbx_1__1__44_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__44_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__44_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__44_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__44_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__44_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__44_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__44_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__44_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__44_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__44_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__44_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__44_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__44_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__44_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__44_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__44_ccff_tail),
    .ccff_tail(cbx_1__1__44_ccff_tail),
    .clk_1_N_out(\clk_1_wires[94] ),
    .clk_1_S_out(\clk_1_wires[95] ),
    .clk_1_W_in(\clk_1_wires[93] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[182] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[94] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[95] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[93] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__37_chanx_right_out[0] ,
    \sb_1__1__37_chanx_right_out[1] ,
    \sb_1__1__37_chanx_right_out[2] ,
    \sb_1__1__37_chanx_right_out[3] ,
    \sb_1__1__37_chanx_right_out[4] ,
    \sb_1__1__37_chanx_right_out[5] ,
    \sb_1__1__37_chanx_right_out[6] ,
    \sb_1__1__37_chanx_right_out[7] ,
    \sb_1__1__37_chanx_right_out[8] ,
    \sb_1__1__37_chanx_right_out[9] ,
    \sb_1__1__37_chanx_right_out[10] ,
    \sb_1__1__37_chanx_right_out[11] ,
    \sb_1__1__37_chanx_right_out[12] ,
    \sb_1__1__37_chanx_right_out[13] ,
    \sb_1__1__37_chanx_right_out[14] ,
    \sb_1__1__37_chanx_right_out[15] ,
    \sb_1__1__37_chanx_right_out[16] ,
    \sb_1__1__37_chanx_right_out[17] ,
    \sb_1__1__37_chanx_right_out[18] ,
    \sb_1__1__37_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__44_chanx_left_out[0] ,
    \cbx_1__1__44_chanx_left_out[1] ,
    \cbx_1__1__44_chanx_left_out[2] ,
    \cbx_1__1__44_chanx_left_out[3] ,
    \cbx_1__1__44_chanx_left_out[4] ,
    \cbx_1__1__44_chanx_left_out[5] ,
    \cbx_1__1__44_chanx_left_out[6] ,
    \cbx_1__1__44_chanx_left_out[7] ,
    \cbx_1__1__44_chanx_left_out[8] ,
    \cbx_1__1__44_chanx_left_out[9] ,
    \cbx_1__1__44_chanx_left_out[10] ,
    \cbx_1__1__44_chanx_left_out[11] ,
    \cbx_1__1__44_chanx_left_out[12] ,
    \cbx_1__1__44_chanx_left_out[13] ,
    \cbx_1__1__44_chanx_left_out[14] ,
    \cbx_1__1__44_chanx_left_out[15] ,
    \cbx_1__1__44_chanx_left_out[16] ,
    \cbx_1__1__44_chanx_left_out[17] ,
    \cbx_1__1__44_chanx_left_out[18] ,
    \cbx_1__1__44_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__44_chanx_left_out[0] ,
    \sb_1__1__44_chanx_left_out[1] ,
    \sb_1__1__44_chanx_left_out[2] ,
    \sb_1__1__44_chanx_left_out[3] ,
    \sb_1__1__44_chanx_left_out[4] ,
    \sb_1__1__44_chanx_left_out[5] ,
    \sb_1__1__44_chanx_left_out[6] ,
    \sb_1__1__44_chanx_left_out[7] ,
    \sb_1__1__44_chanx_left_out[8] ,
    \sb_1__1__44_chanx_left_out[9] ,
    \sb_1__1__44_chanx_left_out[10] ,
    \sb_1__1__44_chanx_left_out[11] ,
    \sb_1__1__44_chanx_left_out[12] ,
    \sb_1__1__44_chanx_left_out[13] ,
    \sb_1__1__44_chanx_left_out[14] ,
    \sb_1__1__44_chanx_left_out[15] ,
    \sb_1__1__44_chanx_left_out[16] ,
    \sb_1__1__44_chanx_left_out[17] ,
    \sb_1__1__44_chanx_left_out[18] ,
    \sb_1__1__44_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__44_chanx_right_out[0] ,
    \cbx_1__1__44_chanx_right_out[1] ,
    \cbx_1__1__44_chanx_right_out[2] ,
    \cbx_1__1__44_chanx_right_out[3] ,
    \cbx_1__1__44_chanx_right_out[4] ,
    \cbx_1__1__44_chanx_right_out[5] ,
    \cbx_1__1__44_chanx_right_out[6] ,
    \cbx_1__1__44_chanx_right_out[7] ,
    \cbx_1__1__44_chanx_right_out[8] ,
    \cbx_1__1__44_chanx_right_out[9] ,
    \cbx_1__1__44_chanx_right_out[10] ,
    \cbx_1__1__44_chanx_right_out[11] ,
    \cbx_1__1__44_chanx_right_out[12] ,
    \cbx_1__1__44_chanx_right_out[13] ,
    \cbx_1__1__44_chanx_right_out[14] ,
    \cbx_1__1__44_chanx_right_out[15] ,
    \cbx_1__1__44_chanx_right_out[16] ,
    \cbx_1__1__44_chanx_right_out[17] ,
    \cbx_1__1__44_chanx_right_out[18] ,
    \cbx_1__1__44_chanx_right_out[19] }));
 cbx_1__1_ cbx_7__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[45] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[45] ),
    .SC_IN_TOP(\scff_Wires[119] ),
    .SC_OUT_BOT(\scff_Wires[120] ),
    .bottom_grid_pin_0_(cbx_1__1__45_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__45_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__45_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__45_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__45_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__45_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__45_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__45_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__45_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__45_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__45_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__45_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__45_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__45_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__45_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__45_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__45_ccff_tail),
    .ccff_tail(cbx_1__1__45_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[185] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__38_chanx_right_out[0] ,
    \sb_1__1__38_chanx_right_out[1] ,
    \sb_1__1__38_chanx_right_out[2] ,
    \sb_1__1__38_chanx_right_out[3] ,
    \sb_1__1__38_chanx_right_out[4] ,
    \sb_1__1__38_chanx_right_out[5] ,
    \sb_1__1__38_chanx_right_out[6] ,
    \sb_1__1__38_chanx_right_out[7] ,
    \sb_1__1__38_chanx_right_out[8] ,
    \sb_1__1__38_chanx_right_out[9] ,
    \sb_1__1__38_chanx_right_out[10] ,
    \sb_1__1__38_chanx_right_out[11] ,
    \sb_1__1__38_chanx_right_out[12] ,
    \sb_1__1__38_chanx_right_out[13] ,
    \sb_1__1__38_chanx_right_out[14] ,
    \sb_1__1__38_chanx_right_out[15] ,
    \sb_1__1__38_chanx_right_out[16] ,
    \sb_1__1__38_chanx_right_out[17] ,
    \sb_1__1__38_chanx_right_out[18] ,
    \sb_1__1__38_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__45_chanx_left_out[0] ,
    \cbx_1__1__45_chanx_left_out[1] ,
    \cbx_1__1__45_chanx_left_out[2] ,
    \cbx_1__1__45_chanx_left_out[3] ,
    \cbx_1__1__45_chanx_left_out[4] ,
    \cbx_1__1__45_chanx_left_out[5] ,
    \cbx_1__1__45_chanx_left_out[6] ,
    \cbx_1__1__45_chanx_left_out[7] ,
    \cbx_1__1__45_chanx_left_out[8] ,
    \cbx_1__1__45_chanx_left_out[9] ,
    \cbx_1__1__45_chanx_left_out[10] ,
    \cbx_1__1__45_chanx_left_out[11] ,
    \cbx_1__1__45_chanx_left_out[12] ,
    \cbx_1__1__45_chanx_left_out[13] ,
    \cbx_1__1__45_chanx_left_out[14] ,
    \cbx_1__1__45_chanx_left_out[15] ,
    \cbx_1__1__45_chanx_left_out[16] ,
    \cbx_1__1__45_chanx_left_out[17] ,
    \cbx_1__1__45_chanx_left_out[18] ,
    \cbx_1__1__45_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__45_chanx_left_out[0] ,
    \sb_1__1__45_chanx_left_out[1] ,
    \sb_1__1__45_chanx_left_out[2] ,
    \sb_1__1__45_chanx_left_out[3] ,
    \sb_1__1__45_chanx_left_out[4] ,
    \sb_1__1__45_chanx_left_out[5] ,
    \sb_1__1__45_chanx_left_out[6] ,
    \sb_1__1__45_chanx_left_out[7] ,
    \sb_1__1__45_chanx_left_out[8] ,
    \sb_1__1__45_chanx_left_out[9] ,
    \sb_1__1__45_chanx_left_out[10] ,
    \sb_1__1__45_chanx_left_out[11] ,
    \sb_1__1__45_chanx_left_out[12] ,
    \sb_1__1__45_chanx_left_out[13] ,
    \sb_1__1__45_chanx_left_out[14] ,
    \sb_1__1__45_chanx_left_out[15] ,
    \sb_1__1__45_chanx_left_out[16] ,
    \sb_1__1__45_chanx_left_out[17] ,
    \sb_1__1__45_chanx_left_out[18] ,
    \sb_1__1__45_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__45_chanx_right_out[0] ,
    \cbx_1__1__45_chanx_right_out[1] ,
    \cbx_1__1__45_chanx_right_out[2] ,
    \cbx_1__1__45_chanx_right_out[3] ,
    \cbx_1__1__45_chanx_right_out[4] ,
    \cbx_1__1__45_chanx_right_out[5] ,
    \cbx_1__1__45_chanx_right_out[6] ,
    \cbx_1__1__45_chanx_right_out[7] ,
    \cbx_1__1__45_chanx_right_out[8] ,
    \cbx_1__1__45_chanx_right_out[9] ,
    \cbx_1__1__45_chanx_right_out[10] ,
    \cbx_1__1__45_chanx_right_out[11] ,
    \cbx_1__1__45_chanx_right_out[12] ,
    \cbx_1__1__45_chanx_right_out[13] ,
    \cbx_1__1__45_chanx_right_out[14] ,
    \cbx_1__1__45_chanx_right_out[15] ,
    \cbx_1__1__45_chanx_right_out[16] ,
    \cbx_1__1__45_chanx_right_out[17] ,
    \cbx_1__1__45_chanx_right_out[18] ,
    \cbx_1__1__45_chanx_right_out[19] }));
 cbx_1__1_ cbx_7__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[46] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[46] ),
    .SC_IN_TOP(\scff_Wires[117] ),
    .SC_OUT_BOT(\scff_Wires[118] ),
    .bottom_grid_pin_0_(cbx_1__1__46_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__46_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__46_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__46_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__46_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__46_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__46_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__46_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__46_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__46_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__46_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__46_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__46_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__46_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__46_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__46_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__46_ccff_tail),
    .ccff_tail(cbx_1__1__46_ccff_tail),
    .clk_1_N_out(\clk_1_wires[101] ),
    .clk_1_S_out(\clk_1_wires[102] ),
    .clk_1_W_in(\clk_1_wires[100] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[188] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[101] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[102] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[100] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__39_chanx_right_out[0] ,
    \sb_1__1__39_chanx_right_out[1] ,
    \sb_1__1__39_chanx_right_out[2] ,
    \sb_1__1__39_chanx_right_out[3] ,
    \sb_1__1__39_chanx_right_out[4] ,
    \sb_1__1__39_chanx_right_out[5] ,
    \sb_1__1__39_chanx_right_out[6] ,
    \sb_1__1__39_chanx_right_out[7] ,
    \sb_1__1__39_chanx_right_out[8] ,
    \sb_1__1__39_chanx_right_out[9] ,
    \sb_1__1__39_chanx_right_out[10] ,
    \sb_1__1__39_chanx_right_out[11] ,
    \sb_1__1__39_chanx_right_out[12] ,
    \sb_1__1__39_chanx_right_out[13] ,
    \sb_1__1__39_chanx_right_out[14] ,
    \sb_1__1__39_chanx_right_out[15] ,
    \sb_1__1__39_chanx_right_out[16] ,
    \sb_1__1__39_chanx_right_out[17] ,
    \sb_1__1__39_chanx_right_out[18] ,
    \sb_1__1__39_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__46_chanx_left_out[0] ,
    \cbx_1__1__46_chanx_left_out[1] ,
    \cbx_1__1__46_chanx_left_out[2] ,
    \cbx_1__1__46_chanx_left_out[3] ,
    \cbx_1__1__46_chanx_left_out[4] ,
    \cbx_1__1__46_chanx_left_out[5] ,
    \cbx_1__1__46_chanx_left_out[6] ,
    \cbx_1__1__46_chanx_left_out[7] ,
    \cbx_1__1__46_chanx_left_out[8] ,
    \cbx_1__1__46_chanx_left_out[9] ,
    \cbx_1__1__46_chanx_left_out[10] ,
    \cbx_1__1__46_chanx_left_out[11] ,
    \cbx_1__1__46_chanx_left_out[12] ,
    \cbx_1__1__46_chanx_left_out[13] ,
    \cbx_1__1__46_chanx_left_out[14] ,
    \cbx_1__1__46_chanx_left_out[15] ,
    \cbx_1__1__46_chanx_left_out[16] ,
    \cbx_1__1__46_chanx_left_out[17] ,
    \cbx_1__1__46_chanx_left_out[18] ,
    \cbx_1__1__46_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__46_chanx_left_out[0] ,
    \sb_1__1__46_chanx_left_out[1] ,
    \sb_1__1__46_chanx_left_out[2] ,
    \sb_1__1__46_chanx_left_out[3] ,
    \sb_1__1__46_chanx_left_out[4] ,
    \sb_1__1__46_chanx_left_out[5] ,
    \sb_1__1__46_chanx_left_out[6] ,
    \sb_1__1__46_chanx_left_out[7] ,
    \sb_1__1__46_chanx_left_out[8] ,
    \sb_1__1__46_chanx_left_out[9] ,
    \sb_1__1__46_chanx_left_out[10] ,
    \sb_1__1__46_chanx_left_out[11] ,
    \sb_1__1__46_chanx_left_out[12] ,
    \sb_1__1__46_chanx_left_out[13] ,
    \sb_1__1__46_chanx_left_out[14] ,
    \sb_1__1__46_chanx_left_out[15] ,
    \sb_1__1__46_chanx_left_out[16] ,
    \sb_1__1__46_chanx_left_out[17] ,
    \sb_1__1__46_chanx_left_out[18] ,
    \sb_1__1__46_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__46_chanx_right_out[0] ,
    \cbx_1__1__46_chanx_right_out[1] ,
    \cbx_1__1__46_chanx_right_out[2] ,
    \cbx_1__1__46_chanx_right_out[3] ,
    \cbx_1__1__46_chanx_right_out[4] ,
    \cbx_1__1__46_chanx_right_out[5] ,
    \cbx_1__1__46_chanx_right_out[6] ,
    \cbx_1__1__46_chanx_right_out[7] ,
    \cbx_1__1__46_chanx_right_out[8] ,
    \cbx_1__1__46_chanx_right_out[9] ,
    \cbx_1__1__46_chanx_right_out[10] ,
    \cbx_1__1__46_chanx_right_out[11] ,
    \cbx_1__1__46_chanx_right_out[12] ,
    \cbx_1__1__46_chanx_right_out[13] ,
    \cbx_1__1__46_chanx_right_out[14] ,
    \cbx_1__1__46_chanx_right_out[15] ,
    \cbx_1__1__46_chanx_right_out[16] ,
    \cbx_1__1__46_chanx_right_out[17] ,
    \cbx_1__1__46_chanx_right_out[18] ,
    \cbx_1__1__46_chanx_right_out[19] }));
 cbx_1__1_ cbx_7__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[47] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[47] ),
    .SC_IN_TOP(\scff_Wires[115] ),
    .SC_OUT_BOT(\scff_Wires[116] ),
    .bottom_grid_pin_0_(cbx_1__1__47_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__47_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__47_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__47_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__47_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__47_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__47_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__47_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__47_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__47_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__47_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__47_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__47_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__47_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__47_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__47_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__47_ccff_tail),
    .ccff_tail(cbx_1__1__47_ccff_tail),
    .clk_2_E_out(\clk_2_wires[41] ),
    .clk_2_W_in(\clk_2_wires[40] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[191] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[41] ),
    .prog_clk_2_W_in(\prog_clk_2_wires[40] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__40_chanx_right_out[0] ,
    \sb_1__1__40_chanx_right_out[1] ,
    \sb_1__1__40_chanx_right_out[2] ,
    \sb_1__1__40_chanx_right_out[3] ,
    \sb_1__1__40_chanx_right_out[4] ,
    \sb_1__1__40_chanx_right_out[5] ,
    \sb_1__1__40_chanx_right_out[6] ,
    \sb_1__1__40_chanx_right_out[7] ,
    \sb_1__1__40_chanx_right_out[8] ,
    \sb_1__1__40_chanx_right_out[9] ,
    \sb_1__1__40_chanx_right_out[10] ,
    \sb_1__1__40_chanx_right_out[11] ,
    \sb_1__1__40_chanx_right_out[12] ,
    \sb_1__1__40_chanx_right_out[13] ,
    \sb_1__1__40_chanx_right_out[14] ,
    \sb_1__1__40_chanx_right_out[15] ,
    \sb_1__1__40_chanx_right_out[16] ,
    \sb_1__1__40_chanx_right_out[17] ,
    \sb_1__1__40_chanx_right_out[18] ,
    \sb_1__1__40_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__47_chanx_left_out[0] ,
    \cbx_1__1__47_chanx_left_out[1] ,
    \cbx_1__1__47_chanx_left_out[2] ,
    \cbx_1__1__47_chanx_left_out[3] ,
    \cbx_1__1__47_chanx_left_out[4] ,
    \cbx_1__1__47_chanx_left_out[5] ,
    \cbx_1__1__47_chanx_left_out[6] ,
    \cbx_1__1__47_chanx_left_out[7] ,
    \cbx_1__1__47_chanx_left_out[8] ,
    \cbx_1__1__47_chanx_left_out[9] ,
    \cbx_1__1__47_chanx_left_out[10] ,
    \cbx_1__1__47_chanx_left_out[11] ,
    \cbx_1__1__47_chanx_left_out[12] ,
    \cbx_1__1__47_chanx_left_out[13] ,
    \cbx_1__1__47_chanx_left_out[14] ,
    \cbx_1__1__47_chanx_left_out[15] ,
    \cbx_1__1__47_chanx_left_out[16] ,
    \cbx_1__1__47_chanx_left_out[17] ,
    \cbx_1__1__47_chanx_left_out[18] ,
    \cbx_1__1__47_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__47_chanx_left_out[0] ,
    \sb_1__1__47_chanx_left_out[1] ,
    \sb_1__1__47_chanx_left_out[2] ,
    \sb_1__1__47_chanx_left_out[3] ,
    \sb_1__1__47_chanx_left_out[4] ,
    \sb_1__1__47_chanx_left_out[5] ,
    \sb_1__1__47_chanx_left_out[6] ,
    \sb_1__1__47_chanx_left_out[7] ,
    \sb_1__1__47_chanx_left_out[8] ,
    \sb_1__1__47_chanx_left_out[9] ,
    \sb_1__1__47_chanx_left_out[10] ,
    \sb_1__1__47_chanx_left_out[11] ,
    \sb_1__1__47_chanx_left_out[12] ,
    \sb_1__1__47_chanx_left_out[13] ,
    \sb_1__1__47_chanx_left_out[14] ,
    \sb_1__1__47_chanx_left_out[15] ,
    \sb_1__1__47_chanx_left_out[16] ,
    \sb_1__1__47_chanx_left_out[17] ,
    \sb_1__1__47_chanx_left_out[18] ,
    \sb_1__1__47_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__47_chanx_right_out[0] ,
    \cbx_1__1__47_chanx_right_out[1] ,
    \cbx_1__1__47_chanx_right_out[2] ,
    \cbx_1__1__47_chanx_right_out[3] ,
    \cbx_1__1__47_chanx_right_out[4] ,
    \cbx_1__1__47_chanx_right_out[5] ,
    \cbx_1__1__47_chanx_right_out[6] ,
    \cbx_1__1__47_chanx_right_out[7] ,
    \cbx_1__1__47_chanx_right_out[8] ,
    \cbx_1__1__47_chanx_right_out[9] ,
    \cbx_1__1__47_chanx_right_out[10] ,
    \cbx_1__1__47_chanx_right_out[11] ,
    \cbx_1__1__47_chanx_right_out[12] ,
    \cbx_1__1__47_chanx_right_out[13] ,
    \cbx_1__1__47_chanx_right_out[14] ,
    \cbx_1__1__47_chanx_right_out[15] ,
    \cbx_1__1__47_chanx_right_out[16] ,
    \cbx_1__1__47_chanx_right_out[17] ,
    \cbx_1__1__47_chanx_right_out[18] ,
    \cbx_1__1__47_chanx_right_out[19] }));
 cbx_1__1_ cbx_7__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[48] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[48] ),
    .SC_IN_TOP(\scff_Wires[113] ),
    .SC_OUT_BOT(\scff_Wires[114] ),
    .bottom_grid_pin_0_(cbx_1__1__48_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__48_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__48_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__48_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__48_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__48_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__48_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__48_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__48_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__48_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__48_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__48_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__48_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__48_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__48_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__48_bottom_grid_pin_9_),
    .ccff_head(sb_1__1__48_ccff_tail),
    .ccff_tail(cbx_1__1__48_ccff_tail),
    .clk_1_N_out(\clk_1_wires[108] ),
    .clk_1_S_out(\clk_1_wires[109] ),
    .clk_1_W_in(\clk_1_wires[107] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[194] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[108] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[109] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[107] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__41_chanx_right_out[0] ,
    \sb_1__1__41_chanx_right_out[1] ,
    \sb_1__1__41_chanx_right_out[2] ,
    \sb_1__1__41_chanx_right_out[3] ,
    \sb_1__1__41_chanx_right_out[4] ,
    \sb_1__1__41_chanx_right_out[5] ,
    \sb_1__1__41_chanx_right_out[6] ,
    \sb_1__1__41_chanx_right_out[7] ,
    \sb_1__1__41_chanx_right_out[8] ,
    \sb_1__1__41_chanx_right_out[9] ,
    \sb_1__1__41_chanx_right_out[10] ,
    \sb_1__1__41_chanx_right_out[11] ,
    \sb_1__1__41_chanx_right_out[12] ,
    \sb_1__1__41_chanx_right_out[13] ,
    \sb_1__1__41_chanx_right_out[14] ,
    \sb_1__1__41_chanx_right_out[15] ,
    \sb_1__1__41_chanx_right_out[16] ,
    \sb_1__1__41_chanx_right_out[17] ,
    \sb_1__1__41_chanx_right_out[18] ,
    \sb_1__1__41_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__48_chanx_left_out[0] ,
    \cbx_1__1__48_chanx_left_out[1] ,
    \cbx_1__1__48_chanx_left_out[2] ,
    \cbx_1__1__48_chanx_left_out[3] ,
    \cbx_1__1__48_chanx_left_out[4] ,
    \cbx_1__1__48_chanx_left_out[5] ,
    \cbx_1__1__48_chanx_left_out[6] ,
    \cbx_1__1__48_chanx_left_out[7] ,
    \cbx_1__1__48_chanx_left_out[8] ,
    \cbx_1__1__48_chanx_left_out[9] ,
    \cbx_1__1__48_chanx_left_out[10] ,
    \cbx_1__1__48_chanx_left_out[11] ,
    \cbx_1__1__48_chanx_left_out[12] ,
    \cbx_1__1__48_chanx_left_out[13] ,
    \cbx_1__1__48_chanx_left_out[14] ,
    \cbx_1__1__48_chanx_left_out[15] ,
    \cbx_1__1__48_chanx_left_out[16] ,
    \cbx_1__1__48_chanx_left_out[17] ,
    \cbx_1__1__48_chanx_left_out[18] ,
    \cbx_1__1__48_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__1__48_chanx_left_out[0] ,
    \sb_1__1__48_chanx_left_out[1] ,
    \sb_1__1__48_chanx_left_out[2] ,
    \sb_1__1__48_chanx_left_out[3] ,
    \sb_1__1__48_chanx_left_out[4] ,
    \sb_1__1__48_chanx_left_out[5] ,
    \sb_1__1__48_chanx_left_out[6] ,
    \sb_1__1__48_chanx_left_out[7] ,
    \sb_1__1__48_chanx_left_out[8] ,
    \sb_1__1__48_chanx_left_out[9] ,
    \sb_1__1__48_chanx_left_out[10] ,
    \sb_1__1__48_chanx_left_out[11] ,
    \sb_1__1__48_chanx_left_out[12] ,
    \sb_1__1__48_chanx_left_out[13] ,
    \sb_1__1__48_chanx_left_out[14] ,
    \sb_1__1__48_chanx_left_out[15] ,
    \sb_1__1__48_chanx_left_out[16] ,
    \sb_1__1__48_chanx_left_out[17] ,
    \sb_1__1__48_chanx_left_out[18] ,
    \sb_1__1__48_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__48_chanx_right_out[0] ,
    \cbx_1__1__48_chanx_right_out[1] ,
    \cbx_1__1__48_chanx_right_out[2] ,
    \cbx_1__1__48_chanx_right_out[3] ,
    \cbx_1__1__48_chanx_right_out[4] ,
    \cbx_1__1__48_chanx_right_out[5] ,
    \cbx_1__1__48_chanx_right_out[6] ,
    \cbx_1__1__48_chanx_right_out[7] ,
    \cbx_1__1__48_chanx_right_out[8] ,
    \cbx_1__1__48_chanx_right_out[9] ,
    \cbx_1__1__48_chanx_right_out[10] ,
    \cbx_1__1__48_chanx_right_out[11] ,
    \cbx_1__1__48_chanx_right_out[12] ,
    \cbx_1__1__48_chanx_right_out[13] ,
    \cbx_1__1__48_chanx_right_out[14] ,
    \cbx_1__1__48_chanx_right_out[15] ,
    \cbx_1__1__48_chanx_right_out[16] ,
    \cbx_1__1__48_chanx_right_out[17] ,
    \cbx_1__1__48_chanx_right_out[18] ,
    \cbx_1__1__48_chanx_right_out[19] }));
 cbx_1__2_ cbx_7__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_TOP(\scff_Wires[111] ),
    .SC_OUT_BOT(\scff_Wires[112] ),
    .bottom_grid_pin_0_(cbx_1__8__6_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__6_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__6_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__6_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__6_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__6_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__6_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__6_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__6_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__6_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__6_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__6_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__6_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__6_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__6_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__6_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__6_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_6_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_6_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_1__8__6_ccff_tail),
    .ccff_tail(grid_io_top_6_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]),
    .prog_clk_0_S_in(\prog_clk_0_wires[197] ),
    .top_grid_pin_0_(cbx_1__8__6_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__8__5_chanx_right_out[0] ,
    \sb_1__8__5_chanx_right_out[1] ,
    \sb_1__8__5_chanx_right_out[2] ,
    \sb_1__8__5_chanx_right_out[3] ,
    \sb_1__8__5_chanx_right_out[4] ,
    \sb_1__8__5_chanx_right_out[5] ,
    \sb_1__8__5_chanx_right_out[6] ,
    \sb_1__8__5_chanx_right_out[7] ,
    \sb_1__8__5_chanx_right_out[8] ,
    \sb_1__8__5_chanx_right_out[9] ,
    \sb_1__8__5_chanx_right_out[10] ,
    \sb_1__8__5_chanx_right_out[11] ,
    \sb_1__8__5_chanx_right_out[12] ,
    \sb_1__8__5_chanx_right_out[13] ,
    \sb_1__8__5_chanx_right_out[14] ,
    \sb_1__8__5_chanx_right_out[15] ,
    \sb_1__8__5_chanx_right_out[16] ,
    \sb_1__8__5_chanx_right_out[17] ,
    \sb_1__8__5_chanx_right_out[18] ,
    \sb_1__8__5_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__6_chanx_left_out[0] ,
    \cbx_1__8__6_chanx_left_out[1] ,
    \cbx_1__8__6_chanx_left_out[2] ,
    \cbx_1__8__6_chanx_left_out[3] ,
    \cbx_1__8__6_chanx_left_out[4] ,
    \cbx_1__8__6_chanx_left_out[5] ,
    \cbx_1__8__6_chanx_left_out[6] ,
    \cbx_1__8__6_chanx_left_out[7] ,
    \cbx_1__8__6_chanx_left_out[8] ,
    \cbx_1__8__6_chanx_left_out[9] ,
    \cbx_1__8__6_chanx_left_out[10] ,
    \cbx_1__8__6_chanx_left_out[11] ,
    \cbx_1__8__6_chanx_left_out[12] ,
    \cbx_1__8__6_chanx_left_out[13] ,
    \cbx_1__8__6_chanx_left_out[14] ,
    \cbx_1__8__6_chanx_left_out[15] ,
    \cbx_1__8__6_chanx_left_out[16] ,
    \cbx_1__8__6_chanx_left_out[17] ,
    \cbx_1__8__6_chanx_left_out[18] ,
    \cbx_1__8__6_chanx_left_out[19] }),
    .chanx_right_in({\sb_1__8__6_chanx_left_out[0] ,
    \sb_1__8__6_chanx_left_out[1] ,
    \sb_1__8__6_chanx_left_out[2] ,
    \sb_1__8__6_chanx_left_out[3] ,
    \sb_1__8__6_chanx_left_out[4] ,
    \sb_1__8__6_chanx_left_out[5] ,
    \sb_1__8__6_chanx_left_out[6] ,
    \sb_1__8__6_chanx_left_out[7] ,
    \sb_1__8__6_chanx_left_out[8] ,
    \sb_1__8__6_chanx_left_out[9] ,
    \sb_1__8__6_chanx_left_out[10] ,
    \sb_1__8__6_chanx_left_out[11] ,
    \sb_1__8__6_chanx_left_out[12] ,
    \sb_1__8__6_chanx_left_out[13] ,
    \sb_1__8__6_chanx_left_out[14] ,
    \sb_1__8__6_chanx_left_out[15] ,
    \sb_1__8__6_chanx_left_out[16] ,
    \sb_1__8__6_chanx_left_out[17] ,
    \sb_1__8__6_chanx_left_out[18] ,
    \sb_1__8__6_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__6_chanx_right_out[0] ,
    \cbx_1__8__6_chanx_right_out[1] ,
    \cbx_1__8__6_chanx_right_out[2] ,
    \cbx_1__8__6_chanx_right_out[3] ,
    \cbx_1__8__6_chanx_right_out[4] ,
    \cbx_1__8__6_chanx_right_out[5] ,
    \cbx_1__8__6_chanx_right_out[6] ,
    \cbx_1__8__6_chanx_right_out[7] ,
    \cbx_1__8__6_chanx_right_out[8] ,
    \cbx_1__8__6_chanx_right_out[9] ,
    \cbx_1__8__6_chanx_right_out[10] ,
    \cbx_1__8__6_chanx_right_out[11] ,
    \cbx_1__8__6_chanx_right_out[12] ,
    \cbx_1__8__6_chanx_right_out[13] ,
    \cbx_1__8__6_chanx_right_out[14] ,
    \cbx_1__8__6_chanx_right_out[15] ,
    \cbx_1__8__6_chanx_right_out[16] ,
    \cbx_1__8__6_chanx_right_out[17] ,
    \cbx_1__8__6_chanx_right_out[18] ,
    \cbx_1__8__6_chanx_right_out[19] }));
 cbx_1__0_ cbx_8__0_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[130] ),
    .SC_OUT_TOP(\scff_Wires[131] ),
    .bottom_grid_pin_0_(cbx_1__0__7_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__0__7_bottom_grid_pin_10_),
    .bottom_grid_pin_12_(cbx_1__0__7_bottom_grid_pin_12_),
    .bottom_grid_pin_14_(cbx_1__0__7_bottom_grid_pin_14_),
    .bottom_grid_pin_16_(cbx_1__0__7_bottom_grid_pin_16_),
    .bottom_grid_pin_2_(cbx_1__0__7_bottom_grid_pin_2_),
    .bottom_grid_pin_4_(cbx_1__0__7_bottom_grid_pin_4_),
    .bottom_grid_pin_6_(cbx_1__0__7_bottom_grid_pin_6_),
    .bottom_grid_pin_8_(cbx_1__0__7_bottom_grid_pin_8_),
    .ccff_head(sb_8__0__0_ccff_tail),
    .ccff_tail(grid_io_bottom_0_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[199] ),
    .top_width_0_height_0__pin_0_(cbx_1__0__7_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__0__7_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_0_top_width_0_height_0__pin_11_lower),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_0_top_width_0_height_0__pin_11_upper),
    .top_width_0_height_0__pin_12_(cbx_1__0__7_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_0_top_width_0_height_0__pin_13_lower),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_0_top_width_0_height_0__pin_13_upper),
    .top_width_0_height_0__pin_14_(cbx_1__0__7_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_0_top_width_0_height_0__pin_15_lower),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_0_top_width_0_height_0__pin_15_upper),
    .top_width_0_height_0__pin_16_(cbx_1__0__7_bottom_grid_pin_16_),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_0_top_width_0_height_0__pin_17_lower),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_0_top_width_0_height_0__pin_17_upper),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_0_top_width_0_height_0__pin_1_lower),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_0_top_width_0_height_0__pin_1_upper),
    .top_width_0_height_0__pin_2_(cbx_1__0__7_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_0_top_width_0_height_0__pin_3_lower),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_0_top_width_0_height_0__pin_3_upper),
    .top_width_0_height_0__pin_4_(cbx_1__0__7_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_0_top_width_0_height_0__pin_5_lower),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_0_top_width_0_height_0__pin_5_upper),
    .top_width_0_height_0__pin_6_(cbx_1__0__7_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_0_top_width_0_height_0__pin_7_lower),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_0_top_width_0_height_0__pin_7_upper),
    .top_width_0_height_0__pin_8_(cbx_1__0__7_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_0_top_width_0_height_0__pin_9_lower),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_0_top_width_0_height_0__pin_9_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__0__6_chanx_right_out[0] ,
    \sb_1__0__6_chanx_right_out[1] ,
    \sb_1__0__6_chanx_right_out[2] ,
    \sb_1__0__6_chanx_right_out[3] ,
    \sb_1__0__6_chanx_right_out[4] ,
    \sb_1__0__6_chanx_right_out[5] ,
    \sb_1__0__6_chanx_right_out[6] ,
    \sb_1__0__6_chanx_right_out[7] ,
    \sb_1__0__6_chanx_right_out[8] ,
    \sb_1__0__6_chanx_right_out[9] ,
    \sb_1__0__6_chanx_right_out[10] ,
    \sb_1__0__6_chanx_right_out[11] ,
    \sb_1__0__6_chanx_right_out[12] ,
    \sb_1__0__6_chanx_right_out[13] ,
    \sb_1__0__6_chanx_right_out[14] ,
    \sb_1__0__6_chanx_right_out[15] ,
    \sb_1__0__6_chanx_right_out[16] ,
    \sb_1__0__6_chanx_right_out[17] ,
    \sb_1__0__6_chanx_right_out[18] ,
    \sb_1__0__6_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__0__7_chanx_left_out[0] ,
    \cbx_1__0__7_chanx_left_out[1] ,
    \cbx_1__0__7_chanx_left_out[2] ,
    \cbx_1__0__7_chanx_left_out[3] ,
    \cbx_1__0__7_chanx_left_out[4] ,
    \cbx_1__0__7_chanx_left_out[5] ,
    \cbx_1__0__7_chanx_left_out[6] ,
    \cbx_1__0__7_chanx_left_out[7] ,
    \cbx_1__0__7_chanx_left_out[8] ,
    \cbx_1__0__7_chanx_left_out[9] ,
    \cbx_1__0__7_chanx_left_out[10] ,
    \cbx_1__0__7_chanx_left_out[11] ,
    \cbx_1__0__7_chanx_left_out[12] ,
    \cbx_1__0__7_chanx_left_out[13] ,
    \cbx_1__0__7_chanx_left_out[14] ,
    \cbx_1__0__7_chanx_left_out[15] ,
    \cbx_1__0__7_chanx_left_out[16] ,
    \cbx_1__0__7_chanx_left_out[17] ,
    \cbx_1__0__7_chanx_left_out[18] ,
    \cbx_1__0__7_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__0__0_chanx_left_out[0] ,
    \sb_8__0__0_chanx_left_out[1] ,
    \sb_8__0__0_chanx_left_out[2] ,
    \sb_8__0__0_chanx_left_out[3] ,
    \sb_8__0__0_chanx_left_out[4] ,
    \sb_8__0__0_chanx_left_out[5] ,
    \sb_8__0__0_chanx_left_out[6] ,
    \sb_8__0__0_chanx_left_out[7] ,
    \sb_8__0__0_chanx_left_out[8] ,
    \sb_8__0__0_chanx_left_out[9] ,
    \sb_8__0__0_chanx_left_out[10] ,
    \sb_8__0__0_chanx_left_out[11] ,
    \sb_8__0__0_chanx_left_out[12] ,
    \sb_8__0__0_chanx_left_out[13] ,
    \sb_8__0__0_chanx_left_out[14] ,
    \sb_8__0__0_chanx_left_out[15] ,
    \sb_8__0__0_chanx_left_out[16] ,
    \sb_8__0__0_chanx_left_out[17] ,
    \sb_8__0__0_chanx_left_out[18] ,
    \sb_8__0__0_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__0__7_chanx_right_out[0] ,
    \cbx_1__0__7_chanx_right_out[1] ,
    \cbx_1__0__7_chanx_right_out[2] ,
    \cbx_1__0__7_chanx_right_out[3] ,
    \cbx_1__0__7_chanx_right_out[4] ,
    \cbx_1__0__7_chanx_right_out[5] ,
    \cbx_1__0__7_chanx_right_out[6] ,
    \cbx_1__0__7_chanx_right_out[7] ,
    \cbx_1__0__7_chanx_right_out[8] ,
    \cbx_1__0__7_chanx_right_out[9] ,
    \cbx_1__0__7_chanx_right_out[10] ,
    \cbx_1__0__7_chanx_right_out[11] ,
    \cbx_1__0__7_chanx_right_out[12] ,
    \cbx_1__0__7_chanx_right_out[13] ,
    \cbx_1__0__7_chanx_right_out[14] ,
    \cbx_1__0__7_chanx_right_out[15] ,
    \cbx_1__0__7_chanx_right_out[16] ,
    \cbx_1__0__7_chanx_right_out[17] ,
    \cbx_1__0__7_chanx_right_out[18] ,
    \cbx_1__0__7_chanx_right_out[19] }),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR({gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17],
    gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN({gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17],
    gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]}),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT({gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17],
    gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]}));
 cbx_1__1_ cbx_8__1_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[49] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[49] ),
    .SC_IN_BOT(\scff_Wires[132] ),
    .SC_OUT_TOP(\scff_Wires[133] ),
    .bottom_grid_pin_0_(cbx_1__1__49_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__49_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__49_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__49_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__49_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__49_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__49_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__49_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__49_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__49_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__49_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__49_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__49_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__49_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__49_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__49_bottom_grid_pin_9_),
    .ccff_head(sb_8__1__0_ccff_tail),
    .ccff_tail(cbx_1__1__49_ccff_tail),
    .clk_1_N_out(\clk_1_wires[89] ),
    .clk_1_S_out(\clk_1_wires[90] ),
    .clk_1_W_in(\clk_1_wires[85] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[202] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[89] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[90] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[85] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__42_chanx_right_out[0] ,
    \sb_1__1__42_chanx_right_out[1] ,
    \sb_1__1__42_chanx_right_out[2] ,
    \sb_1__1__42_chanx_right_out[3] ,
    \sb_1__1__42_chanx_right_out[4] ,
    \sb_1__1__42_chanx_right_out[5] ,
    \sb_1__1__42_chanx_right_out[6] ,
    \sb_1__1__42_chanx_right_out[7] ,
    \sb_1__1__42_chanx_right_out[8] ,
    \sb_1__1__42_chanx_right_out[9] ,
    \sb_1__1__42_chanx_right_out[10] ,
    \sb_1__1__42_chanx_right_out[11] ,
    \sb_1__1__42_chanx_right_out[12] ,
    \sb_1__1__42_chanx_right_out[13] ,
    \sb_1__1__42_chanx_right_out[14] ,
    \sb_1__1__42_chanx_right_out[15] ,
    \sb_1__1__42_chanx_right_out[16] ,
    \sb_1__1__42_chanx_right_out[17] ,
    \sb_1__1__42_chanx_right_out[18] ,
    \sb_1__1__42_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__49_chanx_left_out[0] ,
    \cbx_1__1__49_chanx_left_out[1] ,
    \cbx_1__1__49_chanx_left_out[2] ,
    \cbx_1__1__49_chanx_left_out[3] ,
    \cbx_1__1__49_chanx_left_out[4] ,
    \cbx_1__1__49_chanx_left_out[5] ,
    \cbx_1__1__49_chanx_left_out[6] ,
    \cbx_1__1__49_chanx_left_out[7] ,
    \cbx_1__1__49_chanx_left_out[8] ,
    \cbx_1__1__49_chanx_left_out[9] ,
    \cbx_1__1__49_chanx_left_out[10] ,
    \cbx_1__1__49_chanx_left_out[11] ,
    \cbx_1__1__49_chanx_left_out[12] ,
    \cbx_1__1__49_chanx_left_out[13] ,
    \cbx_1__1__49_chanx_left_out[14] ,
    \cbx_1__1__49_chanx_left_out[15] ,
    \cbx_1__1__49_chanx_left_out[16] ,
    \cbx_1__1__49_chanx_left_out[17] ,
    \cbx_1__1__49_chanx_left_out[18] ,
    \cbx_1__1__49_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__1__0_chanx_left_out[0] ,
    \sb_8__1__0_chanx_left_out[1] ,
    \sb_8__1__0_chanx_left_out[2] ,
    \sb_8__1__0_chanx_left_out[3] ,
    \sb_8__1__0_chanx_left_out[4] ,
    \sb_8__1__0_chanx_left_out[5] ,
    \sb_8__1__0_chanx_left_out[6] ,
    \sb_8__1__0_chanx_left_out[7] ,
    \sb_8__1__0_chanx_left_out[8] ,
    \sb_8__1__0_chanx_left_out[9] ,
    \sb_8__1__0_chanx_left_out[10] ,
    \sb_8__1__0_chanx_left_out[11] ,
    \sb_8__1__0_chanx_left_out[12] ,
    \sb_8__1__0_chanx_left_out[13] ,
    \sb_8__1__0_chanx_left_out[14] ,
    \sb_8__1__0_chanx_left_out[15] ,
    \sb_8__1__0_chanx_left_out[16] ,
    \sb_8__1__0_chanx_left_out[17] ,
    \sb_8__1__0_chanx_left_out[18] ,
    \sb_8__1__0_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__49_chanx_right_out[0] ,
    \cbx_1__1__49_chanx_right_out[1] ,
    \cbx_1__1__49_chanx_right_out[2] ,
    \cbx_1__1__49_chanx_right_out[3] ,
    \cbx_1__1__49_chanx_right_out[4] ,
    \cbx_1__1__49_chanx_right_out[5] ,
    \cbx_1__1__49_chanx_right_out[6] ,
    \cbx_1__1__49_chanx_right_out[7] ,
    \cbx_1__1__49_chanx_right_out[8] ,
    \cbx_1__1__49_chanx_right_out[9] ,
    \cbx_1__1__49_chanx_right_out[10] ,
    \cbx_1__1__49_chanx_right_out[11] ,
    \cbx_1__1__49_chanx_right_out[12] ,
    \cbx_1__1__49_chanx_right_out[13] ,
    \cbx_1__1__49_chanx_right_out[14] ,
    \cbx_1__1__49_chanx_right_out[15] ,
    \cbx_1__1__49_chanx_right_out[16] ,
    \cbx_1__1__49_chanx_right_out[17] ,
    \cbx_1__1__49_chanx_right_out[18] ,
    \cbx_1__1__49_chanx_right_out[19] }));
 cbx_1__1_ cbx_8__2_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[50] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[50] ),
    .SC_IN_BOT(\scff_Wires[134] ),
    .SC_OUT_TOP(\scff_Wires[135] ),
    .bottom_grid_pin_0_(cbx_1__1__50_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__50_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__50_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__50_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__50_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__50_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__50_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__50_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__50_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__50_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__50_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__50_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__50_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__50_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__50_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__50_bottom_grid_pin_9_),
    .ccff_head(sb_8__1__1_ccff_tail),
    .ccff_tail(cbx_1__1__50_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[205] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__43_chanx_right_out[0] ,
    \sb_1__1__43_chanx_right_out[1] ,
    \sb_1__1__43_chanx_right_out[2] ,
    \sb_1__1__43_chanx_right_out[3] ,
    \sb_1__1__43_chanx_right_out[4] ,
    \sb_1__1__43_chanx_right_out[5] ,
    \sb_1__1__43_chanx_right_out[6] ,
    \sb_1__1__43_chanx_right_out[7] ,
    \sb_1__1__43_chanx_right_out[8] ,
    \sb_1__1__43_chanx_right_out[9] ,
    \sb_1__1__43_chanx_right_out[10] ,
    \sb_1__1__43_chanx_right_out[11] ,
    \sb_1__1__43_chanx_right_out[12] ,
    \sb_1__1__43_chanx_right_out[13] ,
    \sb_1__1__43_chanx_right_out[14] ,
    \sb_1__1__43_chanx_right_out[15] ,
    \sb_1__1__43_chanx_right_out[16] ,
    \sb_1__1__43_chanx_right_out[17] ,
    \sb_1__1__43_chanx_right_out[18] ,
    \sb_1__1__43_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__50_chanx_left_out[0] ,
    \cbx_1__1__50_chanx_left_out[1] ,
    \cbx_1__1__50_chanx_left_out[2] ,
    \cbx_1__1__50_chanx_left_out[3] ,
    \cbx_1__1__50_chanx_left_out[4] ,
    \cbx_1__1__50_chanx_left_out[5] ,
    \cbx_1__1__50_chanx_left_out[6] ,
    \cbx_1__1__50_chanx_left_out[7] ,
    \cbx_1__1__50_chanx_left_out[8] ,
    \cbx_1__1__50_chanx_left_out[9] ,
    \cbx_1__1__50_chanx_left_out[10] ,
    \cbx_1__1__50_chanx_left_out[11] ,
    \cbx_1__1__50_chanx_left_out[12] ,
    \cbx_1__1__50_chanx_left_out[13] ,
    \cbx_1__1__50_chanx_left_out[14] ,
    \cbx_1__1__50_chanx_left_out[15] ,
    \cbx_1__1__50_chanx_left_out[16] ,
    \cbx_1__1__50_chanx_left_out[17] ,
    \cbx_1__1__50_chanx_left_out[18] ,
    \cbx_1__1__50_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__1__1_chanx_left_out[0] ,
    \sb_8__1__1_chanx_left_out[1] ,
    \sb_8__1__1_chanx_left_out[2] ,
    \sb_8__1__1_chanx_left_out[3] ,
    \sb_8__1__1_chanx_left_out[4] ,
    \sb_8__1__1_chanx_left_out[5] ,
    \sb_8__1__1_chanx_left_out[6] ,
    \sb_8__1__1_chanx_left_out[7] ,
    \sb_8__1__1_chanx_left_out[8] ,
    \sb_8__1__1_chanx_left_out[9] ,
    \sb_8__1__1_chanx_left_out[10] ,
    \sb_8__1__1_chanx_left_out[11] ,
    \sb_8__1__1_chanx_left_out[12] ,
    \sb_8__1__1_chanx_left_out[13] ,
    \sb_8__1__1_chanx_left_out[14] ,
    \sb_8__1__1_chanx_left_out[15] ,
    \sb_8__1__1_chanx_left_out[16] ,
    \sb_8__1__1_chanx_left_out[17] ,
    \sb_8__1__1_chanx_left_out[18] ,
    \sb_8__1__1_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__50_chanx_right_out[0] ,
    \cbx_1__1__50_chanx_right_out[1] ,
    \cbx_1__1__50_chanx_right_out[2] ,
    \cbx_1__1__50_chanx_right_out[3] ,
    \cbx_1__1__50_chanx_right_out[4] ,
    \cbx_1__1__50_chanx_right_out[5] ,
    \cbx_1__1__50_chanx_right_out[6] ,
    \cbx_1__1__50_chanx_right_out[7] ,
    \cbx_1__1__50_chanx_right_out[8] ,
    \cbx_1__1__50_chanx_right_out[9] ,
    \cbx_1__1__50_chanx_right_out[10] ,
    \cbx_1__1__50_chanx_right_out[11] ,
    \cbx_1__1__50_chanx_right_out[12] ,
    \cbx_1__1__50_chanx_right_out[13] ,
    \cbx_1__1__50_chanx_right_out[14] ,
    \cbx_1__1__50_chanx_right_out[15] ,
    \cbx_1__1__50_chanx_right_out[16] ,
    \cbx_1__1__50_chanx_right_out[17] ,
    \cbx_1__1__50_chanx_right_out[18] ,
    \cbx_1__1__50_chanx_right_out[19] }));
 cbx_1__1_ cbx_8__3_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[51] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[51] ),
    .SC_IN_BOT(\scff_Wires[136] ),
    .SC_OUT_TOP(\scff_Wires[137] ),
    .bottom_grid_pin_0_(cbx_1__1__51_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__51_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__51_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__51_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__51_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__51_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__51_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__51_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__51_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__51_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__51_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__51_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__51_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__51_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__51_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__51_bottom_grid_pin_9_),
    .ccff_head(sb_8__1__2_ccff_tail),
    .ccff_tail(cbx_1__1__51_ccff_tail),
    .clk_1_N_out(\clk_1_wires[96] ),
    .clk_1_S_out(\clk_1_wires[97] ),
    .clk_1_W_in(\clk_1_wires[92] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[208] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[96] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[97] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[92] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__44_chanx_right_out[0] ,
    \sb_1__1__44_chanx_right_out[1] ,
    \sb_1__1__44_chanx_right_out[2] ,
    \sb_1__1__44_chanx_right_out[3] ,
    \sb_1__1__44_chanx_right_out[4] ,
    \sb_1__1__44_chanx_right_out[5] ,
    \sb_1__1__44_chanx_right_out[6] ,
    \sb_1__1__44_chanx_right_out[7] ,
    \sb_1__1__44_chanx_right_out[8] ,
    \sb_1__1__44_chanx_right_out[9] ,
    \sb_1__1__44_chanx_right_out[10] ,
    \sb_1__1__44_chanx_right_out[11] ,
    \sb_1__1__44_chanx_right_out[12] ,
    \sb_1__1__44_chanx_right_out[13] ,
    \sb_1__1__44_chanx_right_out[14] ,
    \sb_1__1__44_chanx_right_out[15] ,
    \sb_1__1__44_chanx_right_out[16] ,
    \sb_1__1__44_chanx_right_out[17] ,
    \sb_1__1__44_chanx_right_out[18] ,
    \sb_1__1__44_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__51_chanx_left_out[0] ,
    \cbx_1__1__51_chanx_left_out[1] ,
    \cbx_1__1__51_chanx_left_out[2] ,
    \cbx_1__1__51_chanx_left_out[3] ,
    \cbx_1__1__51_chanx_left_out[4] ,
    \cbx_1__1__51_chanx_left_out[5] ,
    \cbx_1__1__51_chanx_left_out[6] ,
    \cbx_1__1__51_chanx_left_out[7] ,
    \cbx_1__1__51_chanx_left_out[8] ,
    \cbx_1__1__51_chanx_left_out[9] ,
    \cbx_1__1__51_chanx_left_out[10] ,
    \cbx_1__1__51_chanx_left_out[11] ,
    \cbx_1__1__51_chanx_left_out[12] ,
    \cbx_1__1__51_chanx_left_out[13] ,
    \cbx_1__1__51_chanx_left_out[14] ,
    \cbx_1__1__51_chanx_left_out[15] ,
    \cbx_1__1__51_chanx_left_out[16] ,
    \cbx_1__1__51_chanx_left_out[17] ,
    \cbx_1__1__51_chanx_left_out[18] ,
    \cbx_1__1__51_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__1__2_chanx_left_out[0] ,
    \sb_8__1__2_chanx_left_out[1] ,
    \sb_8__1__2_chanx_left_out[2] ,
    \sb_8__1__2_chanx_left_out[3] ,
    \sb_8__1__2_chanx_left_out[4] ,
    \sb_8__1__2_chanx_left_out[5] ,
    \sb_8__1__2_chanx_left_out[6] ,
    \sb_8__1__2_chanx_left_out[7] ,
    \sb_8__1__2_chanx_left_out[8] ,
    \sb_8__1__2_chanx_left_out[9] ,
    \sb_8__1__2_chanx_left_out[10] ,
    \sb_8__1__2_chanx_left_out[11] ,
    \sb_8__1__2_chanx_left_out[12] ,
    \sb_8__1__2_chanx_left_out[13] ,
    \sb_8__1__2_chanx_left_out[14] ,
    \sb_8__1__2_chanx_left_out[15] ,
    \sb_8__1__2_chanx_left_out[16] ,
    \sb_8__1__2_chanx_left_out[17] ,
    \sb_8__1__2_chanx_left_out[18] ,
    \sb_8__1__2_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__51_chanx_right_out[0] ,
    \cbx_1__1__51_chanx_right_out[1] ,
    \cbx_1__1__51_chanx_right_out[2] ,
    \cbx_1__1__51_chanx_right_out[3] ,
    \cbx_1__1__51_chanx_right_out[4] ,
    \cbx_1__1__51_chanx_right_out[5] ,
    \cbx_1__1__51_chanx_right_out[6] ,
    \cbx_1__1__51_chanx_right_out[7] ,
    \cbx_1__1__51_chanx_right_out[8] ,
    \cbx_1__1__51_chanx_right_out[9] ,
    \cbx_1__1__51_chanx_right_out[10] ,
    \cbx_1__1__51_chanx_right_out[11] ,
    \cbx_1__1__51_chanx_right_out[12] ,
    \cbx_1__1__51_chanx_right_out[13] ,
    \cbx_1__1__51_chanx_right_out[14] ,
    \cbx_1__1__51_chanx_right_out[15] ,
    \cbx_1__1__51_chanx_right_out[16] ,
    \cbx_1__1__51_chanx_right_out[17] ,
    \cbx_1__1__51_chanx_right_out[18] ,
    \cbx_1__1__51_chanx_right_out[19] }));
 cbx_1__1_ cbx_8__4_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[52] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[52] ),
    .SC_IN_BOT(\scff_Wires[138] ),
    .SC_OUT_TOP(\scff_Wires[139] ),
    .bottom_grid_pin_0_(cbx_1__1__52_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__52_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__52_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__52_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__52_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__52_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__52_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__52_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__52_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__52_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__52_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__52_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__52_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__52_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__52_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__52_bottom_grid_pin_9_),
    .ccff_head(sb_8__1__3_ccff_tail),
    .ccff_tail(cbx_1__1__52_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[211] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__45_chanx_right_out[0] ,
    \sb_1__1__45_chanx_right_out[1] ,
    \sb_1__1__45_chanx_right_out[2] ,
    \sb_1__1__45_chanx_right_out[3] ,
    \sb_1__1__45_chanx_right_out[4] ,
    \sb_1__1__45_chanx_right_out[5] ,
    \sb_1__1__45_chanx_right_out[6] ,
    \sb_1__1__45_chanx_right_out[7] ,
    \sb_1__1__45_chanx_right_out[8] ,
    \sb_1__1__45_chanx_right_out[9] ,
    \sb_1__1__45_chanx_right_out[10] ,
    \sb_1__1__45_chanx_right_out[11] ,
    \sb_1__1__45_chanx_right_out[12] ,
    \sb_1__1__45_chanx_right_out[13] ,
    \sb_1__1__45_chanx_right_out[14] ,
    \sb_1__1__45_chanx_right_out[15] ,
    \sb_1__1__45_chanx_right_out[16] ,
    \sb_1__1__45_chanx_right_out[17] ,
    \sb_1__1__45_chanx_right_out[18] ,
    \sb_1__1__45_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__52_chanx_left_out[0] ,
    \cbx_1__1__52_chanx_left_out[1] ,
    \cbx_1__1__52_chanx_left_out[2] ,
    \cbx_1__1__52_chanx_left_out[3] ,
    \cbx_1__1__52_chanx_left_out[4] ,
    \cbx_1__1__52_chanx_left_out[5] ,
    \cbx_1__1__52_chanx_left_out[6] ,
    \cbx_1__1__52_chanx_left_out[7] ,
    \cbx_1__1__52_chanx_left_out[8] ,
    \cbx_1__1__52_chanx_left_out[9] ,
    \cbx_1__1__52_chanx_left_out[10] ,
    \cbx_1__1__52_chanx_left_out[11] ,
    \cbx_1__1__52_chanx_left_out[12] ,
    \cbx_1__1__52_chanx_left_out[13] ,
    \cbx_1__1__52_chanx_left_out[14] ,
    \cbx_1__1__52_chanx_left_out[15] ,
    \cbx_1__1__52_chanx_left_out[16] ,
    \cbx_1__1__52_chanx_left_out[17] ,
    \cbx_1__1__52_chanx_left_out[18] ,
    \cbx_1__1__52_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__1__3_chanx_left_out[0] ,
    \sb_8__1__3_chanx_left_out[1] ,
    \sb_8__1__3_chanx_left_out[2] ,
    \sb_8__1__3_chanx_left_out[3] ,
    \sb_8__1__3_chanx_left_out[4] ,
    \sb_8__1__3_chanx_left_out[5] ,
    \sb_8__1__3_chanx_left_out[6] ,
    \sb_8__1__3_chanx_left_out[7] ,
    \sb_8__1__3_chanx_left_out[8] ,
    \sb_8__1__3_chanx_left_out[9] ,
    \sb_8__1__3_chanx_left_out[10] ,
    \sb_8__1__3_chanx_left_out[11] ,
    \sb_8__1__3_chanx_left_out[12] ,
    \sb_8__1__3_chanx_left_out[13] ,
    \sb_8__1__3_chanx_left_out[14] ,
    \sb_8__1__3_chanx_left_out[15] ,
    \sb_8__1__3_chanx_left_out[16] ,
    \sb_8__1__3_chanx_left_out[17] ,
    \sb_8__1__3_chanx_left_out[18] ,
    \sb_8__1__3_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__52_chanx_right_out[0] ,
    \cbx_1__1__52_chanx_right_out[1] ,
    \cbx_1__1__52_chanx_right_out[2] ,
    \cbx_1__1__52_chanx_right_out[3] ,
    \cbx_1__1__52_chanx_right_out[4] ,
    \cbx_1__1__52_chanx_right_out[5] ,
    \cbx_1__1__52_chanx_right_out[6] ,
    \cbx_1__1__52_chanx_right_out[7] ,
    \cbx_1__1__52_chanx_right_out[8] ,
    \cbx_1__1__52_chanx_right_out[9] ,
    \cbx_1__1__52_chanx_right_out[10] ,
    \cbx_1__1__52_chanx_right_out[11] ,
    \cbx_1__1__52_chanx_right_out[12] ,
    \cbx_1__1__52_chanx_right_out[13] ,
    \cbx_1__1__52_chanx_right_out[14] ,
    \cbx_1__1__52_chanx_right_out[15] ,
    \cbx_1__1__52_chanx_right_out[16] ,
    \cbx_1__1__52_chanx_right_out[17] ,
    \cbx_1__1__52_chanx_right_out[18] ,
    \cbx_1__1__52_chanx_right_out[19] }));
 cbx_1__1_ cbx_8__5_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[53] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[53] ),
    .SC_IN_BOT(\scff_Wires[140] ),
    .SC_OUT_TOP(\scff_Wires[141] ),
    .bottom_grid_pin_0_(cbx_1__1__53_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__53_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__53_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__53_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__53_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__53_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__53_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__53_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__53_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__53_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__53_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__53_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__53_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__53_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__53_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__53_bottom_grid_pin_9_),
    .ccff_head(sb_8__1__4_ccff_tail),
    .ccff_tail(cbx_1__1__53_ccff_tail),
    .clk_1_N_out(\clk_1_wires[103] ),
    .clk_1_S_out(\clk_1_wires[104] ),
    .clk_1_W_in(\clk_1_wires[99] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[214] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[103] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[104] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[99] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__46_chanx_right_out[0] ,
    \sb_1__1__46_chanx_right_out[1] ,
    \sb_1__1__46_chanx_right_out[2] ,
    \sb_1__1__46_chanx_right_out[3] ,
    \sb_1__1__46_chanx_right_out[4] ,
    \sb_1__1__46_chanx_right_out[5] ,
    \sb_1__1__46_chanx_right_out[6] ,
    \sb_1__1__46_chanx_right_out[7] ,
    \sb_1__1__46_chanx_right_out[8] ,
    \sb_1__1__46_chanx_right_out[9] ,
    \sb_1__1__46_chanx_right_out[10] ,
    \sb_1__1__46_chanx_right_out[11] ,
    \sb_1__1__46_chanx_right_out[12] ,
    \sb_1__1__46_chanx_right_out[13] ,
    \sb_1__1__46_chanx_right_out[14] ,
    \sb_1__1__46_chanx_right_out[15] ,
    \sb_1__1__46_chanx_right_out[16] ,
    \sb_1__1__46_chanx_right_out[17] ,
    \sb_1__1__46_chanx_right_out[18] ,
    \sb_1__1__46_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__53_chanx_left_out[0] ,
    \cbx_1__1__53_chanx_left_out[1] ,
    \cbx_1__1__53_chanx_left_out[2] ,
    \cbx_1__1__53_chanx_left_out[3] ,
    \cbx_1__1__53_chanx_left_out[4] ,
    \cbx_1__1__53_chanx_left_out[5] ,
    \cbx_1__1__53_chanx_left_out[6] ,
    \cbx_1__1__53_chanx_left_out[7] ,
    \cbx_1__1__53_chanx_left_out[8] ,
    \cbx_1__1__53_chanx_left_out[9] ,
    \cbx_1__1__53_chanx_left_out[10] ,
    \cbx_1__1__53_chanx_left_out[11] ,
    \cbx_1__1__53_chanx_left_out[12] ,
    \cbx_1__1__53_chanx_left_out[13] ,
    \cbx_1__1__53_chanx_left_out[14] ,
    \cbx_1__1__53_chanx_left_out[15] ,
    \cbx_1__1__53_chanx_left_out[16] ,
    \cbx_1__1__53_chanx_left_out[17] ,
    \cbx_1__1__53_chanx_left_out[18] ,
    \cbx_1__1__53_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__1__4_chanx_left_out[0] ,
    \sb_8__1__4_chanx_left_out[1] ,
    \sb_8__1__4_chanx_left_out[2] ,
    \sb_8__1__4_chanx_left_out[3] ,
    \sb_8__1__4_chanx_left_out[4] ,
    \sb_8__1__4_chanx_left_out[5] ,
    \sb_8__1__4_chanx_left_out[6] ,
    \sb_8__1__4_chanx_left_out[7] ,
    \sb_8__1__4_chanx_left_out[8] ,
    \sb_8__1__4_chanx_left_out[9] ,
    \sb_8__1__4_chanx_left_out[10] ,
    \sb_8__1__4_chanx_left_out[11] ,
    \sb_8__1__4_chanx_left_out[12] ,
    \sb_8__1__4_chanx_left_out[13] ,
    \sb_8__1__4_chanx_left_out[14] ,
    \sb_8__1__4_chanx_left_out[15] ,
    \sb_8__1__4_chanx_left_out[16] ,
    \sb_8__1__4_chanx_left_out[17] ,
    \sb_8__1__4_chanx_left_out[18] ,
    \sb_8__1__4_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__53_chanx_right_out[0] ,
    \cbx_1__1__53_chanx_right_out[1] ,
    \cbx_1__1__53_chanx_right_out[2] ,
    \cbx_1__1__53_chanx_right_out[3] ,
    \cbx_1__1__53_chanx_right_out[4] ,
    \cbx_1__1__53_chanx_right_out[5] ,
    \cbx_1__1__53_chanx_right_out[6] ,
    \cbx_1__1__53_chanx_right_out[7] ,
    \cbx_1__1__53_chanx_right_out[8] ,
    \cbx_1__1__53_chanx_right_out[9] ,
    \cbx_1__1__53_chanx_right_out[10] ,
    \cbx_1__1__53_chanx_right_out[11] ,
    \cbx_1__1__53_chanx_right_out[12] ,
    \cbx_1__1__53_chanx_right_out[13] ,
    \cbx_1__1__53_chanx_right_out[14] ,
    \cbx_1__1__53_chanx_right_out[15] ,
    \cbx_1__1__53_chanx_right_out[16] ,
    \cbx_1__1__53_chanx_right_out[17] ,
    \cbx_1__1__53_chanx_right_out[18] ,
    \cbx_1__1__53_chanx_right_out[19] }));
 cbx_1__1_ cbx_8__6_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[54] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[54] ),
    .SC_IN_BOT(\scff_Wires[142] ),
    .SC_OUT_TOP(\scff_Wires[143] ),
    .bottom_grid_pin_0_(cbx_1__1__54_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__54_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__54_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__54_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__54_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__54_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__54_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__54_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__54_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__54_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__54_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__54_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__54_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__54_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__54_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__54_bottom_grid_pin_9_),
    .ccff_head(sb_8__1__5_ccff_tail),
    .ccff_tail(cbx_1__1__54_ccff_tail),
    .prog_clk_0_N_in(\prog_clk_0_wires[217] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__47_chanx_right_out[0] ,
    \sb_1__1__47_chanx_right_out[1] ,
    \sb_1__1__47_chanx_right_out[2] ,
    \sb_1__1__47_chanx_right_out[3] ,
    \sb_1__1__47_chanx_right_out[4] ,
    \sb_1__1__47_chanx_right_out[5] ,
    \sb_1__1__47_chanx_right_out[6] ,
    \sb_1__1__47_chanx_right_out[7] ,
    \sb_1__1__47_chanx_right_out[8] ,
    \sb_1__1__47_chanx_right_out[9] ,
    \sb_1__1__47_chanx_right_out[10] ,
    \sb_1__1__47_chanx_right_out[11] ,
    \sb_1__1__47_chanx_right_out[12] ,
    \sb_1__1__47_chanx_right_out[13] ,
    \sb_1__1__47_chanx_right_out[14] ,
    \sb_1__1__47_chanx_right_out[15] ,
    \sb_1__1__47_chanx_right_out[16] ,
    \sb_1__1__47_chanx_right_out[17] ,
    \sb_1__1__47_chanx_right_out[18] ,
    \sb_1__1__47_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__54_chanx_left_out[0] ,
    \cbx_1__1__54_chanx_left_out[1] ,
    \cbx_1__1__54_chanx_left_out[2] ,
    \cbx_1__1__54_chanx_left_out[3] ,
    \cbx_1__1__54_chanx_left_out[4] ,
    \cbx_1__1__54_chanx_left_out[5] ,
    \cbx_1__1__54_chanx_left_out[6] ,
    \cbx_1__1__54_chanx_left_out[7] ,
    \cbx_1__1__54_chanx_left_out[8] ,
    \cbx_1__1__54_chanx_left_out[9] ,
    \cbx_1__1__54_chanx_left_out[10] ,
    \cbx_1__1__54_chanx_left_out[11] ,
    \cbx_1__1__54_chanx_left_out[12] ,
    \cbx_1__1__54_chanx_left_out[13] ,
    \cbx_1__1__54_chanx_left_out[14] ,
    \cbx_1__1__54_chanx_left_out[15] ,
    \cbx_1__1__54_chanx_left_out[16] ,
    \cbx_1__1__54_chanx_left_out[17] ,
    \cbx_1__1__54_chanx_left_out[18] ,
    \cbx_1__1__54_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__1__5_chanx_left_out[0] ,
    \sb_8__1__5_chanx_left_out[1] ,
    \sb_8__1__5_chanx_left_out[2] ,
    \sb_8__1__5_chanx_left_out[3] ,
    \sb_8__1__5_chanx_left_out[4] ,
    \sb_8__1__5_chanx_left_out[5] ,
    \sb_8__1__5_chanx_left_out[6] ,
    \sb_8__1__5_chanx_left_out[7] ,
    \sb_8__1__5_chanx_left_out[8] ,
    \sb_8__1__5_chanx_left_out[9] ,
    \sb_8__1__5_chanx_left_out[10] ,
    \sb_8__1__5_chanx_left_out[11] ,
    \sb_8__1__5_chanx_left_out[12] ,
    \sb_8__1__5_chanx_left_out[13] ,
    \sb_8__1__5_chanx_left_out[14] ,
    \sb_8__1__5_chanx_left_out[15] ,
    \sb_8__1__5_chanx_left_out[16] ,
    \sb_8__1__5_chanx_left_out[17] ,
    \sb_8__1__5_chanx_left_out[18] ,
    \sb_8__1__5_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__54_chanx_right_out[0] ,
    \cbx_1__1__54_chanx_right_out[1] ,
    \cbx_1__1__54_chanx_right_out[2] ,
    \cbx_1__1__54_chanx_right_out[3] ,
    \cbx_1__1__54_chanx_right_out[4] ,
    \cbx_1__1__54_chanx_right_out[5] ,
    \cbx_1__1__54_chanx_right_out[6] ,
    \cbx_1__1__54_chanx_right_out[7] ,
    \cbx_1__1__54_chanx_right_out[8] ,
    \cbx_1__1__54_chanx_right_out[9] ,
    \cbx_1__1__54_chanx_right_out[10] ,
    \cbx_1__1__54_chanx_right_out[11] ,
    \cbx_1__1__54_chanx_right_out[12] ,
    \cbx_1__1__54_chanx_right_out[13] ,
    \cbx_1__1__54_chanx_right_out[14] ,
    \cbx_1__1__54_chanx_right_out[15] ,
    \cbx_1__1__54_chanx_right_out[16] ,
    \cbx_1__1__54_chanx_right_out[17] ,
    \cbx_1__1__54_chanx_right_out[18] ,
    \cbx_1__1__54_chanx_right_out[19] }));
 cbx_1__1_ cbx_8__7_ (.REGIN_FEEDTHROUGH(\regin_feedthrough_wires[55] ),
    .REGOUT_FEEDTHROUGH(\regout_feedthrough_wires[55] ),
    .SC_IN_BOT(\scff_Wires[144] ),
    .SC_OUT_TOP(\scff_Wires[145] ),
    .bottom_grid_pin_0_(cbx_1__1__55_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__1__55_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__1__55_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__1__55_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__1__55_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__1__55_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__1__55_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__1__55_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__1__55_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__1__55_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__1__55_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__1__55_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__1__55_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__1__55_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__1__55_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__1__55_bottom_grid_pin_9_),
    .ccff_head(sb_8__1__6_ccff_tail),
    .ccff_tail(cbx_1__1__55_ccff_tail),
    .clk_1_N_out(\clk_1_wires[110] ),
    .clk_1_S_out(\clk_1_wires[111] ),
    .clk_1_W_in(\clk_1_wires[106] ),
    .prog_clk_0_N_in(\prog_clk_0_wires[220] ),
    .prog_clk_1_N_out(\prog_clk_1_wires[110] ),
    .prog_clk_1_S_out(\prog_clk_1_wires[111] ),
    .prog_clk_1_W_in(\prog_clk_1_wires[106] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__1__48_chanx_right_out[0] ,
    \sb_1__1__48_chanx_right_out[1] ,
    \sb_1__1__48_chanx_right_out[2] ,
    \sb_1__1__48_chanx_right_out[3] ,
    \sb_1__1__48_chanx_right_out[4] ,
    \sb_1__1__48_chanx_right_out[5] ,
    \sb_1__1__48_chanx_right_out[6] ,
    \sb_1__1__48_chanx_right_out[7] ,
    \sb_1__1__48_chanx_right_out[8] ,
    \sb_1__1__48_chanx_right_out[9] ,
    \sb_1__1__48_chanx_right_out[10] ,
    \sb_1__1__48_chanx_right_out[11] ,
    \sb_1__1__48_chanx_right_out[12] ,
    \sb_1__1__48_chanx_right_out[13] ,
    \sb_1__1__48_chanx_right_out[14] ,
    \sb_1__1__48_chanx_right_out[15] ,
    \sb_1__1__48_chanx_right_out[16] ,
    \sb_1__1__48_chanx_right_out[17] ,
    \sb_1__1__48_chanx_right_out[18] ,
    \sb_1__1__48_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__1__55_chanx_left_out[0] ,
    \cbx_1__1__55_chanx_left_out[1] ,
    \cbx_1__1__55_chanx_left_out[2] ,
    \cbx_1__1__55_chanx_left_out[3] ,
    \cbx_1__1__55_chanx_left_out[4] ,
    \cbx_1__1__55_chanx_left_out[5] ,
    \cbx_1__1__55_chanx_left_out[6] ,
    \cbx_1__1__55_chanx_left_out[7] ,
    \cbx_1__1__55_chanx_left_out[8] ,
    \cbx_1__1__55_chanx_left_out[9] ,
    \cbx_1__1__55_chanx_left_out[10] ,
    \cbx_1__1__55_chanx_left_out[11] ,
    \cbx_1__1__55_chanx_left_out[12] ,
    \cbx_1__1__55_chanx_left_out[13] ,
    \cbx_1__1__55_chanx_left_out[14] ,
    \cbx_1__1__55_chanx_left_out[15] ,
    \cbx_1__1__55_chanx_left_out[16] ,
    \cbx_1__1__55_chanx_left_out[17] ,
    \cbx_1__1__55_chanx_left_out[18] ,
    \cbx_1__1__55_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__1__6_chanx_left_out[0] ,
    \sb_8__1__6_chanx_left_out[1] ,
    \sb_8__1__6_chanx_left_out[2] ,
    \sb_8__1__6_chanx_left_out[3] ,
    \sb_8__1__6_chanx_left_out[4] ,
    \sb_8__1__6_chanx_left_out[5] ,
    \sb_8__1__6_chanx_left_out[6] ,
    \sb_8__1__6_chanx_left_out[7] ,
    \sb_8__1__6_chanx_left_out[8] ,
    \sb_8__1__6_chanx_left_out[9] ,
    \sb_8__1__6_chanx_left_out[10] ,
    \sb_8__1__6_chanx_left_out[11] ,
    \sb_8__1__6_chanx_left_out[12] ,
    \sb_8__1__6_chanx_left_out[13] ,
    \sb_8__1__6_chanx_left_out[14] ,
    \sb_8__1__6_chanx_left_out[15] ,
    \sb_8__1__6_chanx_left_out[16] ,
    \sb_8__1__6_chanx_left_out[17] ,
    \sb_8__1__6_chanx_left_out[18] ,
    \sb_8__1__6_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__1__55_chanx_right_out[0] ,
    \cbx_1__1__55_chanx_right_out[1] ,
    \cbx_1__1__55_chanx_right_out[2] ,
    \cbx_1__1__55_chanx_right_out[3] ,
    \cbx_1__1__55_chanx_right_out[4] ,
    \cbx_1__1__55_chanx_right_out[5] ,
    \cbx_1__1__55_chanx_right_out[6] ,
    \cbx_1__1__55_chanx_right_out[7] ,
    \cbx_1__1__55_chanx_right_out[8] ,
    \cbx_1__1__55_chanx_right_out[9] ,
    \cbx_1__1__55_chanx_right_out[10] ,
    \cbx_1__1__55_chanx_right_out[11] ,
    \cbx_1__1__55_chanx_right_out[12] ,
    \cbx_1__1__55_chanx_right_out[13] ,
    \cbx_1__1__55_chanx_right_out[14] ,
    \cbx_1__1__55_chanx_right_out[15] ,
    \cbx_1__1__55_chanx_right_out[16] ,
    \cbx_1__1__55_chanx_right_out[17] ,
    \cbx_1__1__55_chanx_right_out[18] ,
    \cbx_1__1__55_chanx_right_out[19] }));
 cbx_1__2_ cbx_8__8_ (.IO_ISOL_N(IO_ISOL_N),
    .SC_IN_BOT(\scff_Wires[146] ),
    .SC_OUT_TOP(\scff_Wires[147] ),
    .bottom_grid_pin_0_(cbx_1__8__7_bottom_grid_pin_0_),
    .bottom_grid_pin_10_(cbx_1__8__7_bottom_grid_pin_10_),
    .bottom_grid_pin_11_(cbx_1__8__7_bottom_grid_pin_11_),
    .bottom_grid_pin_12_(cbx_1__8__7_bottom_grid_pin_12_),
    .bottom_grid_pin_13_(cbx_1__8__7_bottom_grid_pin_13_),
    .bottom_grid_pin_14_(cbx_1__8__7_bottom_grid_pin_14_),
    .bottom_grid_pin_15_(cbx_1__8__7_bottom_grid_pin_15_),
    .bottom_grid_pin_1_(cbx_1__8__7_bottom_grid_pin_1_),
    .bottom_grid_pin_2_(cbx_1__8__7_bottom_grid_pin_2_),
    .bottom_grid_pin_3_(cbx_1__8__7_bottom_grid_pin_3_),
    .bottom_grid_pin_4_(cbx_1__8__7_bottom_grid_pin_4_),
    .bottom_grid_pin_5_(cbx_1__8__7_bottom_grid_pin_5_),
    .bottom_grid_pin_6_(cbx_1__8__7_bottom_grid_pin_6_),
    .bottom_grid_pin_7_(cbx_1__8__7_bottom_grid_pin_7_),
    .bottom_grid_pin_8_(cbx_1__8__7_bottom_grid_pin_8_),
    .bottom_grid_pin_9_(cbx_1__8__7_bottom_grid_pin_9_),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__7_top_grid_pin_0_),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_7_bottom_width_0_height_0__pin_1_lower),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_7_bottom_width_0_height_0__pin_1_upper),
    .ccff_head(sb_8__8__0_ccff_tail),
    .ccff_tail(grid_io_top_7_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]),
    .prog_clk_0_S_in(\prog_clk_0_wires[223] ),
    .top_grid_pin_0_(cbx_1__8__7_top_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\sb_1__8__6_chanx_right_out[0] ,
    \sb_1__8__6_chanx_right_out[1] ,
    \sb_1__8__6_chanx_right_out[2] ,
    \sb_1__8__6_chanx_right_out[3] ,
    \sb_1__8__6_chanx_right_out[4] ,
    \sb_1__8__6_chanx_right_out[5] ,
    \sb_1__8__6_chanx_right_out[6] ,
    \sb_1__8__6_chanx_right_out[7] ,
    \sb_1__8__6_chanx_right_out[8] ,
    \sb_1__8__6_chanx_right_out[9] ,
    \sb_1__8__6_chanx_right_out[10] ,
    \sb_1__8__6_chanx_right_out[11] ,
    \sb_1__8__6_chanx_right_out[12] ,
    \sb_1__8__6_chanx_right_out[13] ,
    \sb_1__8__6_chanx_right_out[14] ,
    \sb_1__8__6_chanx_right_out[15] ,
    \sb_1__8__6_chanx_right_out[16] ,
    \sb_1__8__6_chanx_right_out[17] ,
    \sb_1__8__6_chanx_right_out[18] ,
    \sb_1__8__6_chanx_right_out[19] }),
    .chanx_left_out({\cbx_1__8__7_chanx_left_out[0] ,
    \cbx_1__8__7_chanx_left_out[1] ,
    \cbx_1__8__7_chanx_left_out[2] ,
    \cbx_1__8__7_chanx_left_out[3] ,
    \cbx_1__8__7_chanx_left_out[4] ,
    \cbx_1__8__7_chanx_left_out[5] ,
    \cbx_1__8__7_chanx_left_out[6] ,
    \cbx_1__8__7_chanx_left_out[7] ,
    \cbx_1__8__7_chanx_left_out[8] ,
    \cbx_1__8__7_chanx_left_out[9] ,
    \cbx_1__8__7_chanx_left_out[10] ,
    \cbx_1__8__7_chanx_left_out[11] ,
    \cbx_1__8__7_chanx_left_out[12] ,
    \cbx_1__8__7_chanx_left_out[13] ,
    \cbx_1__8__7_chanx_left_out[14] ,
    \cbx_1__8__7_chanx_left_out[15] ,
    \cbx_1__8__7_chanx_left_out[16] ,
    \cbx_1__8__7_chanx_left_out[17] ,
    \cbx_1__8__7_chanx_left_out[18] ,
    \cbx_1__8__7_chanx_left_out[19] }),
    .chanx_right_in({\sb_8__8__0_chanx_left_out[0] ,
    \sb_8__8__0_chanx_left_out[1] ,
    \sb_8__8__0_chanx_left_out[2] ,
    \sb_8__8__0_chanx_left_out[3] ,
    \sb_8__8__0_chanx_left_out[4] ,
    \sb_8__8__0_chanx_left_out[5] ,
    \sb_8__8__0_chanx_left_out[6] ,
    \sb_8__8__0_chanx_left_out[7] ,
    \sb_8__8__0_chanx_left_out[8] ,
    \sb_8__8__0_chanx_left_out[9] ,
    \sb_8__8__0_chanx_left_out[10] ,
    \sb_8__8__0_chanx_left_out[11] ,
    \sb_8__8__0_chanx_left_out[12] ,
    \sb_8__8__0_chanx_left_out[13] ,
    \sb_8__8__0_chanx_left_out[14] ,
    \sb_8__8__0_chanx_left_out[15] ,
    \sb_8__8__0_chanx_left_out[16] ,
    \sb_8__8__0_chanx_left_out[17] ,
    \sb_8__8__0_chanx_left_out[18] ,
    \sb_8__8__0_chanx_left_out[19] }),
    .chanx_right_out({\cbx_1__8__7_chanx_right_out[0] ,
    \cbx_1__8__7_chanx_right_out[1] ,
    \cbx_1__8__7_chanx_right_out[2] ,
    \cbx_1__8__7_chanx_right_out[3] ,
    \cbx_1__8__7_chanx_right_out[4] ,
    \cbx_1__8__7_chanx_right_out[5] ,
    \cbx_1__8__7_chanx_right_out[6] ,
    \cbx_1__8__7_chanx_right_out[7] ,
    \cbx_1__8__7_chanx_right_out[8] ,
    \cbx_1__8__7_chanx_right_out[9] ,
    \cbx_1__8__7_chanx_right_out[10] ,
    \cbx_1__8__7_chanx_right_out[11] ,
    \cbx_1__8__7_chanx_right_out[12] ,
    \cbx_1__8__7_chanx_right_out[13] ,
    \cbx_1__8__7_chanx_right_out[14] ,
    \cbx_1__8__7_chanx_right_out[15] ,
    \cbx_1__8__7_chanx_right_out[16] ,
    \cbx_1__8__7_chanx_right_out[17] ,
    \cbx_1__8__7_chanx_right_out[18] ,
    \cbx_1__8__7_chanx_right_out[19] }));
 cby_0__1_ cby_0__1_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__1__0_ccff_tail),
    .ccff_tail(grid_io_left_0_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]),
    .left_grid_pin_0_(cby_0__1__0_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[3] ),
    .right_width_0_height_0__pin_0_(cby_0__1__0_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_0_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_0_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__0__0_chany_top_out[0] ,
    \sb_0__0__0_chany_top_out[1] ,
    \sb_0__0__0_chany_top_out[2] ,
    \sb_0__0__0_chany_top_out[3] ,
    \sb_0__0__0_chany_top_out[4] ,
    \sb_0__0__0_chany_top_out[5] ,
    \sb_0__0__0_chany_top_out[6] ,
    \sb_0__0__0_chany_top_out[7] ,
    \sb_0__0__0_chany_top_out[8] ,
    \sb_0__0__0_chany_top_out[9] ,
    \sb_0__0__0_chany_top_out[10] ,
    \sb_0__0__0_chany_top_out[11] ,
    \sb_0__0__0_chany_top_out[12] ,
    \sb_0__0__0_chany_top_out[13] ,
    \sb_0__0__0_chany_top_out[14] ,
    \sb_0__0__0_chany_top_out[15] ,
    \sb_0__0__0_chany_top_out[16] ,
    \sb_0__0__0_chany_top_out[17] ,
    \sb_0__0__0_chany_top_out[18] ,
    \sb_0__0__0_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__0_chany_bottom_out[0] ,
    \cby_0__1__0_chany_bottom_out[1] ,
    \cby_0__1__0_chany_bottom_out[2] ,
    \cby_0__1__0_chany_bottom_out[3] ,
    \cby_0__1__0_chany_bottom_out[4] ,
    \cby_0__1__0_chany_bottom_out[5] ,
    \cby_0__1__0_chany_bottom_out[6] ,
    \cby_0__1__0_chany_bottom_out[7] ,
    \cby_0__1__0_chany_bottom_out[8] ,
    \cby_0__1__0_chany_bottom_out[9] ,
    \cby_0__1__0_chany_bottom_out[10] ,
    \cby_0__1__0_chany_bottom_out[11] ,
    \cby_0__1__0_chany_bottom_out[12] ,
    \cby_0__1__0_chany_bottom_out[13] ,
    \cby_0__1__0_chany_bottom_out[14] ,
    \cby_0__1__0_chany_bottom_out[15] ,
    \cby_0__1__0_chany_bottom_out[16] ,
    \cby_0__1__0_chany_bottom_out[17] ,
    \cby_0__1__0_chany_bottom_out[18] ,
    \cby_0__1__0_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__1__0_chany_bottom_out[0] ,
    \sb_0__1__0_chany_bottom_out[1] ,
    \sb_0__1__0_chany_bottom_out[2] ,
    \sb_0__1__0_chany_bottom_out[3] ,
    \sb_0__1__0_chany_bottom_out[4] ,
    \sb_0__1__0_chany_bottom_out[5] ,
    \sb_0__1__0_chany_bottom_out[6] ,
    \sb_0__1__0_chany_bottom_out[7] ,
    \sb_0__1__0_chany_bottom_out[8] ,
    \sb_0__1__0_chany_bottom_out[9] ,
    \sb_0__1__0_chany_bottom_out[10] ,
    \sb_0__1__0_chany_bottom_out[11] ,
    \sb_0__1__0_chany_bottom_out[12] ,
    \sb_0__1__0_chany_bottom_out[13] ,
    \sb_0__1__0_chany_bottom_out[14] ,
    \sb_0__1__0_chany_bottom_out[15] ,
    \sb_0__1__0_chany_bottom_out[16] ,
    \sb_0__1__0_chany_bottom_out[17] ,
    \sb_0__1__0_chany_bottom_out[18] ,
    \sb_0__1__0_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__0_chany_top_out[0] ,
    \cby_0__1__0_chany_top_out[1] ,
    \cby_0__1__0_chany_top_out[2] ,
    \cby_0__1__0_chany_top_out[3] ,
    \cby_0__1__0_chany_top_out[4] ,
    \cby_0__1__0_chany_top_out[5] ,
    \cby_0__1__0_chany_top_out[6] ,
    \cby_0__1__0_chany_top_out[7] ,
    \cby_0__1__0_chany_top_out[8] ,
    \cby_0__1__0_chany_top_out[9] ,
    \cby_0__1__0_chany_top_out[10] ,
    \cby_0__1__0_chany_top_out[11] ,
    \cby_0__1__0_chany_top_out[12] ,
    \cby_0__1__0_chany_top_out[13] ,
    \cby_0__1__0_chany_top_out[14] ,
    \cby_0__1__0_chany_top_out[15] ,
    \cby_0__1__0_chany_top_out[16] ,
    \cby_0__1__0_chany_top_out[17] ,
    \cby_0__1__0_chany_top_out[18] ,
    \cby_0__1__0_chany_top_out[19] }));
 cby_0__1_ cby_0__2_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__1__1_ccff_tail),
    .ccff_tail(grid_io_left_1_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]),
    .left_grid_pin_0_(cby_0__1__1_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[9] ),
    .right_width_0_height_0__pin_0_(cby_0__1__1_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_1_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_1_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__1__0_chany_top_out[0] ,
    \sb_0__1__0_chany_top_out[1] ,
    \sb_0__1__0_chany_top_out[2] ,
    \sb_0__1__0_chany_top_out[3] ,
    \sb_0__1__0_chany_top_out[4] ,
    \sb_0__1__0_chany_top_out[5] ,
    \sb_0__1__0_chany_top_out[6] ,
    \sb_0__1__0_chany_top_out[7] ,
    \sb_0__1__0_chany_top_out[8] ,
    \sb_0__1__0_chany_top_out[9] ,
    \sb_0__1__0_chany_top_out[10] ,
    \sb_0__1__0_chany_top_out[11] ,
    \sb_0__1__0_chany_top_out[12] ,
    \sb_0__1__0_chany_top_out[13] ,
    \sb_0__1__0_chany_top_out[14] ,
    \sb_0__1__0_chany_top_out[15] ,
    \sb_0__1__0_chany_top_out[16] ,
    \sb_0__1__0_chany_top_out[17] ,
    \sb_0__1__0_chany_top_out[18] ,
    \sb_0__1__0_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__1_chany_bottom_out[0] ,
    \cby_0__1__1_chany_bottom_out[1] ,
    \cby_0__1__1_chany_bottom_out[2] ,
    \cby_0__1__1_chany_bottom_out[3] ,
    \cby_0__1__1_chany_bottom_out[4] ,
    \cby_0__1__1_chany_bottom_out[5] ,
    \cby_0__1__1_chany_bottom_out[6] ,
    \cby_0__1__1_chany_bottom_out[7] ,
    \cby_0__1__1_chany_bottom_out[8] ,
    \cby_0__1__1_chany_bottom_out[9] ,
    \cby_0__1__1_chany_bottom_out[10] ,
    \cby_0__1__1_chany_bottom_out[11] ,
    \cby_0__1__1_chany_bottom_out[12] ,
    \cby_0__1__1_chany_bottom_out[13] ,
    \cby_0__1__1_chany_bottom_out[14] ,
    \cby_0__1__1_chany_bottom_out[15] ,
    \cby_0__1__1_chany_bottom_out[16] ,
    \cby_0__1__1_chany_bottom_out[17] ,
    \cby_0__1__1_chany_bottom_out[18] ,
    \cby_0__1__1_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__1__1_chany_bottom_out[0] ,
    \sb_0__1__1_chany_bottom_out[1] ,
    \sb_0__1__1_chany_bottom_out[2] ,
    \sb_0__1__1_chany_bottom_out[3] ,
    \sb_0__1__1_chany_bottom_out[4] ,
    \sb_0__1__1_chany_bottom_out[5] ,
    \sb_0__1__1_chany_bottom_out[6] ,
    \sb_0__1__1_chany_bottom_out[7] ,
    \sb_0__1__1_chany_bottom_out[8] ,
    \sb_0__1__1_chany_bottom_out[9] ,
    \sb_0__1__1_chany_bottom_out[10] ,
    \sb_0__1__1_chany_bottom_out[11] ,
    \sb_0__1__1_chany_bottom_out[12] ,
    \sb_0__1__1_chany_bottom_out[13] ,
    \sb_0__1__1_chany_bottom_out[14] ,
    \sb_0__1__1_chany_bottom_out[15] ,
    \sb_0__1__1_chany_bottom_out[16] ,
    \sb_0__1__1_chany_bottom_out[17] ,
    \sb_0__1__1_chany_bottom_out[18] ,
    \sb_0__1__1_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__1_chany_top_out[0] ,
    \cby_0__1__1_chany_top_out[1] ,
    \cby_0__1__1_chany_top_out[2] ,
    \cby_0__1__1_chany_top_out[3] ,
    \cby_0__1__1_chany_top_out[4] ,
    \cby_0__1__1_chany_top_out[5] ,
    \cby_0__1__1_chany_top_out[6] ,
    \cby_0__1__1_chany_top_out[7] ,
    \cby_0__1__1_chany_top_out[8] ,
    \cby_0__1__1_chany_top_out[9] ,
    \cby_0__1__1_chany_top_out[10] ,
    \cby_0__1__1_chany_top_out[11] ,
    \cby_0__1__1_chany_top_out[12] ,
    \cby_0__1__1_chany_top_out[13] ,
    \cby_0__1__1_chany_top_out[14] ,
    \cby_0__1__1_chany_top_out[15] ,
    \cby_0__1__1_chany_top_out[16] ,
    \cby_0__1__1_chany_top_out[17] ,
    \cby_0__1__1_chany_top_out[18] ,
    \cby_0__1__1_chany_top_out[19] }));
 cby_0__1_ cby_0__3_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__1__2_ccff_tail),
    .ccff_tail(grid_io_left_2_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]),
    .left_grid_pin_0_(cby_0__1__2_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[14] ),
    .right_width_0_height_0__pin_0_(cby_0__1__2_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_2_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_2_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__1__1_chany_top_out[0] ,
    \sb_0__1__1_chany_top_out[1] ,
    \sb_0__1__1_chany_top_out[2] ,
    \sb_0__1__1_chany_top_out[3] ,
    \sb_0__1__1_chany_top_out[4] ,
    \sb_0__1__1_chany_top_out[5] ,
    \sb_0__1__1_chany_top_out[6] ,
    \sb_0__1__1_chany_top_out[7] ,
    \sb_0__1__1_chany_top_out[8] ,
    \sb_0__1__1_chany_top_out[9] ,
    \sb_0__1__1_chany_top_out[10] ,
    \sb_0__1__1_chany_top_out[11] ,
    \sb_0__1__1_chany_top_out[12] ,
    \sb_0__1__1_chany_top_out[13] ,
    \sb_0__1__1_chany_top_out[14] ,
    \sb_0__1__1_chany_top_out[15] ,
    \sb_0__1__1_chany_top_out[16] ,
    \sb_0__1__1_chany_top_out[17] ,
    \sb_0__1__1_chany_top_out[18] ,
    \sb_0__1__1_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__2_chany_bottom_out[0] ,
    \cby_0__1__2_chany_bottom_out[1] ,
    \cby_0__1__2_chany_bottom_out[2] ,
    \cby_0__1__2_chany_bottom_out[3] ,
    \cby_0__1__2_chany_bottom_out[4] ,
    \cby_0__1__2_chany_bottom_out[5] ,
    \cby_0__1__2_chany_bottom_out[6] ,
    \cby_0__1__2_chany_bottom_out[7] ,
    \cby_0__1__2_chany_bottom_out[8] ,
    \cby_0__1__2_chany_bottom_out[9] ,
    \cby_0__1__2_chany_bottom_out[10] ,
    \cby_0__1__2_chany_bottom_out[11] ,
    \cby_0__1__2_chany_bottom_out[12] ,
    \cby_0__1__2_chany_bottom_out[13] ,
    \cby_0__1__2_chany_bottom_out[14] ,
    \cby_0__1__2_chany_bottom_out[15] ,
    \cby_0__1__2_chany_bottom_out[16] ,
    \cby_0__1__2_chany_bottom_out[17] ,
    \cby_0__1__2_chany_bottom_out[18] ,
    \cby_0__1__2_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__1__2_chany_bottom_out[0] ,
    \sb_0__1__2_chany_bottom_out[1] ,
    \sb_0__1__2_chany_bottom_out[2] ,
    \sb_0__1__2_chany_bottom_out[3] ,
    \sb_0__1__2_chany_bottom_out[4] ,
    \sb_0__1__2_chany_bottom_out[5] ,
    \sb_0__1__2_chany_bottom_out[6] ,
    \sb_0__1__2_chany_bottom_out[7] ,
    \sb_0__1__2_chany_bottom_out[8] ,
    \sb_0__1__2_chany_bottom_out[9] ,
    \sb_0__1__2_chany_bottom_out[10] ,
    \sb_0__1__2_chany_bottom_out[11] ,
    \sb_0__1__2_chany_bottom_out[12] ,
    \sb_0__1__2_chany_bottom_out[13] ,
    \sb_0__1__2_chany_bottom_out[14] ,
    \sb_0__1__2_chany_bottom_out[15] ,
    \sb_0__1__2_chany_bottom_out[16] ,
    \sb_0__1__2_chany_bottom_out[17] ,
    \sb_0__1__2_chany_bottom_out[18] ,
    \sb_0__1__2_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__2_chany_top_out[0] ,
    \cby_0__1__2_chany_top_out[1] ,
    \cby_0__1__2_chany_top_out[2] ,
    \cby_0__1__2_chany_top_out[3] ,
    \cby_0__1__2_chany_top_out[4] ,
    \cby_0__1__2_chany_top_out[5] ,
    \cby_0__1__2_chany_top_out[6] ,
    \cby_0__1__2_chany_top_out[7] ,
    \cby_0__1__2_chany_top_out[8] ,
    \cby_0__1__2_chany_top_out[9] ,
    \cby_0__1__2_chany_top_out[10] ,
    \cby_0__1__2_chany_top_out[11] ,
    \cby_0__1__2_chany_top_out[12] ,
    \cby_0__1__2_chany_top_out[13] ,
    \cby_0__1__2_chany_top_out[14] ,
    \cby_0__1__2_chany_top_out[15] ,
    \cby_0__1__2_chany_top_out[16] ,
    \cby_0__1__2_chany_top_out[17] ,
    \cby_0__1__2_chany_top_out[18] ,
    \cby_0__1__2_chany_top_out[19] }));
 cby_0__1_ cby_0__4_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__1__3_ccff_tail),
    .ccff_tail(grid_io_left_3_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]),
    .left_grid_pin_0_(cby_0__1__3_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[19] ),
    .right_width_0_height_0__pin_0_(cby_0__1__3_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_3_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_3_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__1__2_chany_top_out[0] ,
    \sb_0__1__2_chany_top_out[1] ,
    \sb_0__1__2_chany_top_out[2] ,
    \sb_0__1__2_chany_top_out[3] ,
    \sb_0__1__2_chany_top_out[4] ,
    \sb_0__1__2_chany_top_out[5] ,
    \sb_0__1__2_chany_top_out[6] ,
    \sb_0__1__2_chany_top_out[7] ,
    \sb_0__1__2_chany_top_out[8] ,
    \sb_0__1__2_chany_top_out[9] ,
    \sb_0__1__2_chany_top_out[10] ,
    \sb_0__1__2_chany_top_out[11] ,
    \sb_0__1__2_chany_top_out[12] ,
    \sb_0__1__2_chany_top_out[13] ,
    \sb_0__1__2_chany_top_out[14] ,
    \sb_0__1__2_chany_top_out[15] ,
    \sb_0__1__2_chany_top_out[16] ,
    \sb_0__1__2_chany_top_out[17] ,
    \sb_0__1__2_chany_top_out[18] ,
    \sb_0__1__2_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__3_chany_bottom_out[0] ,
    \cby_0__1__3_chany_bottom_out[1] ,
    \cby_0__1__3_chany_bottom_out[2] ,
    \cby_0__1__3_chany_bottom_out[3] ,
    \cby_0__1__3_chany_bottom_out[4] ,
    \cby_0__1__3_chany_bottom_out[5] ,
    \cby_0__1__3_chany_bottom_out[6] ,
    \cby_0__1__3_chany_bottom_out[7] ,
    \cby_0__1__3_chany_bottom_out[8] ,
    \cby_0__1__3_chany_bottom_out[9] ,
    \cby_0__1__3_chany_bottom_out[10] ,
    \cby_0__1__3_chany_bottom_out[11] ,
    \cby_0__1__3_chany_bottom_out[12] ,
    \cby_0__1__3_chany_bottom_out[13] ,
    \cby_0__1__3_chany_bottom_out[14] ,
    \cby_0__1__3_chany_bottom_out[15] ,
    \cby_0__1__3_chany_bottom_out[16] ,
    \cby_0__1__3_chany_bottom_out[17] ,
    \cby_0__1__3_chany_bottom_out[18] ,
    \cby_0__1__3_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__1__3_chany_bottom_out[0] ,
    \sb_0__1__3_chany_bottom_out[1] ,
    \sb_0__1__3_chany_bottom_out[2] ,
    \sb_0__1__3_chany_bottom_out[3] ,
    \sb_0__1__3_chany_bottom_out[4] ,
    \sb_0__1__3_chany_bottom_out[5] ,
    \sb_0__1__3_chany_bottom_out[6] ,
    \sb_0__1__3_chany_bottom_out[7] ,
    \sb_0__1__3_chany_bottom_out[8] ,
    \sb_0__1__3_chany_bottom_out[9] ,
    \sb_0__1__3_chany_bottom_out[10] ,
    \sb_0__1__3_chany_bottom_out[11] ,
    \sb_0__1__3_chany_bottom_out[12] ,
    \sb_0__1__3_chany_bottom_out[13] ,
    \sb_0__1__3_chany_bottom_out[14] ,
    \sb_0__1__3_chany_bottom_out[15] ,
    \sb_0__1__3_chany_bottom_out[16] ,
    \sb_0__1__3_chany_bottom_out[17] ,
    \sb_0__1__3_chany_bottom_out[18] ,
    \sb_0__1__3_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__3_chany_top_out[0] ,
    \cby_0__1__3_chany_top_out[1] ,
    \cby_0__1__3_chany_top_out[2] ,
    \cby_0__1__3_chany_top_out[3] ,
    \cby_0__1__3_chany_top_out[4] ,
    \cby_0__1__3_chany_top_out[5] ,
    \cby_0__1__3_chany_top_out[6] ,
    \cby_0__1__3_chany_top_out[7] ,
    \cby_0__1__3_chany_top_out[8] ,
    \cby_0__1__3_chany_top_out[9] ,
    \cby_0__1__3_chany_top_out[10] ,
    \cby_0__1__3_chany_top_out[11] ,
    \cby_0__1__3_chany_top_out[12] ,
    \cby_0__1__3_chany_top_out[13] ,
    \cby_0__1__3_chany_top_out[14] ,
    \cby_0__1__3_chany_top_out[15] ,
    \cby_0__1__3_chany_top_out[16] ,
    \cby_0__1__3_chany_top_out[17] ,
    \cby_0__1__3_chany_top_out[18] ,
    \cby_0__1__3_chany_top_out[19] }));
 cby_0__1_ cby_0__5_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__1__4_ccff_tail),
    .ccff_tail(grid_io_left_4_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]),
    .left_grid_pin_0_(cby_0__1__4_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[24] ),
    .right_width_0_height_0__pin_0_(cby_0__1__4_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_4_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_4_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__1__3_chany_top_out[0] ,
    \sb_0__1__3_chany_top_out[1] ,
    \sb_0__1__3_chany_top_out[2] ,
    \sb_0__1__3_chany_top_out[3] ,
    \sb_0__1__3_chany_top_out[4] ,
    \sb_0__1__3_chany_top_out[5] ,
    \sb_0__1__3_chany_top_out[6] ,
    \sb_0__1__3_chany_top_out[7] ,
    \sb_0__1__3_chany_top_out[8] ,
    \sb_0__1__3_chany_top_out[9] ,
    \sb_0__1__3_chany_top_out[10] ,
    \sb_0__1__3_chany_top_out[11] ,
    \sb_0__1__3_chany_top_out[12] ,
    \sb_0__1__3_chany_top_out[13] ,
    \sb_0__1__3_chany_top_out[14] ,
    \sb_0__1__3_chany_top_out[15] ,
    \sb_0__1__3_chany_top_out[16] ,
    \sb_0__1__3_chany_top_out[17] ,
    \sb_0__1__3_chany_top_out[18] ,
    \sb_0__1__3_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__4_chany_bottom_out[0] ,
    \cby_0__1__4_chany_bottom_out[1] ,
    \cby_0__1__4_chany_bottom_out[2] ,
    \cby_0__1__4_chany_bottom_out[3] ,
    \cby_0__1__4_chany_bottom_out[4] ,
    \cby_0__1__4_chany_bottom_out[5] ,
    \cby_0__1__4_chany_bottom_out[6] ,
    \cby_0__1__4_chany_bottom_out[7] ,
    \cby_0__1__4_chany_bottom_out[8] ,
    \cby_0__1__4_chany_bottom_out[9] ,
    \cby_0__1__4_chany_bottom_out[10] ,
    \cby_0__1__4_chany_bottom_out[11] ,
    \cby_0__1__4_chany_bottom_out[12] ,
    \cby_0__1__4_chany_bottom_out[13] ,
    \cby_0__1__4_chany_bottom_out[14] ,
    \cby_0__1__4_chany_bottom_out[15] ,
    \cby_0__1__4_chany_bottom_out[16] ,
    \cby_0__1__4_chany_bottom_out[17] ,
    \cby_0__1__4_chany_bottom_out[18] ,
    \cby_0__1__4_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__1__4_chany_bottom_out[0] ,
    \sb_0__1__4_chany_bottom_out[1] ,
    \sb_0__1__4_chany_bottom_out[2] ,
    \sb_0__1__4_chany_bottom_out[3] ,
    \sb_0__1__4_chany_bottom_out[4] ,
    \sb_0__1__4_chany_bottom_out[5] ,
    \sb_0__1__4_chany_bottom_out[6] ,
    \sb_0__1__4_chany_bottom_out[7] ,
    \sb_0__1__4_chany_bottom_out[8] ,
    \sb_0__1__4_chany_bottom_out[9] ,
    \sb_0__1__4_chany_bottom_out[10] ,
    \sb_0__1__4_chany_bottom_out[11] ,
    \sb_0__1__4_chany_bottom_out[12] ,
    \sb_0__1__4_chany_bottom_out[13] ,
    \sb_0__1__4_chany_bottom_out[14] ,
    \sb_0__1__4_chany_bottom_out[15] ,
    \sb_0__1__4_chany_bottom_out[16] ,
    \sb_0__1__4_chany_bottom_out[17] ,
    \sb_0__1__4_chany_bottom_out[18] ,
    \sb_0__1__4_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__4_chany_top_out[0] ,
    \cby_0__1__4_chany_top_out[1] ,
    \cby_0__1__4_chany_top_out[2] ,
    \cby_0__1__4_chany_top_out[3] ,
    \cby_0__1__4_chany_top_out[4] ,
    \cby_0__1__4_chany_top_out[5] ,
    \cby_0__1__4_chany_top_out[6] ,
    \cby_0__1__4_chany_top_out[7] ,
    \cby_0__1__4_chany_top_out[8] ,
    \cby_0__1__4_chany_top_out[9] ,
    \cby_0__1__4_chany_top_out[10] ,
    \cby_0__1__4_chany_top_out[11] ,
    \cby_0__1__4_chany_top_out[12] ,
    \cby_0__1__4_chany_top_out[13] ,
    \cby_0__1__4_chany_top_out[14] ,
    \cby_0__1__4_chany_top_out[15] ,
    \cby_0__1__4_chany_top_out[16] ,
    \cby_0__1__4_chany_top_out[17] ,
    \cby_0__1__4_chany_top_out[18] ,
    \cby_0__1__4_chany_top_out[19] }));
 cby_0__1_ cby_0__6_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__1__5_ccff_tail),
    .ccff_tail(grid_io_left_5_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]),
    .left_grid_pin_0_(cby_0__1__5_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[29] ),
    .right_width_0_height_0__pin_0_(cby_0__1__5_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_5_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_5_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__1__4_chany_top_out[0] ,
    \sb_0__1__4_chany_top_out[1] ,
    \sb_0__1__4_chany_top_out[2] ,
    \sb_0__1__4_chany_top_out[3] ,
    \sb_0__1__4_chany_top_out[4] ,
    \sb_0__1__4_chany_top_out[5] ,
    \sb_0__1__4_chany_top_out[6] ,
    \sb_0__1__4_chany_top_out[7] ,
    \sb_0__1__4_chany_top_out[8] ,
    \sb_0__1__4_chany_top_out[9] ,
    \sb_0__1__4_chany_top_out[10] ,
    \sb_0__1__4_chany_top_out[11] ,
    \sb_0__1__4_chany_top_out[12] ,
    \sb_0__1__4_chany_top_out[13] ,
    \sb_0__1__4_chany_top_out[14] ,
    \sb_0__1__4_chany_top_out[15] ,
    \sb_0__1__4_chany_top_out[16] ,
    \sb_0__1__4_chany_top_out[17] ,
    \sb_0__1__4_chany_top_out[18] ,
    \sb_0__1__4_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__5_chany_bottom_out[0] ,
    \cby_0__1__5_chany_bottom_out[1] ,
    \cby_0__1__5_chany_bottom_out[2] ,
    \cby_0__1__5_chany_bottom_out[3] ,
    \cby_0__1__5_chany_bottom_out[4] ,
    \cby_0__1__5_chany_bottom_out[5] ,
    \cby_0__1__5_chany_bottom_out[6] ,
    \cby_0__1__5_chany_bottom_out[7] ,
    \cby_0__1__5_chany_bottom_out[8] ,
    \cby_0__1__5_chany_bottom_out[9] ,
    \cby_0__1__5_chany_bottom_out[10] ,
    \cby_0__1__5_chany_bottom_out[11] ,
    \cby_0__1__5_chany_bottom_out[12] ,
    \cby_0__1__5_chany_bottom_out[13] ,
    \cby_0__1__5_chany_bottom_out[14] ,
    \cby_0__1__5_chany_bottom_out[15] ,
    \cby_0__1__5_chany_bottom_out[16] ,
    \cby_0__1__5_chany_bottom_out[17] ,
    \cby_0__1__5_chany_bottom_out[18] ,
    \cby_0__1__5_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__1__5_chany_bottom_out[0] ,
    \sb_0__1__5_chany_bottom_out[1] ,
    \sb_0__1__5_chany_bottom_out[2] ,
    \sb_0__1__5_chany_bottom_out[3] ,
    \sb_0__1__5_chany_bottom_out[4] ,
    \sb_0__1__5_chany_bottom_out[5] ,
    \sb_0__1__5_chany_bottom_out[6] ,
    \sb_0__1__5_chany_bottom_out[7] ,
    \sb_0__1__5_chany_bottom_out[8] ,
    \sb_0__1__5_chany_bottom_out[9] ,
    \sb_0__1__5_chany_bottom_out[10] ,
    \sb_0__1__5_chany_bottom_out[11] ,
    \sb_0__1__5_chany_bottom_out[12] ,
    \sb_0__1__5_chany_bottom_out[13] ,
    \sb_0__1__5_chany_bottom_out[14] ,
    \sb_0__1__5_chany_bottom_out[15] ,
    \sb_0__1__5_chany_bottom_out[16] ,
    \sb_0__1__5_chany_bottom_out[17] ,
    \sb_0__1__5_chany_bottom_out[18] ,
    \sb_0__1__5_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__5_chany_top_out[0] ,
    \cby_0__1__5_chany_top_out[1] ,
    \cby_0__1__5_chany_top_out[2] ,
    \cby_0__1__5_chany_top_out[3] ,
    \cby_0__1__5_chany_top_out[4] ,
    \cby_0__1__5_chany_top_out[5] ,
    \cby_0__1__5_chany_top_out[6] ,
    \cby_0__1__5_chany_top_out[7] ,
    \cby_0__1__5_chany_top_out[8] ,
    \cby_0__1__5_chany_top_out[9] ,
    \cby_0__1__5_chany_top_out[10] ,
    \cby_0__1__5_chany_top_out[11] ,
    \cby_0__1__5_chany_top_out[12] ,
    \cby_0__1__5_chany_top_out[13] ,
    \cby_0__1__5_chany_top_out[14] ,
    \cby_0__1__5_chany_top_out[15] ,
    \cby_0__1__5_chany_top_out[16] ,
    \cby_0__1__5_chany_top_out[17] ,
    \cby_0__1__5_chany_top_out[18] ,
    \cby_0__1__5_chany_top_out[19] }));
 cby_0__1_ cby_0__7_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__1__6_ccff_tail),
    .ccff_tail(grid_io_left_6_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]),
    .left_grid_pin_0_(cby_0__1__6_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[34] ),
    .right_width_0_height_0__pin_0_(cby_0__1__6_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_6_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_6_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__1__5_chany_top_out[0] ,
    \sb_0__1__5_chany_top_out[1] ,
    \sb_0__1__5_chany_top_out[2] ,
    \sb_0__1__5_chany_top_out[3] ,
    \sb_0__1__5_chany_top_out[4] ,
    \sb_0__1__5_chany_top_out[5] ,
    \sb_0__1__5_chany_top_out[6] ,
    \sb_0__1__5_chany_top_out[7] ,
    \sb_0__1__5_chany_top_out[8] ,
    \sb_0__1__5_chany_top_out[9] ,
    \sb_0__1__5_chany_top_out[10] ,
    \sb_0__1__5_chany_top_out[11] ,
    \sb_0__1__5_chany_top_out[12] ,
    \sb_0__1__5_chany_top_out[13] ,
    \sb_0__1__5_chany_top_out[14] ,
    \sb_0__1__5_chany_top_out[15] ,
    \sb_0__1__5_chany_top_out[16] ,
    \sb_0__1__5_chany_top_out[17] ,
    \sb_0__1__5_chany_top_out[18] ,
    \sb_0__1__5_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__6_chany_bottom_out[0] ,
    \cby_0__1__6_chany_bottom_out[1] ,
    \cby_0__1__6_chany_bottom_out[2] ,
    \cby_0__1__6_chany_bottom_out[3] ,
    \cby_0__1__6_chany_bottom_out[4] ,
    \cby_0__1__6_chany_bottom_out[5] ,
    \cby_0__1__6_chany_bottom_out[6] ,
    \cby_0__1__6_chany_bottom_out[7] ,
    \cby_0__1__6_chany_bottom_out[8] ,
    \cby_0__1__6_chany_bottom_out[9] ,
    \cby_0__1__6_chany_bottom_out[10] ,
    \cby_0__1__6_chany_bottom_out[11] ,
    \cby_0__1__6_chany_bottom_out[12] ,
    \cby_0__1__6_chany_bottom_out[13] ,
    \cby_0__1__6_chany_bottom_out[14] ,
    \cby_0__1__6_chany_bottom_out[15] ,
    \cby_0__1__6_chany_bottom_out[16] ,
    \cby_0__1__6_chany_bottom_out[17] ,
    \cby_0__1__6_chany_bottom_out[18] ,
    \cby_0__1__6_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__1__6_chany_bottom_out[0] ,
    \sb_0__1__6_chany_bottom_out[1] ,
    \sb_0__1__6_chany_bottom_out[2] ,
    \sb_0__1__6_chany_bottom_out[3] ,
    \sb_0__1__6_chany_bottom_out[4] ,
    \sb_0__1__6_chany_bottom_out[5] ,
    \sb_0__1__6_chany_bottom_out[6] ,
    \sb_0__1__6_chany_bottom_out[7] ,
    \sb_0__1__6_chany_bottom_out[8] ,
    \sb_0__1__6_chany_bottom_out[9] ,
    \sb_0__1__6_chany_bottom_out[10] ,
    \sb_0__1__6_chany_bottom_out[11] ,
    \sb_0__1__6_chany_bottom_out[12] ,
    \sb_0__1__6_chany_bottom_out[13] ,
    \sb_0__1__6_chany_bottom_out[14] ,
    \sb_0__1__6_chany_bottom_out[15] ,
    \sb_0__1__6_chany_bottom_out[16] ,
    \sb_0__1__6_chany_bottom_out[17] ,
    \sb_0__1__6_chany_bottom_out[18] ,
    \sb_0__1__6_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__6_chany_top_out[0] ,
    \cby_0__1__6_chany_top_out[1] ,
    \cby_0__1__6_chany_top_out[2] ,
    \cby_0__1__6_chany_top_out[3] ,
    \cby_0__1__6_chany_top_out[4] ,
    \cby_0__1__6_chany_top_out[5] ,
    \cby_0__1__6_chany_top_out[6] ,
    \cby_0__1__6_chany_top_out[7] ,
    \cby_0__1__6_chany_top_out[8] ,
    \cby_0__1__6_chany_top_out[9] ,
    \cby_0__1__6_chany_top_out[10] ,
    \cby_0__1__6_chany_top_out[11] ,
    \cby_0__1__6_chany_top_out[12] ,
    \cby_0__1__6_chany_top_out[13] ,
    \cby_0__1__6_chany_top_out[14] ,
    \cby_0__1__6_chany_top_out[15] ,
    \cby_0__1__6_chany_top_out[16] ,
    \cby_0__1__6_chany_top_out[17] ,
    \cby_0__1__6_chany_top_out[18] ,
    \cby_0__1__6_chany_top_out[19] }));
 cby_0__1_ cby_0__8_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(sb_0__8__0_ccff_tail),
    .ccff_tail(grid_io_left_7_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]),
    .left_grid_pin_0_(cby_0__1__7_left_grid_pin_0_),
    .prog_clk_0_E_in(\prog_clk_0_wires[41] ),
    .right_width_0_height_0__pin_0_(cby_0__1__7_left_grid_pin_0_),
    .right_width_0_height_0__pin_1_lower(grid_io_left_7_right_width_0_height_0__pin_1_lower),
    .right_width_0_height_0__pin_1_upper(grid_io_left_7_right_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_0__1__6_chany_top_out[0] ,
    \sb_0__1__6_chany_top_out[1] ,
    \sb_0__1__6_chany_top_out[2] ,
    \sb_0__1__6_chany_top_out[3] ,
    \sb_0__1__6_chany_top_out[4] ,
    \sb_0__1__6_chany_top_out[5] ,
    \sb_0__1__6_chany_top_out[6] ,
    \sb_0__1__6_chany_top_out[7] ,
    \sb_0__1__6_chany_top_out[8] ,
    \sb_0__1__6_chany_top_out[9] ,
    \sb_0__1__6_chany_top_out[10] ,
    \sb_0__1__6_chany_top_out[11] ,
    \sb_0__1__6_chany_top_out[12] ,
    \sb_0__1__6_chany_top_out[13] ,
    \sb_0__1__6_chany_top_out[14] ,
    \sb_0__1__6_chany_top_out[15] ,
    \sb_0__1__6_chany_top_out[16] ,
    \sb_0__1__6_chany_top_out[17] ,
    \sb_0__1__6_chany_top_out[18] ,
    \sb_0__1__6_chany_top_out[19] }),
    .chany_bottom_out({\cby_0__1__7_chany_bottom_out[0] ,
    \cby_0__1__7_chany_bottom_out[1] ,
    \cby_0__1__7_chany_bottom_out[2] ,
    \cby_0__1__7_chany_bottom_out[3] ,
    \cby_0__1__7_chany_bottom_out[4] ,
    \cby_0__1__7_chany_bottom_out[5] ,
    \cby_0__1__7_chany_bottom_out[6] ,
    \cby_0__1__7_chany_bottom_out[7] ,
    \cby_0__1__7_chany_bottom_out[8] ,
    \cby_0__1__7_chany_bottom_out[9] ,
    \cby_0__1__7_chany_bottom_out[10] ,
    \cby_0__1__7_chany_bottom_out[11] ,
    \cby_0__1__7_chany_bottom_out[12] ,
    \cby_0__1__7_chany_bottom_out[13] ,
    \cby_0__1__7_chany_bottom_out[14] ,
    \cby_0__1__7_chany_bottom_out[15] ,
    \cby_0__1__7_chany_bottom_out[16] ,
    \cby_0__1__7_chany_bottom_out[17] ,
    \cby_0__1__7_chany_bottom_out[18] ,
    \cby_0__1__7_chany_bottom_out[19] }),
    .chany_top_in({\sb_0__8__0_chany_bottom_out[0] ,
    \sb_0__8__0_chany_bottom_out[1] ,
    \sb_0__8__0_chany_bottom_out[2] ,
    \sb_0__8__0_chany_bottom_out[3] ,
    \sb_0__8__0_chany_bottom_out[4] ,
    \sb_0__8__0_chany_bottom_out[5] ,
    \sb_0__8__0_chany_bottom_out[6] ,
    \sb_0__8__0_chany_bottom_out[7] ,
    \sb_0__8__0_chany_bottom_out[8] ,
    \sb_0__8__0_chany_bottom_out[9] ,
    \sb_0__8__0_chany_bottom_out[10] ,
    \sb_0__8__0_chany_bottom_out[11] ,
    \sb_0__8__0_chany_bottom_out[12] ,
    \sb_0__8__0_chany_bottom_out[13] ,
    \sb_0__8__0_chany_bottom_out[14] ,
    \sb_0__8__0_chany_bottom_out[15] ,
    \sb_0__8__0_chany_bottom_out[16] ,
    \sb_0__8__0_chany_bottom_out[17] ,
    \sb_0__8__0_chany_bottom_out[18] ,
    \sb_0__8__0_chany_bottom_out[19] }),
    .chany_top_out({\cby_0__1__7_chany_top_out[0] ,
    \cby_0__1__7_chany_top_out[1] ,
    \cby_0__1__7_chany_top_out[2] ,
    \cby_0__1__7_chany_top_out[3] ,
    \cby_0__1__7_chany_top_out[4] ,
    \cby_0__1__7_chany_top_out[5] ,
    \cby_0__1__7_chany_top_out[6] ,
    \cby_0__1__7_chany_top_out[7] ,
    \cby_0__1__7_chany_top_out[8] ,
    \cby_0__1__7_chany_top_out[9] ,
    \cby_0__1__7_chany_top_out[10] ,
    \cby_0__1__7_chany_top_out[11] ,
    \cby_0__1__7_chany_top_out[12] ,
    \cby_0__1__7_chany_top_out[13] ,
    \cby_0__1__7_chany_top_out[14] ,
    \cby_0__1__7_chany_top_out[15] ,
    \cby_0__1__7_chany_top_out[16] ,
    \cby_0__1__7_chany_top_out[17] ,
    \cby_0__1__7_chany_top_out[18] ,
    \cby_0__1__7_chany_top_out[19] }));
 cby_1__1_ cby_1__1_ (.Test_en_E_in(\Test_enWires[18] ),
    .Test_en_S_in(\Test_enWires[18] ),
    .Test_en_W_in(\Test_enWires[18] ),
    .Test_en_W_out(\Test_enWires[16] ),
    .ccff_head(grid_clb_0_ccff_tail),
    .ccff_tail(cby_1__1__0_ccff_tail),
    .left_grid_pin_16_(cby_1__1__0_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__0_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__0_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__0_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__0_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__0_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__0_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__0_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__0_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__0_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__0_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__0_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__0_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__0_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__0_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__0_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[2] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[1] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__0__0_chany_top_out[0] ,
    \sb_1__0__0_chany_top_out[1] ,
    \sb_1__0__0_chany_top_out[2] ,
    \sb_1__0__0_chany_top_out[3] ,
    \sb_1__0__0_chany_top_out[4] ,
    \sb_1__0__0_chany_top_out[5] ,
    \sb_1__0__0_chany_top_out[6] ,
    \sb_1__0__0_chany_top_out[7] ,
    \sb_1__0__0_chany_top_out[8] ,
    \sb_1__0__0_chany_top_out[9] ,
    \sb_1__0__0_chany_top_out[10] ,
    \sb_1__0__0_chany_top_out[11] ,
    \sb_1__0__0_chany_top_out[12] ,
    \sb_1__0__0_chany_top_out[13] ,
    \sb_1__0__0_chany_top_out[14] ,
    \sb_1__0__0_chany_top_out[15] ,
    \sb_1__0__0_chany_top_out[16] ,
    \sb_1__0__0_chany_top_out[17] ,
    \sb_1__0__0_chany_top_out[18] ,
    \sb_1__0__0_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__0_chany_bottom_out[0] ,
    \cby_1__1__0_chany_bottom_out[1] ,
    \cby_1__1__0_chany_bottom_out[2] ,
    \cby_1__1__0_chany_bottom_out[3] ,
    \cby_1__1__0_chany_bottom_out[4] ,
    \cby_1__1__0_chany_bottom_out[5] ,
    \cby_1__1__0_chany_bottom_out[6] ,
    \cby_1__1__0_chany_bottom_out[7] ,
    \cby_1__1__0_chany_bottom_out[8] ,
    \cby_1__1__0_chany_bottom_out[9] ,
    \cby_1__1__0_chany_bottom_out[10] ,
    \cby_1__1__0_chany_bottom_out[11] ,
    \cby_1__1__0_chany_bottom_out[12] ,
    \cby_1__1__0_chany_bottom_out[13] ,
    \cby_1__1__0_chany_bottom_out[14] ,
    \cby_1__1__0_chany_bottom_out[15] ,
    \cby_1__1__0_chany_bottom_out[16] ,
    \cby_1__1__0_chany_bottom_out[17] ,
    \cby_1__1__0_chany_bottom_out[18] ,
    \cby_1__1__0_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__0_chany_bottom_out[0] ,
    \sb_1__1__0_chany_bottom_out[1] ,
    \sb_1__1__0_chany_bottom_out[2] ,
    \sb_1__1__0_chany_bottom_out[3] ,
    \sb_1__1__0_chany_bottom_out[4] ,
    \sb_1__1__0_chany_bottom_out[5] ,
    \sb_1__1__0_chany_bottom_out[6] ,
    \sb_1__1__0_chany_bottom_out[7] ,
    \sb_1__1__0_chany_bottom_out[8] ,
    \sb_1__1__0_chany_bottom_out[9] ,
    \sb_1__1__0_chany_bottom_out[10] ,
    \sb_1__1__0_chany_bottom_out[11] ,
    \sb_1__1__0_chany_bottom_out[12] ,
    \sb_1__1__0_chany_bottom_out[13] ,
    \sb_1__1__0_chany_bottom_out[14] ,
    \sb_1__1__0_chany_bottom_out[15] ,
    \sb_1__1__0_chany_bottom_out[16] ,
    \sb_1__1__0_chany_bottom_out[17] ,
    \sb_1__1__0_chany_bottom_out[18] ,
    \sb_1__1__0_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__0_chany_top_out[0] ,
    \cby_1__1__0_chany_top_out[1] ,
    \cby_1__1__0_chany_top_out[2] ,
    \cby_1__1__0_chany_top_out[3] ,
    \cby_1__1__0_chany_top_out[4] ,
    \cby_1__1__0_chany_top_out[5] ,
    \cby_1__1__0_chany_top_out[6] ,
    \cby_1__1__0_chany_top_out[7] ,
    \cby_1__1__0_chany_top_out[8] ,
    \cby_1__1__0_chany_top_out[9] ,
    \cby_1__1__0_chany_top_out[10] ,
    \cby_1__1__0_chany_top_out[11] ,
    \cby_1__1__0_chany_top_out[12] ,
    \cby_1__1__0_chany_top_out[13] ,
    \cby_1__1__0_chany_top_out[14] ,
    \cby_1__1__0_chany_top_out[15] ,
    \cby_1__1__0_chany_top_out[16] ,
    \cby_1__1__0_chany_top_out[17] ,
    \cby_1__1__0_chany_top_out[18] ,
    \cby_1__1__0_chany_top_out[19] }));
 cby_1__1_ cby_1__2_ (.Test_en_E_in(\Test_enWires[32] ),
    .Test_en_S_in(\Test_enWires[32] ),
    .Test_en_W_in(\Test_enWires[32] ),
    .Test_en_W_out(\Test_enWires[30] ),
    .ccff_head(grid_clb_1_ccff_tail),
    .ccff_tail(cby_1__1__1_ccff_tail),
    .clk_2_S_in(\clk_2_wires[7] ),
    .clk_2_S_out(\clk_2_wires[8] ),
    .left_grid_pin_16_(cby_1__1__1_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__1_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__1_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__1_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__1_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__1_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__1_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__1_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__1_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__1_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__1_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__1_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__1_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__1_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__1_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__1_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[8] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[7] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[7] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[8] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__0_chany_top_out[0] ,
    \sb_1__1__0_chany_top_out[1] ,
    \sb_1__1__0_chany_top_out[2] ,
    \sb_1__1__0_chany_top_out[3] ,
    \sb_1__1__0_chany_top_out[4] ,
    \sb_1__1__0_chany_top_out[5] ,
    \sb_1__1__0_chany_top_out[6] ,
    \sb_1__1__0_chany_top_out[7] ,
    \sb_1__1__0_chany_top_out[8] ,
    \sb_1__1__0_chany_top_out[9] ,
    \sb_1__1__0_chany_top_out[10] ,
    \sb_1__1__0_chany_top_out[11] ,
    \sb_1__1__0_chany_top_out[12] ,
    \sb_1__1__0_chany_top_out[13] ,
    \sb_1__1__0_chany_top_out[14] ,
    \sb_1__1__0_chany_top_out[15] ,
    \sb_1__1__0_chany_top_out[16] ,
    \sb_1__1__0_chany_top_out[17] ,
    \sb_1__1__0_chany_top_out[18] ,
    \sb_1__1__0_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__1_chany_bottom_out[0] ,
    \cby_1__1__1_chany_bottom_out[1] ,
    \cby_1__1__1_chany_bottom_out[2] ,
    \cby_1__1__1_chany_bottom_out[3] ,
    \cby_1__1__1_chany_bottom_out[4] ,
    \cby_1__1__1_chany_bottom_out[5] ,
    \cby_1__1__1_chany_bottom_out[6] ,
    \cby_1__1__1_chany_bottom_out[7] ,
    \cby_1__1__1_chany_bottom_out[8] ,
    \cby_1__1__1_chany_bottom_out[9] ,
    \cby_1__1__1_chany_bottom_out[10] ,
    \cby_1__1__1_chany_bottom_out[11] ,
    \cby_1__1__1_chany_bottom_out[12] ,
    \cby_1__1__1_chany_bottom_out[13] ,
    \cby_1__1__1_chany_bottom_out[14] ,
    \cby_1__1__1_chany_bottom_out[15] ,
    \cby_1__1__1_chany_bottom_out[16] ,
    \cby_1__1__1_chany_bottom_out[17] ,
    \cby_1__1__1_chany_bottom_out[18] ,
    \cby_1__1__1_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__1_chany_bottom_out[0] ,
    \sb_1__1__1_chany_bottom_out[1] ,
    \sb_1__1__1_chany_bottom_out[2] ,
    \sb_1__1__1_chany_bottom_out[3] ,
    \sb_1__1__1_chany_bottom_out[4] ,
    \sb_1__1__1_chany_bottom_out[5] ,
    \sb_1__1__1_chany_bottom_out[6] ,
    \sb_1__1__1_chany_bottom_out[7] ,
    \sb_1__1__1_chany_bottom_out[8] ,
    \sb_1__1__1_chany_bottom_out[9] ,
    \sb_1__1__1_chany_bottom_out[10] ,
    \sb_1__1__1_chany_bottom_out[11] ,
    \sb_1__1__1_chany_bottom_out[12] ,
    \sb_1__1__1_chany_bottom_out[13] ,
    \sb_1__1__1_chany_bottom_out[14] ,
    \sb_1__1__1_chany_bottom_out[15] ,
    \sb_1__1__1_chany_bottom_out[16] ,
    \sb_1__1__1_chany_bottom_out[17] ,
    \sb_1__1__1_chany_bottom_out[18] ,
    \sb_1__1__1_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__1_chany_top_out[0] ,
    \cby_1__1__1_chany_top_out[1] ,
    \cby_1__1__1_chany_top_out[2] ,
    \cby_1__1__1_chany_top_out[3] ,
    \cby_1__1__1_chany_top_out[4] ,
    \cby_1__1__1_chany_top_out[5] ,
    \cby_1__1__1_chany_top_out[6] ,
    \cby_1__1__1_chany_top_out[7] ,
    \cby_1__1__1_chany_top_out[8] ,
    \cby_1__1__1_chany_top_out[9] ,
    \cby_1__1__1_chany_top_out[10] ,
    \cby_1__1__1_chany_top_out[11] ,
    \cby_1__1__1_chany_top_out[12] ,
    \cby_1__1__1_chany_top_out[13] ,
    \cby_1__1__1_chany_top_out[14] ,
    \cby_1__1__1_chany_top_out[15] ,
    \cby_1__1__1_chany_top_out[16] ,
    \cby_1__1__1_chany_top_out[17] ,
    \cby_1__1__1_chany_top_out[18] ,
    \cby_1__1__1_chany_top_out[19] }));
 cby_1__1_ cby_1__3_ (.Test_en_E_in(\Test_enWires[46] ),
    .Test_en_S_in(\Test_enWires[46] ),
    .Test_en_W_in(\Test_enWires[46] ),
    .Test_en_W_out(\Test_enWires[44] ),
    .ccff_head(grid_clb_2_ccff_tail),
    .ccff_tail(cby_1__1__2_ccff_tail),
    .clk_2_N_out(\clk_2_wires[6] ),
    .clk_2_S_in(\clk_2_wires[5] ),
    .left_grid_pin_16_(cby_1__1__2_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__2_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__2_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__2_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__2_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__2_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__2_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__2_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__2_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__2_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__2_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__2_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__2_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__2_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__2_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__2_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[13] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[12] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[6] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[5] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__1_chany_top_out[0] ,
    \sb_1__1__1_chany_top_out[1] ,
    \sb_1__1__1_chany_top_out[2] ,
    \sb_1__1__1_chany_top_out[3] ,
    \sb_1__1__1_chany_top_out[4] ,
    \sb_1__1__1_chany_top_out[5] ,
    \sb_1__1__1_chany_top_out[6] ,
    \sb_1__1__1_chany_top_out[7] ,
    \sb_1__1__1_chany_top_out[8] ,
    \sb_1__1__1_chany_top_out[9] ,
    \sb_1__1__1_chany_top_out[10] ,
    \sb_1__1__1_chany_top_out[11] ,
    \sb_1__1__1_chany_top_out[12] ,
    \sb_1__1__1_chany_top_out[13] ,
    \sb_1__1__1_chany_top_out[14] ,
    \sb_1__1__1_chany_top_out[15] ,
    \sb_1__1__1_chany_top_out[16] ,
    \sb_1__1__1_chany_top_out[17] ,
    \sb_1__1__1_chany_top_out[18] ,
    \sb_1__1__1_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__2_chany_bottom_out[0] ,
    \cby_1__1__2_chany_bottom_out[1] ,
    \cby_1__1__2_chany_bottom_out[2] ,
    \cby_1__1__2_chany_bottom_out[3] ,
    \cby_1__1__2_chany_bottom_out[4] ,
    \cby_1__1__2_chany_bottom_out[5] ,
    \cby_1__1__2_chany_bottom_out[6] ,
    \cby_1__1__2_chany_bottom_out[7] ,
    \cby_1__1__2_chany_bottom_out[8] ,
    \cby_1__1__2_chany_bottom_out[9] ,
    \cby_1__1__2_chany_bottom_out[10] ,
    \cby_1__1__2_chany_bottom_out[11] ,
    \cby_1__1__2_chany_bottom_out[12] ,
    \cby_1__1__2_chany_bottom_out[13] ,
    \cby_1__1__2_chany_bottom_out[14] ,
    \cby_1__1__2_chany_bottom_out[15] ,
    \cby_1__1__2_chany_bottom_out[16] ,
    \cby_1__1__2_chany_bottom_out[17] ,
    \cby_1__1__2_chany_bottom_out[18] ,
    \cby_1__1__2_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__2_chany_bottom_out[0] ,
    \sb_1__1__2_chany_bottom_out[1] ,
    \sb_1__1__2_chany_bottom_out[2] ,
    \sb_1__1__2_chany_bottom_out[3] ,
    \sb_1__1__2_chany_bottom_out[4] ,
    \sb_1__1__2_chany_bottom_out[5] ,
    \sb_1__1__2_chany_bottom_out[6] ,
    \sb_1__1__2_chany_bottom_out[7] ,
    \sb_1__1__2_chany_bottom_out[8] ,
    \sb_1__1__2_chany_bottom_out[9] ,
    \sb_1__1__2_chany_bottom_out[10] ,
    \sb_1__1__2_chany_bottom_out[11] ,
    \sb_1__1__2_chany_bottom_out[12] ,
    \sb_1__1__2_chany_bottom_out[13] ,
    \sb_1__1__2_chany_bottom_out[14] ,
    \sb_1__1__2_chany_bottom_out[15] ,
    \sb_1__1__2_chany_bottom_out[16] ,
    \sb_1__1__2_chany_bottom_out[17] ,
    \sb_1__1__2_chany_bottom_out[18] ,
    \sb_1__1__2_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__2_chany_top_out[0] ,
    \cby_1__1__2_chany_top_out[1] ,
    \cby_1__1__2_chany_top_out[2] ,
    \cby_1__1__2_chany_top_out[3] ,
    \cby_1__1__2_chany_top_out[4] ,
    \cby_1__1__2_chany_top_out[5] ,
    \cby_1__1__2_chany_top_out[6] ,
    \cby_1__1__2_chany_top_out[7] ,
    \cby_1__1__2_chany_top_out[8] ,
    \cby_1__1__2_chany_top_out[9] ,
    \cby_1__1__2_chany_top_out[10] ,
    \cby_1__1__2_chany_top_out[11] ,
    \cby_1__1__2_chany_top_out[12] ,
    \cby_1__1__2_chany_top_out[13] ,
    \cby_1__1__2_chany_top_out[14] ,
    \cby_1__1__2_chany_top_out[15] ,
    \cby_1__1__2_chany_top_out[16] ,
    \cby_1__1__2_chany_top_out[17] ,
    \cby_1__1__2_chany_top_out[18] ,
    \cby_1__1__2_chany_top_out[19] }));
 cby_1__1_ cby_1__4_ (.Test_en_E_in(\Test_enWires[60] ),
    .Test_en_S_in(\Test_enWires[60] ),
    .Test_en_W_in(\Test_enWires[60] ),
    .Test_en_W_out(\Test_enWires[58] ),
    .ccff_head(grid_clb_3_ccff_tail),
    .ccff_tail(cby_1__1__3_ccff_tail),
    .left_grid_pin_16_(cby_1__1__3_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__3_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__3_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__3_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__3_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__3_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__3_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__3_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__3_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__3_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__3_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__3_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__3_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__3_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__3_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__3_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[18] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[17] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__2_chany_top_out[0] ,
    \sb_1__1__2_chany_top_out[1] ,
    \sb_1__1__2_chany_top_out[2] ,
    \sb_1__1__2_chany_top_out[3] ,
    \sb_1__1__2_chany_top_out[4] ,
    \sb_1__1__2_chany_top_out[5] ,
    \sb_1__1__2_chany_top_out[6] ,
    \sb_1__1__2_chany_top_out[7] ,
    \sb_1__1__2_chany_top_out[8] ,
    \sb_1__1__2_chany_top_out[9] ,
    \sb_1__1__2_chany_top_out[10] ,
    \sb_1__1__2_chany_top_out[11] ,
    \sb_1__1__2_chany_top_out[12] ,
    \sb_1__1__2_chany_top_out[13] ,
    \sb_1__1__2_chany_top_out[14] ,
    \sb_1__1__2_chany_top_out[15] ,
    \sb_1__1__2_chany_top_out[16] ,
    \sb_1__1__2_chany_top_out[17] ,
    \sb_1__1__2_chany_top_out[18] ,
    \sb_1__1__2_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__3_chany_bottom_out[0] ,
    \cby_1__1__3_chany_bottom_out[1] ,
    \cby_1__1__3_chany_bottom_out[2] ,
    \cby_1__1__3_chany_bottom_out[3] ,
    \cby_1__1__3_chany_bottom_out[4] ,
    \cby_1__1__3_chany_bottom_out[5] ,
    \cby_1__1__3_chany_bottom_out[6] ,
    \cby_1__1__3_chany_bottom_out[7] ,
    \cby_1__1__3_chany_bottom_out[8] ,
    \cby_1__1__3_chany_bottom_out[9] ,
    \cby_1__1__3_chany_bottom_out[10] ,
    \cby_1__1__3_chany_bottom_out[11] ,
    \cby_1__1__3_chany_bottom_out[12] ,
    \cby_1__1__3_chany_bottom_out[13] ,
    \cby_1__1__3_chany_bottom_out[14] ,
    \cby_1__1__3_chany_bottom_out[15] ,
    \cby_1__1__3_chany_bottom_out[16] ,
    \cby_1__1__3_chany_bottom_out[17] ,
    \cby_1__1__3_chany_bottom_out[18] ,
    \cby_1__1__3_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__3_chany_bottom_out[0] ,
    \sb_1__1__3_chany_bottom_out[1] ,
    \sb_1__1__3_chany_bottom_out[2] ,
    \sb_1__1__3_chany_bottom_out[3] ,
    \sb_1__1__3_chany_bottom_out[4] ,
    \sb_1__1__3_chany_bottom_out[5] ,
    \sb_1__1__3_chany_bottom_out[6] ,
    \sb_1__1__3_chany_bottom_out[7] ,
    \sb_1__1__3_chany_bottom_out[8] ,
    \sb_1__1__3_chany_bottom_out[9] ,
    \sb_1__1__3_chany_bottom_out[10] ,
    \sb_1__1__3_chany_bottom_out[11] ,
    \sb_1__1__3_chany_bottom_out[12] ,
    \sb_1__1__3_chany_bottom_out[13] ,
    \sb_1__1__3_chany_bottom_out[14] ,
    \sb_1__1__3_chany_bottom_out[15] ,
    \sb_1__1__3_chany_bottom_out[16] ,
    \sb_1__1__3_chany_bottom_out[17] ,
    \sb_1__1__3_chany_bottom_out[18] ,
    \sb_1__1__3_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__3_chany_top_out[0] ,
    \cby_1__1__3_chany_top_out[1] ,
    \cby_1__1__3_chany_top_out[2] ,
    \cby_1__1__3_chany_top_out[3] ,
    \cby_1__1__3_chany_top_out[4] ,
    \cby_1__1__3_chany_top_out[5] ,
    \cby_1__1__3_chany_top_out[6] ,
    \cby_1__1__3_chany_top_out[7] ,
    \cby_1__1__3_chany_top_out[8] ,
    \cby_1__1__3_chany_top_out[9] ,
    \cby_1__1__3_chany_top_out[10] ,
    \cby_1__1__3_chany_top_out[11] ,
    \cby_1__1__3_chany_top_out[12] ,
    \cby_1__1__3_chany_top_out[13] ,
    \cby_1__1__3_chany_top_out[14] ,
    \cby_1__1__3_chany_top_out[15] ,
    \cby_1__1__3_chany_top_out[16] ,
    \cby_1__1__3_chany_top_out[17] ,
    \cby_1__1__3_chany_top_out[18] ,
    \cby_1__1__3_chany_top_out[19] }));
 cby_1__1_ cby_1__5_ (.Test_en_E_in(\Test_enWires[74] ),
    .Test_en_S_in(\Test_enWires[74] ),
    .Test_en_W_in(\Test_enWires[74] ),
    .Test_en_W_out(\Test_enWires[72] ),
    .ccff_head(grid_clb_4_ccff_tail),
    .ccff_tail(cby_1__1__4_ccff_tail),
    .left_grid_pin_16_(cby_1__1__4_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__4_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__4_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__4_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__4_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__4_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__4_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__4_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__4_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__4_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__4_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__4_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__4_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__4_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__4_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__4_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[23] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[22] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__3_chany_top_out[0] ,
    \sb_1__1__3_chany_top_out[1] ,
    \sb_1__1__3_chany_top_out[2] ,
    \sb_1__1__3_chany_top_out[3] ,
    \sb_1__1__3_chany_top_out[4] ,
    \sb_1__1__3_chany_top_out[5] ,
    \sb_1__1__3_chany_top_out[6] ,
    \sb_1__1__3_chany_top_out[7] ,
    \sb_1__1__3_chany_top_out[8] ,
    \sb_1__1__3_chany_top_out[9] ,
    \sb_1__1__3_chany_top_out[10] ,
    \sb_1__1__3_chany_top_out[11] ,
    \sb_1__1__3_chany_top_out[12] ,
    \sb_1__1__3_chany_top_out[13] ,
    \sb_1__1__3_chany_top_out[14] ,
    \sb_1__1__3_chany_top_out[15] ,
    \sb_1__1__3_chany_top_out[16] ,
    \sb_1__1__3_chany_top_out[17] ,
    \sb_1__1__3_chany_top_out[18] ,
    \sb_1__1__3_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__4_chany_bottom_out[0] ,
    \cby_1__1__4_chany_bottom_out[1] ,
    \cby_1__1__4_chany_bottom_out[2] ,
    \cby_1__1__4_chany_bottom_out[3] ,
    \cby_1__1__4_chany_bottom_out[4] ,
    \cby_1__1__4_chany_bottom_out[5] ,
    \cby_1__1__4_chany_bottom_out[6] ,
    \cby_1__1__4_chany_bottom_out[7] ,
    \cby_1__1__4_chany_bottom_out[8] ,
    \cby_1__1__4_chany_bottom_out[9] ,
    \cby_1__1__4_chany_bottom_out[10] ,
    \cby_1__1__4_chany_bottom_out[11] ,
    \cby_1__1__4_chany_bottom_out[12] ,
    \cby_1__1__4_chany_bottom_out[13] ,
    \cby_1__1__4_chany_bottom_out[14] ,
    \cby_1__1__4_chany_bottom_out[15] ,
    \cby_1__1__4_chany_bottom_out[16] ,
    \cby_1__1__4_chany_bottom_out[17] ,
    \cby_1__1__4_chany_bottom_out[18] ,
    \cby_1__1__4_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__4_chany_bottom_out[0] ,
    \sb_1__1__4_chany_bottom_out[1] ,
    \sb_1__1__4_chany_bottom_out[2] ,
    \sb_1__1__4_chany_bottom_out[3] ,
    \sb_1__1__4_chany_bottom_out[4] ,
    \sb_1__1__4_chany_bottom_out[5] ,
    \sb_1__1__4_chany_bottom_out[6] ,
    \sb_1__1__4_chany_bottom_out[7] ,
    \sb_1__1__4_chany_bottom_out[8] ,
    \sb_1__1__4_chany_bottom_out[9] ,
    \sb_1__1__4_chany_bottom_out[10] ,
    \sb_1__1__4_chany_bottom_out[11] ,
    \sb_1__1__4_chany_bottom_out[12] ,
    \sb_1__1__4_chany_bottom_out[13] ,
    \sb_1__1__4_chany_bottom_out[14] ,
    \sb_1__1__4_chany_bottom_out[15] ,
    \sb_1__1__4_chany_bottom_out[16] ,
    \sb_1__1__4_chany_bottom_out[17] ,
    \sb_1__1__4_chany_bottom_out[18] ,
    \sb_1__1__4_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__4_chany_top_out[0] ,
    \cby_1__1__4_chany_top_out[1] ,
    \cby_1__1__4_chany_top_out[2] ,
    \cby_1__1__4_chany_top_out[3] ,
    \cby_1__1__4_chany_top_out[4] ,
    \cby_1__1__4_chany_top_out[5] ,
    \cby_1__1__4_chany_top_out[6] ,
    \cby_1__1__4_chany_top_out[7] ,
    \cby_1__1__4_chany_top_out[8] ,
    \cby_1__1__4_chany_top_out[9] ,
    \cby_1__1__4_chany_top_out[10] ,
    \cby_1__1__4_chany_top_out[11] ,
    \cby_1__1__4_chany_top_out[12] ,
    \cby_1__1__4_chany_top_out[13] ,
    \cby_1__1__4_chany_top_out[14] ,
    \cby_1__1__4_chany_top_out[15] ,
    \cby_1__1__4_chany_top_out[16] ,
    \cby_1__1__4_chany_top_out[17] ,
    \cby_1__1__4_chany_top_out[18] ,
    \cby_1__1__4_chany_top_out[19] }));
 cby_1__1_ cby_1__6_ (.Test_en_E_in(\Test_enWires[88] ),
    .Test_en_S_in(\Test_enWires[88] ),
    .Test_en_W_in(\Test_enWires[88] ),
    .Test_en_W_out(\Test_enWires[86] ),
    .ccff_head(grid_clb_5_ccff_tail),
    .ccff_tail(cby_1__1__5_ccff_tail),
    .clk_2_S_in(\clk_2_wires[20] ),
    .clk_2_S_out(\clk_2_wires[21] ),
    .left_grid_pin_16_(cby_1__1__5_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__5_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__5_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__5_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__5_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__5_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__5_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__5_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__5_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__5_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__5_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__5_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__5_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__5_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__5_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__5_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[28] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[27] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[20] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[21] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__4_chany_top_out[0] ,
    \sb_1__1__4_chany_top_out[1] ,
    \sb_1__1__4_chany_top_out[2] ,
    \sb_1__1__4_chany_top_out[3] ,
    \sb_1__1__4_chany_top_out[4] ,
    \sb_1__1__4_chany_top_out[5] ,
    \sb_1__1__4_chany_top_out[6] ,
    \sb_1__1__4_chany_top_out[7] ,
    \sb_1__1__4_chany_top_out[8] ,
    \sb_1__1__4_chany_top_out[9] ,
    \sb_1__1__4_chany_top_out[10] ,
    \sb_1__1__4_chany_top_out[11] ,
    \sb_1__1__4_chany_top_out[12] ,
    \sb_1__1__4_chany_top_out[13] ,
    \sb_1__1__4_chany_top_out[14] ,
    \sb_1__1__4_chany_top_out[15] ,
    \sb_1__1__4_chany_top_out[16] ,
    \sb_1__1__4_chany_top_out[17] ,
    \sb_1__1__4_chany_top_out[18] ,
    \sb_1__1__4_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__5_chany_bottom_out[0] ,
    \cby_1__1__5_chany_bottom_out[1] ,
    \cby_1__1__5_chany_bottom_out[2] ,
    \cby_1__1__5_chany_bottom_out[3] ,
    \cby_1__1__5_chany_bottom_out[4] ,
    \cby_1__1__5_chany_bottom_out[5] ,
    \cby_1__1__5_chany_bottom_out[6] ,
    \cby_1__1__5_chany_bottom_out[7] ,
    \cby_1__1__5_chany_bottom_out[8] ,
    \cby_1__1__5_chany_bottom_out[9] ,
    \cby_1__1__5_chany_bottom_out[10] ,
    \cby_1__1__5_chany_bottom_out[11] ,
    \cby_1__1__5_chany_bottom_out[12] ,
    \cby_1__1__5_chany_bottom_out[13] ,
    \cby_1__1__5_chany_bottom_out[14] ,
    \cby_1__1__5_chany_bottom_out[15] ,
    \cby_1__1__5_chany_bottom_out[16] ,
    \cby_1__1__5_chany_bottom_out[17] ,
    \cby_1__1__5_chany_bottom_out[18] ,
    \cby_1__1__5_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__5_chany_bottom_out[0] ,
    \sb_1__1__5_chany_bottom_out[1] ,
    \sb_1__1__5_chany_bottom_out[2] ,
    \sb_1__1__5_chany_bottom_out[3] ,
    \sb_1__1__5_chany_bottom_out[4] ,
    \sb_1__1__5_chany_bottom_out[5] ,
    \sb_1__1__5_chany_bottom_out[6] ,
    \sb_1__1__5_chany_bottom_out[7] ,
    \sb_1__1__5_chany_bottom_out[8] ,
    \sb_1__1__5_chany_bottom_out[9] ,
    \sb_1__1__5_chany_bottom_out[10] ,
    \sb_1__1__5_chany_bottom_out[11] ,
    \sb_1__1__5_chany_bottom_out[12] ,
    \sb_1__1__5_chany_bottom_out[13] ,
    \sb_1__1__5_chany_bottom_out[14] ,
    \sb_1__1__5_chany_bottom_out[15] ,
    \sb_1__1__5_chany_bottom_out[16] ,
    \sb_1__1__5_chany_bottom_out[17] ,
    \sb_1__1__5_chany_bottom_out[18] ,
    \sb_1__1__5_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__5_chany_top_out[0] ,
    \cby_1__1__5_chany_top_out[1] ,
    \cby_1__1__5_chany_top_out[2] ,
    \cby_1__1__5_chany_top_out[3] ,
    \cby_1__1__5_chany_top_out[4] ,
    \cby_1__1__5_chany_top_out[5] ,
    \cby_1__1__5_chany_top_out[6] ,
    \cby_1__1__5_chany_top_out[7] ,
    \cby_1__1__5_chany_top_out[8] ,
    \cby_1__1__5_chany_top_out[9] ,
    \cby_1__1__5_chany_top_out[10] ,
    \cby_1__1__5_chany_top_out[11] ,
    \cby_1__1__5_chany_top_out[12] ,
    \cby_1__1__5_chany_top_out[13] ,
    \cby_1__1__5_chany_top_out[14] ,
    \cby_1__1__5_chany_top_out[15] ,
    \cby_1__1__5_chany_top_out[16] ,
    \cby_1__1__5_chany_top_out[17] ,
    \cby_1__1__5_chany_top_out[18] ,
    \cby_1__1__5_chany_top_out[19] }));
 cby_1__1_ cby_1__7_ (.Test_en_E_in(\Test_enWires[102] ),
    .Test_en_S_in(\Test_enWires[102] ),
    .Test_en_W_in(\Test_enWires[102] ),
    .Test_en_W_out(\Test_enWires[100] ),
    .ccff_head(grid_clb_6_ccff_tail),
    .ccff_tail(cby_1__1__6_ccff_tail),
    .clk_2_N_out(\clk_2_wires[19] ),
    .clk_2_S_in(\clk_2_wires[18] ),
    .left_grid_pin_16_(cby_1__1__6_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__6_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__6_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__6_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__6_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__6_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__6_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__6_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__6_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__6_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__6_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__6_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__6_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__6_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__6_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__6_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[33] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[32] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[19] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[18] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__5_chany_top_out[0] ,
    \sb_1__1__5_chany_top_out[1] ,
    \sb_1__1__5_chany_top_out[2] ,
    \sb_1__1__5_chany_top_out[3] ,
    \sb_1__1__5_chany_top_out[4] ,
    \sb_1__1__5_chany_top_out[5] ,
    \sb_1__1__5_chany_top_out[6] ,
    \sb_1__1__5_chany_top_out[7] ,
    \sb_1__1__5_chany_top_out[8] ,
    \sb_1__1__5_chany_top_out[9] ,
    \sb_1__1__5_chany_top_out[10] ,
    \sb_1__1__5_chany_top_out[11] ,
    \sb_1__1__5_chany_top_out[12] ,
    \sb_1__1__5_chany_top_out[13] ,
    \sb_1__1__5_chany_top_out[14] ,
    \sb_1__1__5_chany_top_out[15] ,
    \sb_1__1__5_chany_top_out[16] ,
    \sb_1__1__5_chany_top_out[17] ,
    \sb_1__1__5_chany_top_out[18] ,
    \sb_1__1__5_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__6_chany_bottom_out[0] ,
    \cby_1__1__6_chany_bottom_out[1] ,
    \cby_1__1__6_chany_bottom_out[2] ,
    \cby_1__1__6_chany_bottom_out[3] ,
    \cby_1__1__6_chany_bottom_out[4] ,
    \cby_1__1__6_chany_bottom_out[5] ,
    \cby_1__1__6_chany_bottom_out[6] ,
    \cby_1__1__6_chany_bottom_out[7] ,
    \cby_1__1__6_chany_bottom_out[8] ,
    \cby_1__1__6_chany_bottom_out[9] ,
    \cby_1__1__6_chany_bottom_out[10] ,
    \cby_1__1__6_chany_bottom_out[11] ,
    \cby_1__1__6_chany_bottom_out[12] ,
    \cby_1__1__6_chany_bottom_out[13] ,
    \cby_1__1__6_chany_bottom_out[14] ,
    \cby_1__1__6_chany_bottom_out[15] ,
    \cby_1__1__6_chany_bottom_out[16] ,
    \cby_1__1__6_chany_bottom_out[17] ,
    \cby_1__1__6_chany_bottom_out[18] ,
    \cby_1__1__6_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__6_chany_bottom_out[0] ,
    \sb_1__1__6_chany_bottom_out[1] ,
    \sb_1__1__6_chany_bottom_out[2] ,
    \sb_1__1__6_chany_bottom_out[3] ,
    \sb_1__1__6_chany_bottom_out[4] ,
    \sb_1__1__6_chany_bottom_out[5] ,
    \sb_1__1__6_chany_bottom_out[6] ,
    \sb_1__1__6_chany_bottom_out[7] ,
    \sb_1__1__6_chany_bottom_out[8] ,
    \sb_1__1__6_chany_bottom_out[9] ,
    \sb_1__1__6_chany_bottom_out[10] ,
    \sb_1__1__6_chany_bottom_out[11] ,
    \sb_1__1__6_chany_bottom_out[12] ,
    \sb_1__1__6_chany_bottom_out[13] ,
    \sb_1__1__6_chany_bottom_out[14] ,
    \sb_1__1__6_chany_bottom_out[15] ,
    \sb_1__1__6_chany_bottom_out[16] ,
    \sb_1__1__6_chany_bottom_out[17] ,
    \sb_1__1__6_chany_bottom_out[18] ,
    \sb_1__1__6_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__6_chany_top_out[0] ,
    \cby_1__1__6_chany_top_out[1] ,
    \cby_1__1__6_chany_top_out[2] ,
    \cby_1__1__6_chany_top_out[3] ,
    \cby_1__1__6_chany_top_out[4] ,
    \cby_1__1__6_chany_top_out[5] ,
    \cby_1__1__6_chany_top_out[6] ,
    \cby_1__1__6_chany_top_out[7] ,
    \cby_1__1__6_chany_top_out[8] ,
    \cby_1__1__6_chany_top_out[9] ,
    \cby_1__1__6_chany_top_out[10] ,
    \cby_1__1__6_chany_top_out[11] ,
    \cby_1__1__6_chany_top_out[12] ,
    \cby_1__1__6_chany_top_out[13] ,
    \cby_1__1__6_chany_top_out[14] ,
    \cby_1__1__6_chany_top_out[15] ,
    \cby_1__1__6_chany_top_out[16] ,
    \cby_1__1__6_chany_top_out[17] ,
    \cby_1__1__6_chany_top_out[18] ,
    \cby_1__1__6_chany_top_out[19] }));
 cby_1__1_ cby_1__8_ (.Test_en_E_in(\Test_enWires[116] ),
    .Test_en_S_in(\Test_enWires[116] ),
    .Test_en_W_in(\Test_enWires[116] ),
    .Test_en_W_out(\Test_enWires[114] ),
    .ccff_head(grid_clb_7_ccff_tail),
    .ccff_tail(cby_1__1__7_ccff_tail),
    .left_grid_pin_16_(cby_1__1__7_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__7_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__7_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__7_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__7_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__7_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__7_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__7_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__7_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__7_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__7_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__7_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__7_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__7_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__7_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__7_left_grid_pin_31_),
    .prog_clk_0_N_out(\prog_clk_0_wires[40] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[38] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[37] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__6_chany_top_out[0] ,
    \sb_1__1__6_chany_top_out[1] ,
    \sb_1__1__6_chany_top_out[2] ,
    \sb_1__1__6_chany_top_out[3] ,
    \sb_1__1__6_chany_top_out[4] ,
    \sb_1__1__6_chany_top_out[5] ,
    \sb_1__1__6_chany_top_out[6] ,
    \sb_1__1__6_chany_top_out[7] ,
    \sb_1__1__6_chany_top_out[8] ,
    \sb_1__1__6_chany_top_out[9] ,
    \sb_1__1__6_chany_top_out[10] ,
    \sb_1__1__6_chany_top_out[11] ,
    \sb_1__1__6_chany_top_out[12] ,
    \sb_1__1__6_chany_top_out[13] ,
    \sb_1__1__6_chany_top_out[14] ,
    \sb_1__1__6_chany_top_out[15] ,
    \sb_1__1__6_chany_top_out[16] ,
    \sb_1__1__6_chany_top_out[17] ,
    \sb_1__1__6_chany_top_out[18] ,
    \sb_1__1__6_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__7_chany_bottom_out[0] ,
    \cby_1__1__7_chany_bottom_out[1] ,
    \cby_1__1__7_chany_bottom_out[2] ,
    \cby_1__1__7_chany_bottom_out[3] ,
    \cby_1__1__7_chany_bottom_out[4] ,
    \cby_1__1__7_chany_bottom_out[5] ,
    \cby_1__1__7_chany_bottom_out[6] ,
    \cby_1__1__7_chany_bottom_out[7] ,
    \cby_1__1__7_chany_bottom_out[8] ,
    \cby_1__1__7_chany_bottom_out[9] ,
    \cby_1__1__7_chany_bottom_out[10] ,
    \cby_1__1__7_chany_bottom_out[11] ,
    \cby_1__1__7_chany_bottom_out[12] ,
    \cby_1__1__7_chany_bottom_out[13] ,
    \cby_1__1__7_chany_bottom_out[14] ,
    \cby_1__1__7_chany_bottom_out[15] ,
    \cby_1__1__7_chany_bottom_out[16] ,
    \cby_1__1__7_chany_bottom_out[17] ,
    \cby_1__1__7_chany_bottom_out[18] ,
    \cby_1__1__7_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__8__0_chany_bottom_out[0] ,
    \sb_1__8__0_chany_bottom_out[1] ,
    \sb_1__8__0_chany_bottom_out[2] ,
    \sb_1__8__0_chany_bottom_out[3] ,
    \sb_1__8__0_chany_bottom_out[4] ,
    \sb_1__8__0_chany_bottom_out[5] ,
    \sb_1__8__0_chany_bottom_out[6] ,
    \sb_1__8__0_chany_bottom_out[7] ,
    \sb_1__8__0_chany_bottom_out[8] ,
    \sb_1__8__0_chany_bottom_out[9] ,
    \sb_1__8__0_chany_bottom_out[10] ,
    \sb_1__8__0_chany_bottom_out[11] ,
    \sb_1__8__0_chany_bottom_out[12] ,
    \sb_1__8__0_chany_bottom_out[13] ,
    \sb_1__8__0_chany_bottom_out[14] ,
    \sb_1__8__0_chany_bottom_out[15] ,
    \sb_1__8__0_chany_bottom_out[16] ,
    \sb_1__8__0_chany_bottom_out[17] ,
    \sb_1__8__0_chany_bottom_out[18] ,
    \sb_1__8__0_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__7_chany_top_out[0] ,
    \cby_1__1__7_chany_top_out[1] ,
    \cby_1__1__7_chany_top_out[2] ,
    \cby_1__1__7_chany_top_out[3] ,
    \cby_1__1__7_chany_top_out[4] ,
    \cby_1__1__7_chany_top_out[5] ,
    \cby_1__1__7_chany_top_out[6] ,
    \cby_1__1__7_chany_top_out[7] ,
    \cby_1__1__7_chany_top_out[8] ,
    \cby_1__1__7_chany_top_out[9] ,
    \cby_1__1__7_chany_top_out[10] ,
    \cby_1__1__7_chany_top_out[11] ,
    \cby_1__1__7_chany_top_out[12] ,
    \cby_1__1__7_chany_top_out[13] ,
    \cby_1__1__7_chany_top_out[14] ,
    \cby_1__1__7_chany_top_out[15] ,
    \cby_1__1__7_chany_top_out[16] ,
    \cby_1__1__7_chany_top_out[17] ,
    \cby_1__1__7_chany_top_out[18] ,
    \cby_1__1__7_chany_top_out[19] }));
 cby_1__1_ cby_2__1_ (.Test_en_E_in(\Test_enWires[20] ),
    .Test_en_S_in(\Test_enWires[20] ),
    .Test_en_W_in(\Test_enWires[20] ),
    .Test_en_W_out(\Test_enWires[17] ),
    .ccff_head(grid_clb_8_ccff_tail),
    .ccff_tail(cby_1__1__8_ccff_tail),
    .left_grid_pin_16_(cby_1__1__8_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__8_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__8_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__8_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__8_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__8_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__8_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__8_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__8_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__8_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__8_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__8_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__8_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__8_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__8_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__8_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[45] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[44] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__0__1_chany_top_out[0] ,
    \sb_1__0__1_chany_top_out[1] ,
    \sb_1__0__1_chany_top_out[2] ,
    \sb_1__0__1_chany_top_out[3] ,
    \sb_1__0__1_chany_top_out[4] ,
    \sb_1__0__1_chany_top_out[5] ,
    \sb_1__0__1_chany_top_out[6] ,
    \sb_1__0__1_chany_top_out[7] ,
    \sb_1__0__1_chany_top_out[8] ,
    \sb_1__0__1_chany_top_out[9] ,
    \sb_1__0__1_chany_top_out[10] ,
    \sb_1__0__1_chany_top_out[11] ,
    \sb_1__0__1_chany_top_out[12] ,
    \sb_1__0__1_chany_top_out[13] ,
    \sb_1__0__1_chany_top_out[14] ,
    \sb_1__0__1_chany_top_out[15] ,
    \sb_1__0__1_chany_top_out[16] ,
    \sb_1__0__1_chany_top_out[17] ,
    \sb_1__0__1_chany_top_out[18] ,
    \sb_1__0__1_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__8_chany_bottom_out[0] ,
    \cby_1__1__8_chany_bottom_out[1] ,
    \cby_1__1__8_chany_bottom_out[2] ,
    \cby_1__1__8_chany_bottom_out[3] ,
    \cby_1__1__8_chany_bottom_out[4] ,
    \cby_1__1__8_chany_bottom_out[5] ,
    \cby_1__1__8_chany_bottom_out[6] ,
    \cby_1__1__8_chany_bottom_out[7] ,
    \cby_1__1__8_chany_bottom_out[8] ,
    \cby_1__1__8_chany_bottom_out[9] ,
    \cby_1__1__8_chany_bottom_out[10] ,
    \cby_1__1__8_chany_bottom_out[11] ,
    \cby_1__1__8_chany_bottom_out[12] ,
    \cby_1__1__8_chany_bottom_out[13] ,
    \cby_1__1__8_chany_bottom_out[14] ,
    \cby_1__1__8_chany_bottom_out[15] ,
    \cby_1__1__8_chany_bottom_out[16] ,
    \cby_1__1__8_chany_bottom_out[17] ,
    \cby_1__1__8_chany_bottom_out[18] ,
    \cby_1__1__8_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__7_chany_bottom_out[0] ,
    \sb_1__1__7_chany_bottom_out[1] ,
    \sb_1__1__7_chany_bottom_out[2] ,
    \sb_1__1__7_chany_bottom_out[3] ,
    \sb_1__1__7_chany_bottom_out[4] ,
    \sb_1__1__7_chany_bottom_out[5] ,
    \sb_1__1__7_chany_bottom_out[6] ,
    \sb_1__1__7_chany_bottom_out[7] ,
    \sb_1__1__7_chany_bottom_out[8] ,
    \sb_1__1__7_chany_bottom_out[9] ,
    \sb_1__1__7_chany_bottom_out[10] ,
    \sb_1__1__7_chany_bottom_out[11] ,
    \sb_1__1__7_chany_bottom_out[12] ,
    \sb_1__1__7_chany_bottom_out[13] ,
    \sb_1__1__7_chany_bottom_out[14] ,
    \sb_1__1__7_chany_bottom_out[15] ,
    \sb_1__1__7_chany_bottom_out[16] ,
    \sb_1__1__7_chany_bottom_out[17] ,
    \sb_1__1__7_chany_bottom_out[18] ,
    \sb_1__1__7_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__8_chany_top_out[0] ,
    \cby_1__1__8_chany_top_out[1] ,
    \cby_1__1__8_chany_top_out[2] ,
    \cby_1__1__8_chany_top_out[3] ,
    \cby_1__1__8_chany_top_out[4] ,
    \cby_1__1__8_chany_top_out[5] ,
    \cby_1__1__8_chany_top_out[6] ,
    \cby_1__1__8_chany_top_out[7] ,
    \cby_1__1__8_chany_top_out[8] ,
    \cby_1__1__8_chany_top_out[9] ,
    \cby_1__1__8_chany_top_out[10] ,
    \cby_1__1__8_chany_top_out[11] ,
    \cby_1__1__8_chany_top_out[12] ,
    \cby_1__1__8_chany_top_out[13] ,
    \cby_1__1__8_chany_top_out[14] ,
    \cby_1__1__8_chany_top_out[15] ,
    \cby_1__1__8_chany_top_out[16] ,
    \cby_1__1__8_chany_top_out[17] ,
    \cby_1__1__8_chany_top_out[18] ,
    \cby_1__1__8_chany_top_out[19] }));
 cby_1__1_ cby_2__2_ (.Test_en_E_in(\Test_enWires[34] ),
    .Test_en_S_in(\Test_enWires[34] ),
    .Test_en_W_in(\Test_enWires[34] ),
    .Test_en_W_out(\Test_enWires[31] ),
    .ccff_head(grid_clb_9_ccff_tail),
    .ccff_tail(cby_1__1__9_ccff_tail),
    .left_grid_pin_16_(cby_1__1__9_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__9_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__9_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__9_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__9_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__9_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__9_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__9_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__9_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__9_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__9_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__9_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__9_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__9_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__9_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__9_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[48] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[47] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__7_chany_top_out[0] ,
    \sb_1__1__7_chany_top_out[1] ,
    \sb_1__1__7_chany_top_out[2] ,
    \sb_1__1__7_chany_top_out[3] ,
    \sb_1__1__7_chany_top_out[4] ,
    \sb_1__1__7_chany_top_out[5] ,
    \sb_1__1__7_chany_top_out[6] ,
    \sb_1__1__7_chany_top_out[7] ,
    \sb_1__1__7_chany_top_out[8] ,
    \sb_1__1__7_chany_top_out[9] ,
    \sb_1__1__7_chany_top_out[10] ,
    \sb_1__1__7_chany_top_out[11] ,
    \sb_1__1__7_chany_top_out[12] ,
    \sb_1__1__7_chany_top_out[13] ,
    \sb_1__1__7_chany_top_out[14] ,
    \sb_1__1__7_chany_top_out[15] ,
    \sb_1__1__7_chany_top_out[16] ,
    \sb_1__1__7_chany_top_out[17] ,
    \sb_1__1__7_chany_top_out[18] ,
    \sb_1__1__7_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__9_chany_bottom_out[0] ,
    \cby_1__1__9_chany_bottom_out[1] ,
    \cby_1__1__9_chany_bottom_out[2] ,
    \cby_1__1__9_chany_bottom_out[3] ,
    \cby_1__1__9_chany_bottom_out[4] ,
    \cby_1__1__9_chany_bottom_out[5] ,
    \cby_1__1__9_chany_bottom_out[6] ,
    \cby_1__1__9_chany_bottom_out[7] ,
    \cby_1__1__9_chany_bottom_out[8] ,
    \cby_1__1__9_chany_bottom_out[9] ,
    \cby_1__1__9_chany_bottom_out[10] ,
    \cby_1__1__9_chany_bottom_out[11] ,
    \cby_1__1__9_chany_bottom_out[12] ,
    \cby_1__1__9_chany_bottom_out[13] ,
    \cby_1__1__9_chany_bottom_out[14] ,
    \cby_1__1__9_chany_bottom_out[15] ,
    \cby_1__1__9_chany_bottom_out[16] ,
    \cby_1__1__9_chany_bottom_out[17] ,
    \cby_1__1__9_chany_bottom_out[18] ,
    \cby_1__1__9_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__8_chany_bottom_out[0] ,
    \sb_1__1__8_chany_bottom_out[1] ,
    \sb_1__1__8_chany_bottom_out[2] ,
    \sb_1__1__8_chany_bottom_out[3] ,
    \sb_1__1__8_chany_bottom_out[4] ,
    \sb_1__1__8_chany_bottom_out[5] ,
    \sb_1__1__8_chany_bottom_out[6] ,
    \sb_1__1__8_chany_bottom_out[7] ,
    \sb_1__1__8_chany_bottom_out[8] ,
    \sb_1__1__8_chany_bottom_out[9] ,
    \sb_1__1__8_chany_bottom_out[10] ,
    \sb_1__1__8_chany_bottom_out[11] ,
    \sb_1__1__8_chany_bottom_out[12] ,
    \sb_1__1__8_chany_bottom_out[13] ,
    \sb_1__1__8_chany_bottom_out[14] ,
    \sb_1__1__8_chany_bottom_out[15] ,
    \sb_1__1__8_chany_bottom_out[16] ,
    \sb_1__1__8_chany_bottom_out[17] ,
    \sb_1__1__8_chany_bottom_out[18] ,
    \sb_1__1__8_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__9_chany_top_out[0] ,
    \cby_1__1__9_chany_top_out[1] ,
    \cby_1__1__9_chany_top_out[2] ,
    \cby_1__1__9_chany_top_out[3] ,
    \cby_1__1__9_chany_top_out[4] ,
    \cby_1__1__9_chany_top_out[5] ,
    \cby_1__1__9_chany_top_out[6] ,
    \cby_1__1__9_chany_top_out[7] ,
    \cby_1__1__9_chany_top_out[8] ,
    \cby_1__1__9_chany_top_out[9] ,
    \cby_1__1__9_chany_top_out[10] ,
    \cby_1__1__9_chany_top_out[11] ,
    \cby_1__1__9_chany_top_out[12] ,
    \cby_1__1__9_chany_top_out[13] ,
    \cby_1__1__9_chany_top_out[14] ,
    \cby_1__1__9_chany_top_out[15] ,
    \cby_1__1__9_chany_top_out[16] ,
    \cby_1__1__9_chany_top_out[17] ,
    \cby_1__1__9_chany_top_out[18] ,
    \cby_1__1__9_chany_top_out[19] }));
 cby_1__1_ cby_2__3_ (.Test_en_E_in(\Test_enWires[48] ),
    .Test_en_S_in(\Test_enWires[48] ),
    .Test_en_W_in(\Test_enWires[48] ),
    .Test_en_W_out(\Test_enWires[45] ),
    .ccff_head(grid_clb_10_ccff_tail),
    .ccff_tail(cby_1__1__10_ccff_tail),
    .clk_3_S_in(\clk_3_wires[16] ),
    .clk_3_S_out(\clk_3_wires[17] ),
    .left_grid_pin_16_(cby_1__1__10_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__10_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__10_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__10_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__10_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__10_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__10_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__10_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__10_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__10_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__10_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__10_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__10_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__10_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__10_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__10_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[51] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[50] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[16] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[17] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__8_chany_top_out[0] ,
    \sb_1__1__8_chany_top_out[1] ,
    \sb_1__1__8_chany_top_out[2] ,
    \sb_1__1__8_chany_top_out[3] ,
    \sb_1__1__8_chany_top_out[4] ,
    \sb_1__1__8_chany_top_out[5] ,
    \sb_1__1__8_chany_top_out[6] ,
    \sb_1__1__8_chany_top_out[7] ,
    \sb_1__1__8_chany_top_out[8] ,
    \sb_1__1__8_chany_top_out[9] ,
    \sb_1__1__8_chany_top_out[10] ,
    \sb_1__1__8_chany_top_out[11] ,
    \sb_1__1__8_chany_top_out[12] ,
    \sb_1__1__8_chany_top_out[13] ,
    \sb_1__1__8_chany_top_out[14] ,
    \sb_1__1__8_chany_top_out[15] ,
    \sb_1__1__8_chany_top_out[16] ,
    \sb_1__1__8_chany_top_out[17] ,
    \sb_1__1__8_chany_top_out[18] ,
    \sb_1__1__8_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__10_chany_bottom_out[0] ,
    \cby_1__1__10_chany_bottom_out[1] ,
    \cby_1__1__10_chany_bottom_out[2] ,
    \cby_1__1__10_chany_bottom_out[3] ,
    \cby_1__1__10_chany_bottom_out[4] ,
    \cby_1__1__10_chany_bottom_out[5] ,
    \cby_1__1__10_chany_bottom_out[6] ,
    \cby_1__1__10_chany_bottom_out[7] ,
    \cby_1__1__10_chany_bottom_out[8] ,
    \cby_1__1__10_chany_bottom_out[9] ,
    \cby_1__1__10_chany_bottom_out[10] ,
    \cby_1__1__10_chany_bottom_out[11] ,
    \cby_1__1__10_chany_bottom_out[12] ,
    \cby_1__1__10_chany_bottom_out[13] ,
    \cby_1__1__10_chany_bottom_out[14] ,
    \cby_1__1__10_chany_bottom_out[15] ,
    \cby_1__1__10_chany_bottom_out[16] ,
    \cby_1__1__10_chany_bottom_out[17] ,
    \cby_1__1__10_chany_bottom_out[18] ,
    \cby_1__1__10_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__9_chany_bottom_out[0] ,
    \sb_1__1__9_chany_bottom_out[1] ,
    \sb_1__1__9_chany_bottom_out[2] ,
    \sb_1__1__9_chany_bottom_out[3] ,
    \sb_1__1__9_chany_bottom_out[4] ,
    \sb_1__1__9_chany_bottom_out[5] ,
    \sb_1__1__9_chany_bottom_out[6] ,
    \sb_1__1__9_chany_bottom_out[7] ,
    \sb_1__1__9_chany_bottom_out[8] ,
    \sb_1__1__9_chany_bottom_out[9] ,
    \sb_1__1__9_chany_bottom_out[10] ,
    \sb_1__1__9_chany_bottom_out[11] ,
    \sb_1__1__9_chany_bottom_out[12] ,
    \sb_1__1__9_chany_bottom_out[13] ,
    \sb_1__1__9_chany_bottom_out[14] ,
    \sb_1__1__9_chany_bottom_out[15] ,
    \sb_1__1__9_chany_bottom_out[16] ,
    \sb_1__1__9_chany_bottom_out[17] ,
    \sb_1__1__9_chany_bottom_out[18] ,
    \sb_1__1__9_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__10_chany_top_out[0] ,
    \cby_1__1__10_chany_top_out[1] ,
    \cby_1__1__10_chany_top_out[2] ,
    \cby_1__1__10_chany_top_out[3] ,
    \cby_1__1__10_chany_top_out[4] ,
    \cby_1__1__10_chany_top_out[5] ,
    \cby_1__1__10_chany_top_out[6] ,
    \cby_1__1__10_chany_top_out[7] ,
    \cby_1__1__10_chany_top_out[8] ,
    \cby_1__1__10_chany_top_out[9] ,
    \cby_1__1__10_chany_top_out[10] ,
    \cby_1__1__10_chany_top_out[11] ,
    \cby_1__1__10_chany_top_out[12] ,
    \cby_1__1__10_chany_top_out[13] ,
    \cby_1__1__10_chany_top_out[14] ,
    \cby_1__1__10_chany_top_out[15] ,
    \cby_1__1__10_chany_top_out[16] ,
    \cby_1__1__10_chany_top_out[17] ,
    \cby_1__1__10_chany_top_out[18] ,
    \cby_1__1__10_chany_top_out[19] }));
 cby_1__1_ cby_2__4_ (.Test_en_E_in(\Test_enWires[62] ),
    .Test_en_S_in(\Test_enWires[62] ),
    .Test_en_W_in(\Test_enWires[62] ),
    .Test_en_W_out(\Test_enWires[59] ),
    .ccff_head(grid_clb_11_ccff_tail),
    .ccff_tail(cby_1__1__11_ccff_tail),
    .clk_3_S_in(\clk_3_wires[12] ),
    .clk_3_S_out(\clk_3_wires[13] ),
    .left_grid_pin_16_(cby_1__1__11_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__11_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__11_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__11_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__11_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__11_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__11_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__11_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__11_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__11_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__11_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__11_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__11_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__11_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__11_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__11_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[54] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[53] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[12] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[13] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__9_chany_top_out[0] ,
    \sb_1__1__9_chany_top_out[1] ,
    \sb_1__1__9_chany_top_out[2] ,
    \sb_1__1__9_chany_top_out[3] ,
    \sb_1__1__9_chany_top_out[4] ,
    \sb_1__1__9_chany_top_out[5] ,
    \sb_1__1__9_chany_top_out[6] ,
    \sb_1__1__9_chany_top_out[7] ,
    \sb_1__1__9_chany_top_out[8] ,
    \sb_1__1__9_chany_top_out[9] ,
    \sb_1__1__9_chany_top_out[10] ,
    \sb_1__1__9_chany_top_out[11] ,
    \sb_1__1__9_chany_top_out[12] ,
    \sb_1__1__9_chany_top_out[13] ,
    \sb_1__1__9_chany_top_out[14] ,
    \sb_1__1__9_chany_top_out[15] ,
    \sb_1__1__9_chany_top_out[16] ,
    \sb_1__1__9_chany_top_out[17] ,
    \sb_1__1__9_chany_top_out[18] ,
    \sb_1__1__9_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__11_chany_bottom_out[0] ,
    \cby_1__1__11_chany_bottom_out[1] ,
    \cby_1__1__11_chany_bottom_out[2] ,
    \cby_1__1__11_chany_bottom_out[3] ,
    \cby_1__1__11_chany_bottom_out[4] ,
    \cby_1__1__11_chany_bottom_out[5] ,
    \cby_1__1__11_chany_bottom_out[6] ,
    \cby_1__1__11_chany_bottom_out[7] ,
    \cby_1__1__11_chany_bottom_out[8] ,
    \cby_1__1__11_chany_bottom_out[9] ,
    \cby_1__1__11_chany_bottom_out[10] ,
    \cby_1__1__11_chany_bottom_out[11] ,
    \cby_1__1__11_chany_bottom_out[12] ,
    \cby_1__1__11_chany_bottom_out[13] ,
    \cby_1__1__11_chany_bottom_out[14] ,
    \cby_1__1__11_chany_bottom_out[15] ,
    \cby_1__1__11_chany_bottom_out[16] ,
    \cby_1__1__11_chany_bottom_out[17] ,
    \cby_1__1__11_chany_bottom_out[18] ,
    \cby_1__1__11_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__10_chany_bottom_out[0] ,
    \sb_1__1__10_chany_bottom_out[1] ,
    \sb_1__1__10_chany_bottom_out[2] ,
    \sb_1__1__10_chany_bottom_out[3] ,
    \sb_1__1__10_chany_bottom_out[4] ,
    \sb_1__1__10_chany_bottom_out[5] ,
    \sb_1__1__10_chany_bottom_out[6] ,
    \sb_1__1__10_chany_bottom_out[7] ,
    \sb_1__1__10_chany_bottom_out[8] ,
    \sb_1__1__10_chany_bottom_out[9] ,
    \sb_1__1__10_chany_bottom_out[10] ,
    \sb_1__1__10_chany_bottom_out[11] ,
    \sb_1__1__10_chany_bottom_out[12] ,
    \sb_1__1__10_chany_bottom_out[13] ,
    \sb_1__1__10_chany_bottom_out[14] ,
    \sb_1__1__10_chany_bottom_out[15] ,
    \sb_1__1__10_chany_bottom_out[16] ,
    \sb_1__1__10_chany_bottom_out[17] ,
    \sb_1__1__10_chany_bottom_out[18] ,
    \sb_1__1__10_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__11_chany_top_out[0] ,
    \cby_1__1__11_chany_top_out[1] ,
    \cby_1__1__11_chany_top_out[2] ,
    \cby_1__1__11_chany_top_out[3] ,
    \cby_1__1__11_chany_top_out[4] ,
    \cby_1__1__11_chany_top_out[5] ,
    \cby_1__1__11_chany_top_out[6] ,
    \cby_1__1__11_chany_top_out[7] ,
    \cby_1__1__11_chany_top_out[8] ,
    \cby_1__1__11_chany_top_out[9] ,
    \cby_1__1__11_chany_top_out[10] ,
    \cby_1__1__11_chany_top_out[11] ,
    \cby_1__1__11_chany_top_out[12] ,
    \cby_1__1__11_chany_top_out[13] ,
    \cby_1__1__11_chany_top_out[14] ,
    \cby_1__1__11_chany_top_out[15] ,
    \cby_1__1__11_chany_top_out[16] ,
    \cby_1__1__11_chany_top_out[17] ,
    \cby_1__1__11_chany_top_out[18] ,
    \cby_1__1__11_chany_top_out[19] }));
 cby_1__1_ cby_2__5_ (.Test_en_E_in(\Test_enWires[76] ),
    .Test_en_S_in(\Test_enWires[76] ),
    .Test_en_W_in(\Test_enWires[76] ),
    .Test_en_W_out(\Test_enWires[73] ),
    .ccff_head(grid_clb_12_ccff_tail),
    .ccff_tail(cby_1__1__12_ccff_tail),
    .clk_3_N_out(\clk_3_wires[11] ),
    .clk_3_S_in(\clk_3_wires[10] ),
    .left_grid_pin_16_(cby_1__1__12_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__12_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__12_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__12_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__12_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__12_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__12_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__12_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__12_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__12_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__12_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__12_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__12_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__12_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__12_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__12_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[57] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[56] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[11] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[10] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__10_chany_top_out[0] ,
    \sb_1__1__10_chany_top_out[1] ,
    \sb_1__1__10_chany_top_out[2] ,
    \sb_1__1__10_chany_top_out[3] ,
    \sb_1__1__10_chany_top_out[4] ,
    \sb_1__1__10_chany_top_out[5] ,
    \sb_1__1__10_chany_top_out[6] ,
    \sb_1__1__10_chany_top_out[7] ,
    \sb_1__1__10_chany_top_out[8] ,
    \sb_1__1__10_chany_top_out[9] ,
    \sb_1__1__10_chany_top_out[10] ,
    \sb_1__1__10_chany_top_out[11] ,
    \sb_1__1__10_chany_top_out[12] ,
    \sb_1__1__10_chany_top_out[13] ,
    \sb_1__1__10_chany_top_out[14] ,
    \sb_1__1__10_chany_top_out[15] ,
    \sb_1__1__10_chany_top_out[16] ,
    \sb_1__1__10_chany_top_out[17] ,
    \sb_1__1__10_chany_top_out[18] ,
    \sb_1__1__10_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__12_chany_bottom_out[0] ,
    \cby_1__1__12_chany_bottom_out[1] ,
    \cby_1__1__12_chany_bottom_out[2] ,
    \cby_1__1__12_chany_bottom_out[3] ,
    \cby_1__1__12_chany_bottom_out[4] ,
    \cby_1__1__12_chany_bottom_out[5] ,
    \cby_1__1__12_chany_bottom_out[6] ,
    \cby_1__1__12_chany_bottom_out[7] ,
    \cby_1__1__12_chany_bottom_out[8] ,
    \cby_1__1__12_chany_bottom_out[9] ,
    \cby_1__1__12_chany_bottom_out[10] ,
    \cby_1__1__12_chany_bottom_out[11] ,
    \cby_1__1__12_chany_bottom_out[12] ,
    \cby_1__1__12_chany_bottom_out[13] ,
    \cby_1__1__12_chany_bottom_out[14] ,
    \cby_1__1__12_chany_bottom_out[15] ,
    \cby_1__1__12_chany_bottom_out[16] ,
    \cby_1__1__12_chany_bottom_out[17] ,
    \cby_1__1__12_chany_bottom_out[18] ,
    \cby_1__1__12_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__11_chany_bottom_out[0] ,
    \sb_1__1__11_chany_bottom_out[1] ,
    \sb_1__1__11_chany_bottom_out[2] ,
    \sb_1__1__11_chany_bottom_out[3] ,
    \sb_1__1__11_chany_bottom_out[4] ,
    \sb_1__1__11_chany_bottom_out[5] ,
    \sb_1__1__11_chany_bottom_out[6] ,
    \sb_1__1__11_chany_bottom_out[7] ,
    \sb_1__1__11_chany_bottom_out[8] ,
    \sb_1__1__11_chany_bottom_out[9] ,
    \sb_1__1__11_chany_bottom_out[10] ,
    \sb_1__1__11_chany_bottom_out[11] ,
    \sb_1__1__11_chany_bottom_out[12] ,
    \sb_1__1__11_chany_bottom_out[13] ,
    \sb_1__1__11_chany_bottom_out[14] ,
    \sb_1__1__11_chany_bottom_out[15] ,
    \sb_1__1__11_chany_bottom_out[16] ,
    \sb_1__1__11_chany_bottom_out[17] ,
    \sb_1__1__11_chany_bottom_out[18] ,
    \sb_1__1__11_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__12_chany_top_out[0] ,
    \cby_1__1__12_chany_top_out[1] ,
    \cby_1__1__12_chany_top_out[2] ,
    \cby_1__1__12_chany_top_out[3] ,
    \cby_1__1__12_chany_top_out[4] ,
    \cby_1__1__12_chany_top_out[5] ,
    \cby_1__1__12_chany_top_out[6] ,
    \cby_1__1__12_chany_top_out[7] ,
    \cby_1__1__12_chany_top_out[8] ,
    \cby_1__1__12_chany_top_out[9] ,
    \cby_1__1__12_chany_top_out[10] ,
    \cby_1__1__12_chany_top_out[11] ,
    \cby_1__1__12_chany_top_out[12] ,
    \cby_1__1__12_chany_top_out[13] ,
    \cby_1__1__12_chany_top_out[14] ,
    \cby_1__1__12_chany_top_out[15] ,
    \cby_1__1__12_chany_top_out[16] ,
    \cby_1__1__12_chany_top_out[17] ,
    \cby_1__1__12_chany_top_out[18] ,
    \cby_1__1__12_chany_top_out[19] }));
 cby_1__1_ cby_2__6_ (.Test_en_E_in(\Test_enWires[90] ),
    .Test_en_S_in(\Test_enWires[90] ),
    .Test_en_W_in(\Test_enWires[90] ),
    .Test_en_W_out(\Test_enWires[87] ),
    .ccff_head(grid_clb_13_ccff_tail),
    .ccff_tail(cby_1__1__13_ccff_tail),
    .clk_3_N_out(\clk_3_wires[15] ),
    .clk_3_S_in(\clk_3_wires[14] ),
    .left_grid_pin_16_(cby_1__1__13_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__13_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__13_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__13_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__13_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__13_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__13_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__13_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__13_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__13_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__13_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__13_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__13_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__13_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__13_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__13_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[60] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[59] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[15] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[14] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__11_chany_top_out[0] ,
    \sb_1__1__11_chany_top_out[1] ,
    \sb_1__1__11_chany_top_out[2] ,
    \sb_1__1__11_chany_top_out[3] ,
    \sb_1__1__11_chany_top_out[4] ,
    \sb_1__1__11_chany_top_out[5] ,
    \sb_1__1__11_chany_top_out[6] ,
    \sb_1__1__11_chany_top_out[7] ,
    \sb_1__1__11_chany_top_out[8] ,
    \sb_1__1__11_chany_top_out[9] ,
    \sb_1__1__11_chany_top_out[10] ,
    \sb_1__1__11_chany_top_out[11] ,
    \sb_1__1__11_chany_top_out[12] ,
    \sb_1__1__11_chany_top_out[13] ,
    \sb_1__1__11_chany_top_out[14] ,
    \sb_1__1__11_chany_top_out[15] ,
    \sb_1__1__11_chany_top_out[16] ,
    \sb_1__1__11_chany_top_out[17] ,
    \sb_1__1__11_chany_top_out[18] ,
    \sb_1__1__11_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__13_chany_bottom_out[0] ,
    \cby_1__1__13_chany_bottom_out[1] ,
    \cby_1__1__13_chany_bottom_out[2] ,
    \cby_1__1__13_chany_bottom_out[3] ,
    \cby_1__1__13_chany_bottom_out[4] ,
    \cby_1__1__13_chany_bottom_out[5] ,
    \cby_1__1__13_chany_bottom_out[6] ,
    \cby_1__1__13_chany_bottom_out[7] ,
    \cby_1__1__13_chany_bottom_out[8] ,
    \cby_1__1__13_chany_bottom_out[9] ,
    \cby_1__1__13_chany_bottom_out[10] ,
    \cby_1__1__13_chany_bottom_out[11] ,
    \cby_1__1__13_chany_bottom_out[12] ,
    \cby_1__1__13_chany_bottom_out[13] ,
    \cby_1__1__13_chany_bottom_out[14] ,
    \cby_1__1__13_chany_bottom_out[15] ,
    \cby_1__1__13_chany_bottom_out[16] ,
    \cby_1__1__13_chany_bottom_out[17] ,
    \cby_1__1__13_chany_bottom_out[18] ,
    \cby_1__1__13_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__12_chany_bottom_out[0] ,
    \sb_1__1__12_chany_bottom_out[1] ,
    \sb_1__1__12_chany_bottom_out[2] ,
    \sb_1__1__12_chany_bottom_out[3] ,
    \sb_1__1__12_chany_bottom_out[4] ,
    \sb_1__1__12_chany_bottom_out[5] ,
    \sb_1__1__12_chany_bottom_out[6] ,
    \sb_1__1__12_chany_bottom_out[7] ,
    \sb_1__1__12_chany_bottom_out[8] ,
    \sb_1__1__12_chany_bottom_out[9] ,
    \sb_1__1__12_chany_bottom_out[10] ,
    \sb_1__1__12_chany_bottom_out[11] ,
    \sb_1__1__12_chany_bottom_out[12] ,
    \sb_1__1__12_chany_bottom_out[13] ,
    \sb_1__1__12_chany_bottom_out[14] ,
    \sb_1__1__12_chany_bottom_out[15] ,
    \sb_1__1__12_chany_bottom_out[16] ,
    \sb_1__1__12_chany_bottom_out[17] ,
    \sb_1__1__12_chany_bottom_out[18] ,
    \sb_1__1__12_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__13_chany_top_out[0] ,
    \cby_1__1__13_chany_top_out[1] ,
    \cby_1__1__13_chany_top_out[2] ,
    \cby_1__1__13_chany_top_out[3] ,
    \cby_1__1__13_chany_top_out[4] ,
    \cby_1__1__13_chany_top_out[5] ,
    \cby_1__1__13_chany_top_out[6] ,
    \cby_1__1__13_chany_top_out[7] ,
    \cby_1__1__13_chany_top_out[8] ,
    \cby_1__1__13_chany_top_out[9] ,
    \cby_1__1__13_chany_top_out[10] ,
    \cby_1__1__13_chany_top_out[11] ,
    \cby_1__1__13_chany_top_out[12] ,
    \cby_1__1__13_chany_top_out[13] ,
    \cby_1__1__13_chany_top_out[14] ,
    \cby_1__1__13_chany_top_out[15] ,
    \cby_1__1__13_chany_top_out[16] ,
    \cby_1__1__13_chany_top_out[17] ,
    \cby_1__1__13_chany_top_out[18] ,
    \cby_1__1__13_chany_top_out[19] }));
 cby_1__1_ cby_2__7_ (.Test_en_E_in(\Test_enWires[104] ),
    .Test_en_S_in(\Test_enWires[104] ),
    .Test_en_W_in(\Test_enWires[104] ),
    .Test_en_W_out(\Test_enWires[101] ),
    .ccff_head(grid_clb_14_ccff_tail),
    .ccff_tail(cby_1__1__14_ccff_tail),
    .left_grid_pin_16_(cby_1__1__14_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__14_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__14_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__14_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__14_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__14_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__14_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__14_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__14_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__14_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__14_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__14_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__14_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__14_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__14_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__14_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[63] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[62] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__12_chany_top_out[0] ,
    \sb_1__1__12_chany_top_out[1] ,
    \sb_1__1__12_chany_top_out[2] ,
    \sb_1__1__12_chany_top_out[3] ,
    \sb_1__1__12_chany_top_out[4] ,
    \sb_1__1__12_chany_top_out[5] ,
    \sb_1__1__12_chany_top_out[6] ,
    \sb_1__1__12_chany_top_out[7] ,
    \sb_1__1__12_chany_top_out[8] ,
    \sb_1__1__12_chany_top_out[9] ,
    \sb_1__1__12_chany_top_out[10] ,
    \sb_1__1__12_chany_top_out[11] ,
    \sb_1__1__12_chany_top_out[12] ,
    \sb_1__1__12_chany_top_out[13] ,
    \sb_1__1__12_chany_top_out[14] ,
    \sb_1__1__12_chany_top_out[15] ,
    \sb_1__1__12_chany_top_out[16] ,
    \sb_1__1__12_chany_top_out[17] ,
    \sb_1__1__12_chany_top_out[18] ,
    \sb_1__1__12_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__14_chany_bottom_out[0] ,
    \cby_1__1__14_chany_bottom_out[1] ,
    \cby_1__1__14_chany_bottom_out[2] ,
    \cby_1__1__14_chany_bottom_out[3] ,
    \cby_1__1__14_chany_bottom_out[4] ,
    \cby_1__1__14_chany_bottom_out[5] ,
    \cby_1__1__14_chany_bottom_out[6] ,
    \cby_1__1__14_chany_bottom_out[7] ,
    \cby_1__1__14_chany_bottom_out[8] ,
    \cby_1__1__14_chany_bottom_out[9] ,
    \cby_1__1__14_chany_bottom_out[10] ,
    \cby_1__1__14_chany_bottom_out[11] ,
    \cby_1__1__14_chany_bottom_out[12] ,
    \cby_1__1__14_chany_bottom_out[13] ,
    \cby_1__1__14_chany_bottom_out[14] ,
    \cby_1__1__14_chany_bottom_out[15] ,
    \cby_1__1__14_chany_bottom_out[16] ,
    \cby_1__1__14_chany_bottom_out[17] ,
    \cby_1__1__14_chany_bottom_out[18] ,
    \cby_1__1__14_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__13_chany_bottom_out[0] ,
    \sb_1__1__13_chany_bottom_out[1] ,
    \sb_1__1__13_chany_bottom_out[2] ,
    \sb_1__1__13_chany_bottom_out[3] ,
    \sb_1__1__13_chany_bottom_out[4] ,
    \sb_1__1__13_chany_bottom_out[5] ,
    \sb_1__1__13_chany_bottom_out[6] ,
    \sb_1__1__13_chany_bottom_out[7] ,
    \sb_1__1__13_chany_bottom_out[8] ,
    \sb_1__1__13_chany_bottom_out[9] ,
    \sb_1__1__13_chany_bottom_out[10] ,
    \sb_1__1__13_chany_bottom_out[11] ,
    \sb_1__1__13_chany_bottom_out[12] ,
    \sb_1__1__13_chany_bottom_out[13] ,
    \sb_1__1__13_chany_bottom_out[14] ,
    \sb_1__1__13_chany_bottom_out[15] ,
    \sb_1__1__13_chany_bottom_out[16] ,
    \sb_1__1__13_chany_bottom_out[17] ,
    \sb_1__1__13_chany_bottom_out[18] ,
    \sb_1__1__13_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__14_chany_top_out[0] ,
    \cby_1__1__14_chany_top_out[1] ,
    \cby_1__1__14_chany_top_out[2] ,
    \cby_1__1__14_chany_top_out[3] ,
    \cby_1__1__14_chany_top_out[4] ,
    \cby_1__1__14_chany_top_out[5] ,
    \cby_1__1__14_chany_top_out[6] ,
    \cby_1__1__14_chany_top_out[7] ,
    \cby_1__1__14_chany_top_out[8] ,
    \cby_1__1__14_chany_top_out[9] ,
    \cby_1__1__14_chany_top_out[10] ,
    \cby_1__1__14_chany_top_out[11] ,
    \cby_1__1__14_chany_top_out[12] ,
    \cby_1__1__14_chany_top_out[13] ,
    \cby_1__1__14_chany_top_out[14] ,
    \cby_1__1__14_chany_top_out[15] ,
    \cby_1__1__14_chany_top_out[16] ,
    \cby_1__1__14_chany_top_out[17] ,
    \cby_1__1__14_chany_top_out[18] ,
    \cby_1__1__14_chany_top_out[19] }));
 cby_1__1_ cby_2__8_ (.Test_en_E_in(\Test_enWires[118] ),
    .Test_en_S_in(\Test_enWires[118] ),
    .Test_en_W_in(\Test_enWires[118] ),
    .Test_en_W_out(\Test_enWires[115] ),
    .ccff_head(grid_clb_15_ccff_tail),
    .ccff_tail(cby_1__1__15_ccff_tail),
    .left_grid_pin_16_(cby_1__1__15_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__15_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__15_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__15_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__15_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__15_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__15_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__15_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__15_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__15_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__15_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__15_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__15_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__15_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__15_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__15_left_grid_pin_31_),
    .prog_clk_0_N_out(\prog_clk_0_wires[68] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[66] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[65] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__13_chany_top_out[0] ,
    \sb_1__1__13_chany_top_out[1] ,
    \sb_1__1__13_chany_top_out[2] ,
    \sb_1__1__13_chany_top_out[3] ,
    \sb_1__1__13_chany_top_out[4] ,
    \sb_1__1__13_chany_top_out[5] ,
    \sb_1__1__13_chany_top_out[6] ,
    \sb_1__1__13_chany_top_out[7] ,
    \sb_1__1__13_chany_top_out[8] ,
    \sb_1__1__13_chany_top_out[9] ,
    \sb_1__1__13_chany_top_out[10] ,
    \sb_1__1__13_chany_top_out[11] ,
    \sb_1__1__13_chany_top_out[12] ,
    \sb_1__1__13_chany_top_out[13] ,
    \sb_1__1__13_chany_top_out[14] ,
    \sb_1__1__13_chany_top_out[15] ,
    \sb_1__1__13_chany_top_out[16] ,
    \sb_1__1__13_chany_top_out[17] ,
    \sb_1__1__13_chany_top_out[18] ,
    \sb_1__1__13_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__15_chany_bottom_out[0] ,
    \cby_1__1__15_chany_bottom_out[1] ,
    \cby_1__1__15_chany_bottom_out[2] ,
    \cby_1__1__15_chany_bottom_out[3] ,
    \cby_1__1__15_chany_bottom_out[4] ,
    \cby_1__1__15_chany_bottom_out[5] ,
    \cby_1__1__15_chany_bottom_out[6] ,
    \cby_1__1__15_chany_bottom_out[7] ,
    \cby_1__1__15_chany_bottom_out[8] ,
    \cby_1__1__15_chany_bottom_out[9] ,
    \cby_1__1__15_chany_bottom_out[10] ,
    \cby_1__1__15_chany_bottom_out[11] ,
    \cby_1__1__15_chany_bottom_out[12] ,
    \cby_1__1__15_chany_bottom_out[13] ,
    \cby_1__1__15_chany_bottom_out[14] ,
    \cby_1__1__15_chany_bottom_out[15] ,
    \cby_1__1__15_chany_bottom_out[16] ,
    \cby_1__1__15_chany_bottom_out[17] ,
    \cby_1__1__15_chany_bottom_out[18] ,
    \cby_1__1__15_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__8__1_chany_bottom_out[0] ,
    \sb_1__8__1_chany_bottom_out[1] ,
    \sb_1__8__1_chany_bottom_out[2] ,
    \sb_1__8__1_chany_bottom_out[3] ,
    \sb_1__8__1_chany_bottom_out[4] ,
    \sb_1__8__1_chany_bottom_out[5] ,
    \sb_1__8__1_chany_bottom_out[6] ,
    \sb_1__8__1_chany_bottom_out[7] ,
    \sb_1__8__1_chany_bottom_out[8] ,
    \sb_1__8__1_chany_bottom_out[9] ,
    \sb_1__8__1_chany_bottom_out[10] ,
    \sb_1__8__1_chany_bottom_out[11] ,
    \sb_1__8__1_chany_bottom_out[12] ,
    \sb_1__8__1_chany_bottom_out[13] ,
    \sb_1__8__1_chany_bottom_out[14] ,
    \sb_1__8__1_chany_bottom_out[15] ,
    \sb_1__8__1_chany_bottom_out[16] ,
    \sb_1__8__1_chany_bottom_out[17] ,
    \sb_1__8__1_chany_bottom_out[18] ,
    \sb_1__8__1_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__15_chany_top_out[0] ,
    \cby_1__1__15_chany_top_out[1] ,
    \cby_1__1__15_chany_top_out[2] ,
    \cby_1__1__15_chany_top_out[3] ,
    \cby_1__1__15_chany_top_out[4] ,
    \cby_1__1__15_chany_top_out[5] ,
    \cby_1__1__15_chany_top_out[6] ,
    \cby_1__1__15_chany_top_out[7] ,
    \cby_1__1__15_chany_top_out[8] ,
    \cby_1__1__15_chany_top_out[9] ,
    \cby_1__1__15_chany_top_out[10] ,
    \cby_1__1__15_chany_top_out[11] ,
    \cby_1__1__15_chany_top_out[12] ,
    \cby_1__1__15_chany_top_out[13] ,
    \cby_1__1__15_chany_top_out[14] ,
    \cby_1__1__15_chany_top_out[15] ,
    \cby_1__1__15_chany_top_out[16] ,
    \cby_1__1__15_chany_top_out[17] ,
    \cby_1__1__15_chany_top_out[18] ,
    \cby_1__1__15_chany_top_out[19] }));
 cby_1__1_ cby_3__1_ (.Test_en_E_in(\Test_enWires[22] ),
    .Test_en_S_in(\Test_enWires[22] ),
    .Test_en_W_in(\Test_enWires[22] ),
    .Test_en_W_out(\Test_enWires[19] ),
    .ccff_head(grid_clb_16_ccff_tail),
    .ccff_tail(cby_1__1__16_ccff_tail),
    .left_grid_pin_16_(cby_1__1__16_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__16_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__16_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__16_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__16_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__16_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__16_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__16_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__16_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__16_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__16_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__16_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__16_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__16_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__16_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__16_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[71] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[70] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__0__2_chany_top_out[0] ,
    \sb_1__0__2_chany_top_out[1] ,
    \sb_1__0__2_chany_top_out[2] ,
    \sb_1__0__2_chany_top_out[3] ,
    \sb_1__0__2_chany_top_out[4] ,
    \sb_1__0__2_chany_top_out[5] ,
    \sb_1__0__2_chany_top_out[6] ,
    \sb_1__0__2_chany_top_out[7] ,
    \sb_1__0__2_chany_top_out[8] ,
    \sb_1__0__2_chany_top_out[9] ,
    \sb_1__0__2_chany_top_out[10] ,
    \sb_1__0__2_chany_top_out[11] ,
    \sb_1__0__2_chany_top_out[12] ,
    \sb_1__0__2_chany_top_out[13] ,
    \sb_1__0__2_chany_top_out[14] ,
    \sb_1__0__2_chany_top_out[15] ,
    \sb_1__0__2_chany_top_out[16] ,
    \sb_1__0__2_chany_top_out[17] ,
    \sb_1__0__2_chany_top_out[18] ,
    \sb_1__0__2_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__16_chany_bottom_out[0] ,
    \cby_1__1__16_chany_bottom_out[1] ,
    \cby_1__1__16_chany_bottom_out[2] ,
    \cby_1__1__16_chany_bottom_out[3] ,
    \cby_1__1__16_chany_bottom_out[4] ,
    \cby_1__1__16_chany_bottom_out[5] ,
    \cby_1__1__16_chany_bottom_out[6] ,
    \cby_1__1__16_chany_bottom_out[7] ,
    \cby_1__1__16_chany_bottom_out[8] ,
    \cby_1__1__16_chany_bottom_out[9] ,
    \cby_1__1__16_chany_bottom_out[10] ,
    \cby_1__1__16_chany_bottom_out[11] ,
    \cby_1__1__16_chany_bottom_out[12] ,
    \cby_1__1__16_chany_bottom_out[13] ,
    \cby_1__1__16_chany_bottom_out[14] ,
    \cby_1__1__16_chany_bottom_out[15] ,
    \cby_1__1__16_chany_bottom_out[16] ,
    \cby_1__1__16_chany_bottom_out[17] ,
    \cby_1__1__16_chany_bottom_out[18] ,
    \cby_1__1__16_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__14_chany_bottom_out[0] ,
    \sb_1__1__14_chany_bottom_out[1] ,
    \sb_1__1__14_chany_bottom_out[2] ,
    \sb_1__1__14_chany_bottom_out[3] ,
    \sb_1__1__14_chany_bottom_out[4] ,
    \sb_1__1__14_chany_bottom_out[5] ,
    \sb_1__1__14_chany_bottom_out[6] ,
    \sb_1__1__14_chany_bottom_out[7] ,
    \sb_1__1__14_chany_bottom_out[8] ,
    \sb_1__1__14_chany_bottom_out[9] ,
    \sb_1__1__14_chany_bottom_out[10] ,
    \sb_1__1__14_chany_bottom_out[11] ,
    \sb_1__1__14_chany_bottom_out[12] ,
    \sb_1__1__14_chany_bottom_out[13] ,
    \sb_1__1__14_chany_bottom_out[14] ,
    \sb_1__1__14_chany_bottom_out[15] ,
    \sb_1__1__14_chany_bottom_out[16] ,
    \sb_1__1__14_chany_bottom_out[17] ,
    \sb_1__1__14_chany_bottom_out[18] ,
    \sb_1__1__14_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__16_chany_top_out[0] ,
    \cby_1__1__16_chany_top_out[1] ,
    \cby_1__1__16_chany_top_out[2] ,
    \cby_1__1__16_chany_top_out[3] ,
    \cby_1__1__16_chany_top_out[4] ,
    \cby_1__1__16_chany_top_out[5] ,
    \cby_1__1__16_chany_top_out[6] ,
    \cby_1__1__16_chany_top_out[7] ,
    \cby_1__1__16_chany_top_out[8] ,
    \cby_1__1__16_chany_top_out[9] ,
    \cby_1__1__16_chany_top_out[10] ,
    \cby_1__1__16_chany_top_out[11] ,
    \cby_1__1__16_chany_top_out[12] ,
    \cby_1__1__16_chany_top_out[13] ,
    \cby_1__1__16_chany_top_out[14] ,
    \cby_1__1__16_chany_top_out[15] ,
    \cby_1__1__16_chany_top_out[16] ,
    \cby_1__1__16_chany_top_out[17] ,
    \cby_1__1__16_chany_top_out[18] ,
    \cby_1__1__16_chany_top_out[19] }));
 cby_1__1_ cby_3__2_ (.Test_en_E_in(\Test_enWires[36] ),
    .Test_en_S_in(\Test_enWires[36] ),
    .Test_en_W_in(\Test_enWires[36] ),
    .Test_en_W_out(\Test_enWires[33] ),
    .ccff_head(grid_clb_17_ccff_tail),
    .ccff_tail(cby_1__1__17_ccff_tail),
    .clk_2_S_in(\clk_2_wires[11] ),
    .clk_2_S_out(\clk_2_wires[12] ),
    .left_grid_pin_16_(cby_1__1__17_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__17_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__17_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__17_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__17_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__17_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__17_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__17_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__17_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__17_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__17_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__17_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__17_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__17_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__17_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__17_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[74] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[73] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[11] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[12] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__14_chany_top_out[0] ,
    \sb_1__1__14_chany_top_out[1] ,
    \sb_1__1__14_chany_top_out[2] ,
    \sb_1__1__14_chany_top_out[3] ,
    \sb_1__1__14_chany_top_out[4] ,
    \sb_1__1__14_chany_top_out[5] ,
    \sb_1__1__14_chany_top_out[6] ,
    \sb_1__1__14_chany_top_out[7] ,
    \sb_1__1__14_chany_top_out[8] ,
    \sb_1__1__14_chany_top_out[9] ,
    \sb_1__1__14_chany_top_out[10] ,
    \sb_1__1__14_chany_top_out[11] ,
    \sb_1__1__14_chany_top_out[12] ,
    \sb_1__1__14_chany_top_out[13] ,
    \sb_1__1__14_chany_top_out[14] ,
    \sb_1__1__14_chany_top_out[15] ,
    \sb_1__1__14_chany_top_out[16] ,
    \sb_1__1__14_chany_top_out[17] ,
    \sb_1__1__14_chany_top_out[18] ,
    \sb_1__1__14_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__17_chany_bottom_out[0] ,
    \cby_1__1__17_chany_bottom_out[1] ,
    \cby_1__1__17_chany_bottom_out[2] ,
    \cby_1__1__17_chany_bottom_out[3] ,
    \cby_1__1__17_chany_bottom_out[4] ,
    \cby_1__1__17_chany_bottom_out[5] ,
    \cby_1__1__17_chany_bottom_out[6] ,
    \cby_1__1__17_chany_bottom_out[7] ,
    \cby_1__1__17_chany_bottom_out[8] ,
    \cby_1__1__17_chany_bottom_out[9] ,
    \cby_1__1__17_chany_bottom_out[10] ,
    \cby_1__1__17_chany_bottom_out[11] ,
    \cby_1__1__17_chany_bottom_out[12] ,
    \cby_1__1__17_chany_bottom_out[13] ,
    \cby_1__1__17_chany_bottom_out[14] ,
    \cby_1__1__17_chany_bottom_out[15] ,
    \cby_1__1__17_chany_bottom_out[16] ,
    \cby_1__1__17_chany_bottom_out[17] ,
    \cby_1__1__17_chany_bottom_out[18] ,
    \cby_1__1__17_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__15_chany_bottom_out[0] ,
    \sb_1__1__15_chany_bottom_out[1] ,
    \sb_1__1__15_chany_bottom_out[2] ,
    \sb_1__1__15_chany_bottom_out[3] ,
    \sb_1__1__15_chany_bottom_out[4] ,
    \sb_1__1__15_chany_bottom_out[5] ,
    \sb_1__1__15_chany_bottom_out[6] ,
    \sb_1__1__15_chany_bottom_out[7] ,
    \sb_1__1__15_chany_bottom_out[8] ,
    \sb_1__1__15_chany_bottom_out[9] ,
    \sb_1__1__15_chany_bottom_out[10] ,
    \sb_1__1__15_chany_bottom_out[11] ,
    \sb_1__1__15_chany_bottom_out[12] ,
    \sb_1__1__15_chany_bottom_out[13] ,
    \sb_1__1__15_chany_bottom_out[14] ,
    \sb_1__1__15_chany_bottom_out[15] ,
    \sb_1__1__15_chany_bottom_out[16] ,
    \sb_1__1__15_chany_bottom_out[17] ,
    \sb_1__1__15_chany_bottom_out[18] ,
    \sb_1__1__15_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__17_chany_top_out[0] ,
    \cby_1__1__17_chany_top_out[1] ,
    \cby_1__1__17_chany_top_out[2] ,
    \cby_1__1__17_chany_top_out[3] ,
    \cby_1__1__17_chany_top_out[4] ,
    \cby_1__1__17_chany_top_out[5] ,
    \cby_1__1__17_chany_top_out[6] ,
    \cby_1__1__17_chany_top_out[7] ,
    \cby_1__1__17_chany_top_out[8] ,
    \cby_1__1__17_chany_top_out[9] ,
    \cby_1__1__17_chany_top_out[10] ,
    \cby_1__1__17_chany_top_out[11] ,
    \cby_1__1__17_chany_top_out[12] ,
    \cby_1__1__17_chany_top_out[13] ,
    \cby_1__1__17_chany_top_out[14] ,
    \cby_1__1__17_chany_top_out[15] ,
    \cby_1__1__17_chany_top_out[16] ,
    \cby_1__1__17_chany_top_out[17] ,
    \cby_1__1__17_chany_top_out[18] ,
    \cby_1__1__17_chany_top_out[19] }));
 cby_1__1_ cby_3__3_ (.Test_en_E_in(\Test_enWires[50] ),
    .Test_en_S_in(\Test_enWires[50] ),
    .Test_en_W_in(\Test_enWires[50] ),
    .Test_en_W_out(\Test_enWires[47] ),
    .ccff_head(grid_clb_18_ccff_tail),
    .ccff_tail(cby_1__1__18_ccff_tail),
    .clk_2_N_out(\clk_2_wires[10] ),
    .clk_2_S_in(\clk_2_wires[9] ),
    .left_grid_pin_16_(cby_1__1__18_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__18_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__18_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__18_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__18_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__18_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__18_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__18_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__18_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__18_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__18_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__18_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__18_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__18_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__18_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__18_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[77] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[76] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[10] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[9] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__15_chany_top_out[0] ,
    \sb_1__1__15_chany_top_out[1] ,
    \sb_1__1__15_chany_top_out[2] ,
    \sb_1__1__15_chany_top_out[3] ,
    \sb_1__1__15_chany_top_out[4] ,
    \sb_1__1__15_chany_top_out[5] ,
    \sb_1__1__15_chany_top_out[6] ,
    \sb_1__1__15_chany_top_out[7] ,
    \sb_1__1__15_chany_top_out[8] ,
    \sb_1__1__15_chany_top_out[9] ,
    \sb_1__1__15_chany_top_out[10] ,
    \sb_1__1__15_chany_top_out[11] ,
    \sb_1__1__15_chany_top_out[12] ,
    \sb_1__1__15_chany_top_out[13] ,
    \sb_1__1__15_chany_top_out[14] ,
    \sb_1__1__15_chany_top_out[15] ,
    \sb_1__1__15_chany_top_out[16] ,
    \sb_1__1__15_chany_top_out[17] ,
    \sb_1__1__15_chany_top_out[18] ,
    \sb_1__1__15_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__18_chany_bottom_out[0] ,
    \cby_1__1__18_chany_bottom_out[1] ,
    \cby_1__1__18_chany_bottom_out[2] ,
    \cby_1__1__18_chany_bottom_out[3] ,
    \cby_1__1__18_chany_bottom_out[4] ,
    \cby_1__1__18_chany_bottom_out[5] ,
    \cby_1__1__18_chany_bottom_out[6] ,
    \cby_1__1__18_chany_bottom_out[7] ,
    \cby_1__1__18_chany_bottom_out[8] ,
    \cby_1__1__18_chany_bottom_out[9] ,
    \cby_1__1__18_chany_bottom_out[10] ,
    \cby_1__1__18_chany_bottom_out[11] ,
    \cby_1__1__18_chany_bottom_out[12] ,
    \cby_1__1__18_chany_bottom_out[13] ,
    \cby_1__1__18_chany_bottom_out[14] ,
    \cby_1__1__18_chany_bottom_out[15] ,
    \cby_1__1__18_chany_bottom_out[16] ,
    \cby_1__1__18_chany_bottom_out[17] ,
    \cby_1__1__18_chany_bottom_out[18] ,
    \cby_1__1__18_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__16_chany_bottom_out[0] ,
    \sb_1__1__16_chany_bottom_out[1] ,
    \sb_1__1__16_chany_bottom_out[2] ,
    \sb_1__1__16_chany_bottom_out[3] ,
    \sb_1__1__16_chany_bottom_out[4] ,
    \sb_1__1__16_chany_bottom_out[5] ,
    \sb_1__1__16_chany_bottom_out[6] ,
    \sb_1__1__16_chany_bottom_out[7] ,
    \sb_1__1__16_chany_bottom_out[8] ,
    \sb_1__1__16_chany_bottom_out[9] ,
    \sb_1__1__16_chany_bottom_out[10] ,
    \sb_1__1__16_chany_bottom_out[11] ,
    \sb_1__1__16_chany_bottom_out[12] ,
    \sb_1__1__16_chany_bottom_out[13] ,
    \sb_1__1__16_chany_bottom_out[14] ,
    \sb_1__1__16_chany_bottom_out[15] ,
    \sb_1__1__16_chany_bottom_out[16] ,
    \sb_1__1__16_chany_bottom_out[17] ,
    \sb_1__1__16_chany_bottom_out[18] ,
    \sb_1__1__16_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__18_chany_top_out[0] ,
    \cby_1__1__18_chany_top_out[1] ,
    \cby_1__1__18_chany_top_out[2] ,
    \cby_1__1__18_chany_top_out[3] ,
    \cby_1__1__18_chany_top_out[4] ,
    \cby_1__1__18_chany_top_out[5] ,
    \cby_1__1__18_chany_top_out[6] ,
    \cby_1__1__18_chany_top_out[7] ,
    \cby_1__1__18_chany_top_out[8] ,
    \cby_1__1__18_chany_top_out[9] ,
    \cby_1__1__18_chany_top_out[10] ,
    \cby_1__1__18_chany_top_out[11] ,
    \cby_1__1__18_chany_top_out[12] ,
    \cby_1__1__18_chany_top_out[13] ,
    \cby_1__1__18_chany_top_out[14] ,
    \cby_1__1__18_chany_top_out[15] ,
    \cby_1__1__18_chany_top_out[16] ,
    \cby_1__1__18_chany_top_out[17] ,
    \cby_1__1__18_chany_top_out[18] ,
    \cby_1__1__18_chany_top_out[19] }));
 cby_1__1_ cby_3__4_ (.Test_en_E_in(\Test_enWires[64] ),
    .Test_en_S_in(\Test_enWires[64] ),
    .Test_en_W_in(\Test_enWires[64] ),
    .Test_en_W_out(\Test_enWires[61] ),
    .ccff_head(grid_clb_19_ccff_tail),
    .ccff_tail(cby_1__1__19_ccff_tail),
    .left_grid_pin_16_(cby_1__1__19_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__19_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__19_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__19_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__19_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__19_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__19_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__19_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__19_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__19_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__19_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__19_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__19_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__19_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__19_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__19_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[80] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[79] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__16_chany_top_out[0] ,
    \sb_1__1__16_chany_top_out[1] ,
    \sb_1__1__16_chany_top_out[2] ,
    \sb_1__1__16_chany_top_out[3] ,
    \sb_1__1__16_chany_top_out[4] ,
    \sb_1__1__16_chany_top_out[5] ,
    \sb_1__1__16_chany_top_out[6] ,
    \sb_1__1__16_chany_top_out[7] ,
    \sb_1__1__16_chany_top_out[8] ,
    \sb_1__1__16_chany_top_out[9] ,
    \sb_1__1__16_chany_top_out[10] ,
    \sb_1__1__16_chany_top_out[11] ,
    \sb_1__1__16_chany_top_out[12] ,
    \sb_1__1__16_chany_top_out[13] ,
    \sb_1__1__16_chany_top_out[14] ,
    \sb_1__1__16_chany_top_out[15] ,
    \sb_1__1__16_chany_top_out[16] ,
    \sb_1__1__16_chany_top_out[17] ,
    \sb_1__1__16_chany_top_out[18] ,
    \sb_1__1__16_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__19_chany_bottom_out[0] ,
    \cby_1__1__19_chany_bottom_out[1] ,
    \cby_1__1__19_chany_bottom_out[2] ,
    \cby_1__1__19_chany_bottom_out[3] ,
    \cby_1__1__19_chany_bottom_out[4] ,
    \cby_1__1__19_chany_bottom_out[5] ,
    \cby_1__1__19_chany_bottom_out[6] ,
    \cby_1__1__19_chany_bottom_out[7] ,
    \cby_1__1__19_chany_bottom_out[8] ,
    \cby_1__1__19_chany_bottom_out[9] ,
    \cby_1__1__19_chany_bottom_out[10] ,
    \cby_1__1__19_chany_bottom_out[11] ,
    \cby_1__1__19_chany_bottom_out[12] ,
    \cby_1__1__19_chany_bottom_out[13] ,
    \cby_1__1__19_chany_bottom_out[14] ,
    \cby_1__1__19_chany_bottom_out[15] ,
    \cby_1__1__19_chany_bottom_out[16] ,
    \cby_1__1__19_chany_bottom_out[17] ,
    \cby_1__1__19_chany_bottom_out[18] ,
    \cby_1__1__19_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__17_chany_bottom_out[0] ,
    \sb_1__1__17_chany_bottom_out[1] ,
    \sb_1__1__17_chany_bottom_out[2] ,
    \sb_1__1__17_chany_bottom_out[3] ,
    \sb_1__1__17_chany_bottom_out[4] ,
    \sb_1__1__17_chany_bottom_out[5] ,
    \sb_1__1__17_chany_bottom_out[6] ,
    \sb_1__1__17_chany_bottom_out[7] ,
    \sb_1__1__17_chany_bottom_out[8] ,
    \sb_1__1__17_chany_bottom_out[9] ,
    \sb_1__1__17_chany_bottom_out[10] ,
    \sb_1__1__17_chany_bottom_out[11] ,
    \sb_1__1__17_chany_bottom_out[12] ,
    \sb_1__1__17_chany_bottom_out[13] ,
    \sb_1__1__17_chany_bottom_out[14] ,
    \sb_1__1__17_chany_bottom_out[15] ,
    \sb_1__1__17_chany_bottom_out[16] ,
    \sb_1__1__17_chany_bottom_out[17] ,
    \sb_1__1__17_chany_bottom_out[18] ,
    \sb_1__1__17_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__19_chany_top_out[0] ,
    \cby_1__1__19_chany_top_out[1] ,
    \cby_1__1__19_chany_top_out[2] ,
    \cby_1__1__19_chany_top_out[3] ,
    \cby_1__1__19_chany_top_out[4] ,
    \cby_1__1__19_chany_top_out[5] ,
    \cby_1__1__19_chany_top_out[6] ,
    \cby_1__1__19_chany_top_out[7] ,
    \cby_1__1__19_chany_top_out[8] ,
    \cby_1__1__19_chany_top_out[9] ,
    \cby_1__1__19_chany_top_out[10] ,
    \cby_1__1__19_chany_top_out[11] ,
    \cby_1__1__19_chany_top_out[12] ,
    \cby_1__1__19_chany_top_out[13] ,
    \cby_1__1__19_chany_top_out[14] ,
    \cby_1__1__19_chany_top_out[15] ,
    \cby_1__1__19_chany_top_out[16] ,
    \cby_1__1__19_chany_top_out[17] ,
    \cby_1__1__19_chany_top_out[18] ,
    \cby_1__1__19_chany_top_out[19] }));
 cby_1__1_ cby_3__5_ (.Test_en_E_in(\Test_enWires[78] ),
    .Test_en_S_in(\Test_enWires[78] ),
    .Test_en_W_in(\Test_enWires[78] ),
    .Test_en_W_out(\Test_enWires[75] ),
    .ccff_head(grid_clb_20_ccff_tail),
    .ccff_tail(cby_1__1__20_ccff_tail),
    .left_grid_pin_16_(cby_1__1__20_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__20_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__20_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__20_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__20_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__20_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__20_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__20_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__20_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__20_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__20_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__20_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__20_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__20_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__20_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__20_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[83] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[82] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__17_chany_top_out[0] ,
    \sb_1__1__17_chany_top_out[1] ,
    \sb_1__1__17_chany_top_out[2] ,
    \sb_1__1__17_chany_top_out[3] ,
    \sb_1__1__17_chany_top_out[4] ,
    \sb_1__1__17_chany_top_out[5] ,
    \sb_1__1__17_chany_top_out[6] ,
    \sb_1__1__17_chany_top_out[7] ,
    \sb_1__1__17_chany_top_out[8] ,
    \sb_1__1__17_chany_top_out[9] ,
    \sb_1__1__17_chany_top_out[10] ,
    \sb_1__1__17_chany_top_out[11] ,
    \sb_1__1__17_chany_top_out[12] ,
    \sb_1__1__17_chany_top_out[13] ,
    \sb_1__1__17_chany_top_out[14] ,
    \sb_1__1__17_chany_top_out[15] ,
    \sb_1__1__17_chany_top_out[16] ,
    \sb_1__1__17_chany_top_out[17] ,
    \sb_1__1__17_chany_top_out[18] ,
    \sb_1__1__17_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__20_chany_bottom_out[0] ,
    \cby_1__1__20_chany_bottom_out[1] ,
    \cby_1__1__20_chany_bottom_out[2] ,
    \cby_1__1__20_chany_bottom_out[3] ,
    \cby_1__1__20_chany_bottom_out[4] ,
    \cby_1__1__20_chany_bottom_out[5] ,
    \cby_1__1__20_chany_bottom_out[6] ,
    \cby_1__1__20_chany_bottom_out[7] ,
    \cby_1__1__20_chany_bottom_out[8] ,
    \cby_1__1__20_chany_bottom_out[9] ,
    \cby_1__1__20_chany_bottom_out[10] ,
    \cby_1__1__20_chany_bottom_out[11] ,
    \cby_1__1__20_chany_bottom_out[12] ,
    \cby_1__1__20_chany_bottom_out[13] ,
    \cby_1__1__20_chany_bottom_out[14] ,
    \cby_1__1__20_chany_bottom_out[15] ,
    \cby_1__1__20_chany_bottom_out[16] ,
    \cby_1__1__20_chany_bottom_out[17] ,
    \cby_1__1__20_chany_bottom_out[18] ,
    \cby_1__1__20_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__18_chany_bottom_out[0] ,
    \sb_1__1__18_chany_bottom_out[1] ,
    \sb_1__1__18_chany_bottom_out[2] ,
    \sb_1__1__18_chany_bottom_out[3] ,
    \sb_1__1__18_chany_bottom_out[4] ,
    \sb_1__1__18_chany_bottom_out[5] ,
    \sb_1__1__18_chany_bottom_out[6] ,
    \sb_1__1__18_chany_bottom_out[7] ,
    \sb_1__1__18_chany_bottom_out[8] ,
    \sb_1__1__18_chany_bottom_out[9] ,
    \sb_1__1__18_chany_bottom_out[10] ,
    \sb_1__1__18_chany_bottom_out[11] ,
    \sb_1__1__18_chany_bottom_out[12] ,
    \sb_1__1__18_chany_bottom_out[13] ,
    \sb_1__1__18_chany_bottom_out[14] ,
    \sb_1__1__18_chany_bottom_out[15] ,
    \sb_1__1__18_chany_bottom_out[16] ,
    \sb_1__1__18_chany_bottom_out[17] ,
    \sb_1__1__18_chany_bottom_out[18] ,
    \sb_1__1__18_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__20_chany_top_out[0] ,
    \cby_1__1__20_chany_top_out[1] ,
    \cby_1__1__20_chany_top_out[2] ,
    \cby_1__1__20_chany_top_out[3] ,
    \cby_1__1__20_chany_top_out[4] ,
    \cby_1__1__20_chany_top_out[5] ,
    \cby_1__1__20_chany_top_out[6] ,
    \cby_1__1__20_chany_top_out[7] ,
    \cby_1__1__20_chany_top_out[8] ,
    \cby_1__1__20_chany_top_out[9] ,
    \cby_1__1__20_chany_top_out[10] ,
    \cby_1__1__20_chany_top_out[11] ,
    \cby_1__1__20_chany_top_out[12] ,
    \cby_1__1__20_chany_top_out[13] ,
    \cby_1__1__20_chany_top_out[14] ,
    \cby_1__1__20_chany_top_out[15] ,
    \cby_1__1__20_chany_top_out[16] ,
    \cby_1__1__20_chany_top_out[17] ,
    \cby_1__1__20_chany_top_out[18] ,
    \cby_1__1__20_chany_top_out[19] }));
 cby_1__1_ cby_3__6_ (.Test_en_E_in(\Test_enWires[92] ),
    .Test_en_S_in(\Test_enWires[92] ),
    .Test_en_W_in(\Test_enWires[92] ),
    .Test_en_W_out(\Test_enWires[89] ),
    .ccff_head(grid_clb_21_ccff_tail),
    .ccff_tail(cby_1__1__21_ccff_tail),
    .clk_2_S_in(\clk_2_wires[24] ),
    .clk_2_S_out(\clk_2_wires[25] ),
    .left_grid_pin_16_(cby_1__1__21_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__21_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__21_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__21_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__21_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__21_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__21_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__21_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__21_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__21_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__21_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__21_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__21_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__21_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__21_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__21_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[86] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[85] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[24] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[25] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__18_chany_top_out[0] ,
    \sb_1__1__18_chany_top_out[1] ,
    \sb_1__1__18_chany_top_out[2] ,
    \sb_1__1__18_chany_top_out[3] ,
    \sb_1__1__18_chany_top_out[4] ,
    \sb_1__1__18_chany_top_out[5] ,
    \sb_1__1__18_chany_top_out[6] ,
    \sb_1__1__18_chany_top_out[7] ,
    \sb_1__1__18_chany_top_out[8] ,
    \sb_1__1__18_chany_top_out[9] ,
    \sb_1__1__18_chany_top_out[10] ,
    \sb_1__1__18_chany_top_out[11] ,
    \sb_1__1__18_chany_top_out[12] ,
    \sb_1__1__18_chany_top_out[13] ,
    \sb_1__1__18_chany_top_out[14] ,
    \sb_1__1__18_chany_top_out[15] ,
    \sb_1__1__18_chany_top_out[16] ,
    \sb_1__1__18_chany_top_out[17] ,
    \sb_1__1__18_chany_top_out[18] ,
    \sb_1__1__18_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__21_chany_bottom_out[0] ,
    \cby_1__1__21_chany_bottom_out[1] ,
    \cby_1__1__21_chany_bottom_out[2] ,
    \cby_1__1__21_chany_bottom_out[3] ,
    \cby_1__1__21_chany_bottom_out[4] ,
    \cby_1__1__21_chany_bottom_out[5] ,
    \cby_1__1__21_chany_bottom_out[6] ,
    \cby_1__1__21_chany_bottom_out[7] ,
    \cby_1__1__21_chany_bottom_out[8] ,
    \cby_1__1__21_chany_bottom_out[9] ,
    \cby_1__1__21_chany_bottom_out[10] ,
    \cby_1__1__21_chany_bottom_out[11] ,
    \cby_1__1__21_chany_bottom_out[12] ,
    \cby_1__1__21_chany_bottom_out[13] ,
    \cby_1__1__21_chany_bottom_out[14] ,
    \cby_1__1__21_chany_bottom_out[15] ,
    \cby_1__1__21_chany_bottom_out[16] ,
    \cby_1__1__21_chany_bottom_out[17] ,
    \cby_1__1__21_chany_bottom_out[18] ,
    \cby_1__1__21_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__19_chany_bottom_out[0] ,
    \sb_1__1__19_chany_bottom_out[1] ,
    \sb_1__1__19_chany_bottom_out[2] ,
    \sb_1__1__19_chany_bottom_out[3] ,
    \sb_1__1__19_chany_bottom_out[4] ,
    \sb_1__1__19_chany_bottom_out[5] ,
    \sb_1__1__19_chany_bottom_out[6] ,
    \sb_1__1__19_chany_bottom_out[7] ,
    \sb_1__1__19_chany_bottom_out[8] ,
    \sb_1__1__19_chany_bottom_out[9] ,
    \sb_1__1__19_chany_bottom_out[10] ,
    \sb_1__1__19_chany_bottom_out[11] ,
    \sb_1__1__19_chany_bottom_out[12] ,
    \sb_1__1__19_chany_bottom_out[13] ,
    \sb_1__1__19_chany_bottom_out[14] ,
    \sb_1__1__19_chany_bottom_out[15] ,
    \sb_1__1__19_chany_bottom_out[16] ,
    \sb_1__1__19_chany_bottom_out[17] ,
    \sb_1__1__19_chany_bottom_out[18] ,
    \sb_1__1__19_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__21_chany_top_out[0] ,
    \cby_1__1__21_chany_top_out[1] ,
    \cby_1__1__21_chany_top_out[2] ,
    \cby_1__1__21_chany_top_out[3] ,
    \cby_1__1__21_chany_top_out[4] ,
    \cby_1__1__21_chany_top_out[5] ,
    \cby_1__1__21_chany_top_out[6] ,
    \cby_1__1__21_chany_top_out[7] ,
    \cby_1__1__21_chany_top_out[8] ,
    \cby_1__1__21_chany_top_out[9] ,
    \cby_1__1__21_chany_top_out[10] ,
    \cby_1__1__21_chany_top_out[11] ,
    \cby_1__1__21_chany_top_out[12] ,
    \cby_1__1__21_chany_top_out[13] ,
    \cby_1__1__21_chany_top_out[14] ,
    \cby_1__1__21_chany_top_out[15] ,
    \cby_1__1__21_chany_top_out[16] ,
    \cby_1__1__21_chany_top_out[17] ,
    \cby_1__1__21_chany_top_out[18] ,
    \cby_1__1__21_chany_top_out[19] }));
 cby_1__1_ cby_3__7_ (.Test_en_E_in(\Test_enWires[106] ),
    .Test_en_S_in(\Test_enWires[106] ),
    .Test_en_W_in(\Test_enWires[106] ),
    .Test_en_W_out(\Test_enWires[103] ),
    .ccff_head(grid_clb_22_ccff_tail),
    .ccff_tail(cby_1__1__22_ccff_tail),
    .clk_2_N_out(\clk_2_wires[23] ),
    .clk_2_S_in(\clk_2_wires[22] ),
    .left_grid_pin_16_(cby_1__1__22_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__22_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__22_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__22_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__22_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__22_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__22_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__22_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__22_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__22_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__22_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__22_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__22_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__22_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__22_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__22_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[89] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[88] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[23] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[22] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__19_chany_top_out[0] ,
    \sb_1__1__19_chany_top_out[1] ,
    \sb_1__1__19_chany_top_out[2] ,
    \sb_1__1__19_chany_top_out[3] ,
    \sb_1__1__19_chany_top_out[4] ,
    \sb_1__1__19_chany_top_out[5] ,
    \sb_1__1__19_chany_top_out[6] ,
    \sb_1__1__19_chany_top_out[7] ,
    \sb_1__1__19_chany_top_out[8] ,
    \sb_1__1__19_chany_top_out[9] ,
    \sb_1__1__19_chany_top_out[10] ,
    \sb_1__1__19_chany_top_out[11] ,
    \sb_1__1__19_chany_top_out[12] ,
    \sb_1__1__19_chany_top_out[13] ,
    \sb_1__1__19_chany_top_out[14] ,
    \sb_1__1__19_chany_top_out[15] ,
    \sb_1__1__19_chany_top_out[16] ,
    \sb_1__1__19_chany_top_out[17] ,
    \sb_1__1__19_chany_top_out[18] ,
    \sb_1__1__19_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__22_chany_bottom_out[0] ,
    \cby_1__1__22_chany_bottom_out[1] ,
    \cby_1__1__22_chany_bottom_out[2] ,
    \cby_1__1__22_chany_bottom_out[3] ,
    \cby_1__1__22_chany_bottom_out[4] ,
    \cby_1__1__22_chany_bottom_out[5] ,
    \cby_1__1__22_chany_bottom_out[6] ,
    \cby_1__1__22_chany_bottom_out[7] ,
    \cby_1__1__22_chany_bottom_out[8] ,
    \cby_1__1__22_chany_bottom_out[9] ,
    \cby_1__1__22_chany_bottom_out[10] ,
    \cby_1__1__22_chany_bottom_out[11] ,
    \cby_1__1__22_chany_bottom_out[12] ,
    \cby_1__1__22_chany_bottom_out[13] ,
    \cby_1__1__22_chany_bottom_out[14] ,
    \cby_1__1__22_chany_bottom_out[15] ,
    \cby_1__1__22_chany_bottom_out[16] ,
    \cby_1__1__22_chany_bottom_out[17] ,
    \cby_1__1__22_chany_bottom_out[18] ,
    \cby_1__1__22_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__20_chany_bottom_out[0] ,
    \sb_1__1__20_chany_bottom_out[1] ,
    \sb_1__1__20_chany_bottom_out[2] ,
    \sb_1__1__20_chany_bottom_out[3] ,
    \sb_1__1__20_chany_bottom_out[4] ,
    \sb_1__1__20_chany_bottom_out[5] ,
    \sb_1__1__20_chany_bottom_out[6] ,
    \sb_1__1__20_chany_bottom_out[7] ,
    \sb_1__1__20_chany_bottom_out[8] ,
    \sb_1__1__20_chany_bottom_out[9] ,
    \sb_1__1__20_chany_bottom_out[10] ,
    \sb_1__1__20_chany_bottom_out[11] ,
    \sb_1__1__20_chany_bottom_out[12] ,
    \sb_1__1__20_chany_bottom_out[13] ,
    \sb_1__1__20_chany_bottom_out[14] ,
    \sb_1__1__20_chany_bottom_out[15] ,
    \sb_1__1__20_chany_bottom_out[16] ,
    \sb_1__1__20_chany_bottom_out[17] ,
    \sb_1__1__20_chany_bottom_out[18] ,
    \sb_1__1__20_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__22_chany_top_out[0] ,
    \cby_1__1__22_chany_top_out[1] ,
    \cby_1__1__22_chany_top_out[2] ,
    \cby_1__1__22_chany_top_out[3] ,
    \cby_1__1__22_chany_top_out[4] ,
    \cby_1__1__22_chany_top_out[5] ,
    \cby_1__1__22_chany_top_out[6] ,
    \cby_1__1__22_chany_top_out[7] ,
    \cby_1__1__22_chany_top_out[8] ,
    \cby_1__1__22_chany_top_out[9] ,
    \cby_1__1__22_chany_top_out[10] ,
    \cby_1__1__22_chany_top_out[11] ,
    \cby_1__1__22_chany_top_out[12] ,
    \cby_1__1__22_chany_top_out[13] ,
    \cby_1__1__22_chany_top_out[14] ,
    \cby_1__1__22_chany_top_out[15] ,
    \cby_1__1__22_chany_top_out[16] ,
    \cby_1__1__22_chany_top_out[17] ,
    \cby_1__1__22_chany_top_out[18] ,
    \cby_1__1__22_chany_top_out[19] }));
 cby_1__1_ cby_3__8_ (.Test_en_E_in(\Test_enWires[120] ),
    .Test_en_S_in(\Test_enWires[120] ),
    .Test_en_W_in(\Test_enWires[120] ),
    .Test_en_W_out(\Test_enWires[117] ),
    .ccff_head(grid_clb_23_ccff_tail),
    .ccff_tail(cby_1__1__23_ccff_tail),
    .left_grid_pin_16_(cby_1__1__23_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__23_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__23_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__23_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__23_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__23_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__23_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__23_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__23_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__23_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__23_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__23_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__23_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__23_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__23_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__23_left_grid_pin_31_),
    .prog_clk_0_N_out(\prog_clk_0_wires[94] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[92] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[91] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__20_chany_top_out[0] ,
    \sb_1__1__20_chany_top_out[1] ,
    \sb_1__1__20_chany_top_out[2] ,
    \sb_1__1__20_chany_top_out[3] ,
    \sb_1__1__20_chany_top_out[4] ,
    \sb_1__1__20_chany_top_out[5] ,
    \sb_1__1__20_chany_top_out[6] ,
    \sb_1__1__20_chany_top_out[7] ,
    \sb_1__1__20_chany_top_out[8] ,
    \sb_1__1__20_chany_top_out[9] ,
    \sb_1__1__20_chany_top_out[10] ,
    \sb_1__1__20_chany_top_out[11] ,
    \sb_1__1__20_chany_top_out[12] ,
    \sb_1__1__20_chany_top_out[13] ,
    \sb_1__1__20_chany_top_out[14] ,
    \sb_1__1__20_chany_top_out[15] ,
    \sb_1__1__20_chany_top_out[16] ,
    \sb_1__1__20_chany_top_out[17] ,
    \sb_1__1__20_chany_top_out[18] ,
    \sb_1__1__20_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__23_chany_bottom_out[0] ,
    \cby_1__1__23_chany_bottom_out[1] ,
    \cby_1__1__23_chany_bottom_out[2] ,
    \cby_1__1__23_chany_bottom_out[3] ,
    \cby_1__1__23_chany_bottom_out[4] ,
    \cby_1__1__23_chany_bottom_out[5] ,
    \cby_1__1__23_chany_bottom_out[6] ,
    \cby_1__1__23_chany_bottom_out[7] ,
    \cby_1__1__23_chany_bottom_out[8] ,
    \cby_1__1__23_chany_bottom_out[9] ,
    \cby_1__1__23_chany_bottom_out[10] ,
    \cby_1__1__23_chany_bottom_out[11] ,
    \cby_1__1__23_chany_bottom_out[12] ,
    \cby_1__1__23_chany_bottom_out[13] ,
    \cby_1__1__23_chany_bottom_out[14] ,
    \cby_1__1__23_chany_bottom_out[15] ,
    \cby_1__1__23_chany_bottom_out[16] ,
    \cby_1__1__23_chany_bottom_out[17] ,
    \cby_1__1__23_chany_bottom_out[18] ,
    \cby_1__1__23_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__8__2_chany_bottom_out[0] ,
    \sb_1__8__2_chany_bottom_out[1] ,
    \sb_1__8__2_chany_bottom_out[2] ,
    \sb_1__8__2_chany_bottom_out[3] ,
    \sb_1__8__2_chany_bottom_out[4] ,
    \sb_1__8__2_chany_bottom_out[5] ,
    \sb_1__8__2_chany_bottom_out[6] ,
    \sb_1__8__2_chany_bottom_out[7] ,
    \sb_1__8__2_chany_bottom_out[8] ,
    \sb_1__8__2_chany_bottom_out[9] ,
    \sb_1__8__2_chany_bottom_out[10] ,
    \sb_1__8__2_chany_bottom_out[11] ,
    \sb_1__8__2_chany_bottom_out[12] ,
    \sb_1__8__2_chany_bottom_out[13] ,
    \sb_1__8__2_chany_bottom_out[14] ,
    \sb_1__8__2_chany_bottom_out[15] ,
    \sb_1__8__2_chany_bottom_out[16] ,
    \sb_1__8__2_chany_bottom_out[17] ,
    \sb_1__8__2_chany_bottom_out[18] ,
    \sb_1__8__2_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__23_chany_top_out[0] ,
    \cby_1__1__23_chany_top_out[1] ,
    \cby_1__1__23_chany_top_out[2] ,
    \cby_1__1__23_chany_top_out[3] ,
    \cby_1__1__23_chany_top_out[4] ,
    \cby_1__1__23_chany_top_out[5] ,
    \cby_1__1__23_chany_top_out[6] ,
    \cby_1__1__23_chany_top_out[7] ,
    \cby_1__1__23_chany_top_out[8] ,
    \cby_1__1__23_chany_top_out[9] ,
    \cby_1__1__23_chany_top_out[10] ,
    \cby_1__1__23_chany_top_out[11] ,
    \cby_1__1__23_chany_top_out[12] ,
    \cby_1__1__23_chany_top_out[13] ,
    \cby_1__1__23_chany_top_out[14] ,
    \cby_1__1__23_chany_top_out[15] ,
    \cby_1__1__23_chany_top_out[16] ,
    \cby_1__1__23_chany_top_out[17] ,
    \cby_1__1__23_chany_top_out[18] ,
    \cby_1__1__23_chany_top_out[19] }));
 cby_1__1_ cby_4__1_ (.Test_en_E_in(\Test_enWires[1] ),
    .Test_en_E_out(\Test_enWires[23] ),
    .Test_en_N_out(\Test_enWires[2] ),
    .Test_en_S_in(\Test_enWires[1] ),
    .Test_en_W_in(\Test_enWires[1] ),
    .Test_en_W_out(\Test_enWires[21] ),
    .ccff_head(grid_clb_24_ccff_tail),
    .ccff_tail(cby_1__1__24_ccff_tail),
    .clk_3_N_out(\clk_3_wires[27] ),
    .clk_3_S_in(\clk_3_wires[28] ),
    .left_grid_pin_16_(cby_1__1__24_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__24_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__24_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__24_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__24_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__24_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__24_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__24_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__24_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__24_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__24_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__24_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__24_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__24_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__24_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__24_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[97] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[96] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[27] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[28] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__0__3_chany_top_out[0] ,
    \sb_1__0__3_chany_top_out[1] ,
    \sb_1__0__3_chany_top_out[2] ,
    \sb_1__0__3_chany_top_out[3] ,
    \sb_1__0__3_chany_top_out[4] ,
    \sb_1__0__3_chany_top_out[5] ,
    \sb_1__0__3_chany_top_out[6] ,
    \sb_1__0__3_chany_top_out[7] ,
    \sb_1__0__3_chany_top_out[8] ,
    \sb_1__0__3_chany_top_out[9] ,
    \sb_1__0__3_chany_top_out[10] ,
    \sb_1__0__3_chany_top_out[11] ,
    \sb_1__0__3_chany_top_out[12] ,
    \sb_1__0__3_chany_top_out[13] ,
    \sb_1__0__3_chany_top_out[14] ,
    \sb_1__0__3_chany_top_out[15] ,
    \sb_1__0__3_chany_top_out[16] ,
    \sb_1__0__3_chany_top_out[17] ,
    \sb_1__0__3_chany_top_out[18] ,
    \sb_1__0__3_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__24_chany_bottom_out[0] ,
    \cby_1__1__24_chany_bottom_out[1] ,
    \cby_1__1__24_chany_bottom_out[2] ,
    \cby_1__1__24_chany_bottom_out[3] ,
    \cby_1__1__24_chany_bottom_out[4] ,
    \cby_1__1__24_chany_bottom_out[5] ,
    \cby_1__1__24_chany_bottom_out[6] ,
    \cby_1__1__24_chany_bottom_out[7] ,
    \cby_1__1__24_chany_bottom_out[8] ,
    \cby_1__1__24_chany_bottom_out[9] ,
    \cby_1__1__24_chany_bottom_out[10] ,
    \cby_1__1__24_chany_bottom_out[11] ,
    \cby_1__1__24_chany_bottom_out[12] ,
    \cby_1__1__24_chany_bottom_out[13] ,
    \cby_1__1__24_chany_bottom_out[14] ,
    \cby_1__1__24_chany_bottom_out[15] ,
    \cby_1__1__24_chany_bottom_out[16] ,
    \cby_1__1__24_chany_bottom_out[17] ,
    \cby_1__1__24_chany_bottom_out[18] ,
    \cby_1__1__24_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__21_chany_bottom_out[0] ,
    \sb_1__1__21_chany_bottom_out[1] ,
    \sb_1__1__21_chany_bottom_out[2] ,
    \sb_1__1__21_chany_bottom_out[3] ,
    \sb_1__1__21_chany_bottom_out[4] ,
    \sb_1__1__21_chany_bottom_out[5] ,
    \sb_1__1__21_chany_bottom_out[6] ,
    \sb_1__1__21_chany_bottom_out[7] ,
    \sb_1__1__21_chany_bottom_out[8] ,
    \sb_1__1__21_chany_bottom_out[9] ,
    \sb_1__1__21_chany_bottom_out[10] ,
    \sb_1__1__21_chany_bottom_out[11] ,
    \sb_1__1__21_chany_bottom_out[12] ,
    \sb_1__1__21_chany_bottom_out[13] ,
    \sb_1__1__21_chany_bottom_out[14] ,
    \sb_1__1__21_chany_bottom_out[15] ,
    \sb_1__1__21_chany_bottom_out[16] ,
    \sb_1__1__21_chany_bottom_out[17] ,
    \sb_1__1__21_chany_bottom_out[18] ,
    \sb_1__1__21_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__24_chany_top_out[0] ,
    \cby_1__1__24_chany_top_out[1] ,
    \cby_1__1__24_chany_top_out[2] ,
    \cby_1__1__24_chany_top_out[3] ,
    \cby_1__1__24_chany_top_out[4] ,
    \cby_1__1__24_chany_top_out[5] ,
    \cby_1__1__24_chany_top_out[6] ,
    \cby_1__1__24_chany_top_out[7] ,
    \cby_1__1__24_chany_top_out[8] ,
    \cby_1__1__24_chany_top_out[9] ,
    \cby_1__1__24_chany_top_out[10] ,
    \cby_1__1__24_chany_top_out[11] ,
    \cby_1__1__24_chany_top_out[12] ,
    \cby_1__1__24_chany_top_out[13] ,
    \cby_1__1__24_chany_top_out[14] ,
    \cby_1__1__24_chany_top_out[15] ,
    \cby_1__1__24_chany_top_out[16] ,
    \cby_1__1__24_chany_top_out[17] ,
    \cby_1__1__24_chany_top_out[18] ,
    \cby_1__1__24_chany_top_out[19] }));
 cby_1__1_ cby_4__2_ (.Test_en_E_in(\Test_enWires[3] ),
    .Test_en_E_out(\Test_enWires[37] ),
    .Test_en_N_out(\Test_enWires[4] ),
    .Test_en_S_in(\Test_enWires[3] ),
    .Test_en_W_in(\Test_enWires[3] ),
    .Test_en_W_out(\Test_enWires[35] ),
    .ccff_head(grid_clb_25_ccff_tail),
    .ccff_tail(cby_1__1__25_ccff_tail),
    .clk_3_N_out(\clk_3_wires[29] ),
    .clk_3_S_in(\clk_3_wires[30] ),
    .left_grid_pin_16_(cby_1__1__25_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__25_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__25_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__25_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__25_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__25_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__25_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__25_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__25_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__25_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__25_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__25_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__25_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__25_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__25_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__25_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[100] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[99] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[29] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[30] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__21_chany_top_out[0] ,
    \sb_1__1__21_chany_top_out[1] ,
    \sb_1__1__21_chany_top_out[2] ,
    \sb_1__1__21_chany_top_out[3] ,
    \sb_1__1__21_chany_top_out[4] ,
    \sb_1__1__21_chany_top_out[5] ,
    \sb_1__1__21_chany_top_out[6] ,
    \sb_1__1__21_chany_top_out[7] ,
    \sb_1__1__21_chany_top_out[8] ,
    \sb_1__1__21_chany_top_out[9] ,
    \sb_1__1__21_chany_top_out[10] ,
    \sb_1__1__21_chany_top_out[11] ,
    \sb_1__1__21_chany_top_out[12] ,
    \sb_1__1__21_chany_top_out[13] ,
    \sb_1__1__21_chany_top_out[14] ,
    \sb_1__1__21_chany_top_out[15] ,
    \sb_1__1__21_chany_top_out[16] ,
    \sb_1__1__21_chany_top_out[17] ,
    \sb_1__1__21_chany_top_out[18] ,
    \sb_1__1__21_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__25_chany_bottom_out[0] ,
    \cby_1__1__25_chany_bottom_out[1] ,
    \cby_1__1__25_chany_bottom_out[2] ,
    \cby_1__1__25_chany_bottom_out[3] ,
    \cby_1__1__25_chany_bottom_out[4] ,
    \cby_1__1__25_chany_bottom_out[5] ,
    \cby_1__1__25_chany_bottom_out[6] ,
    \cby_1__1__25_chany_bottom_out[7] ,
    \cby_1__1__25_chany_bottom_out[8] ,
    \cby_1__1__25_chany_bottom_out[9] ,
    \cby_1__1__25_chany_bottom_out[10] ,
    \cby_1__1__25_chany_bottom_out[11] ,
    \cby_1__1__25_chany_bottom_out[12] ,
    \cby_1__1__25_chany_bottom_out[13] ,
    \cby_1__1__25_chany_bottom_out[14] ,
    \cby_1__1__25_chany_bottom_out[15] ,
    \cby_1__1__25_chany_bottom_out[16] ,
    \cby_1__1__25_chany_bottom_out[17] ,
    \cby_1__1__25_chany_bottom_out[18] ,
    \cby_1__1__25_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__22_chany_bottom_out[0] ,
    \sb_1__1__22_chany_bottom_out[1] ,
    \sb_1__1__22_chany_bottom_out[2] ,
    \sb_1__1__22_chany_bottom_out[3] ,
    \sb_1__1__22_chany_bottom_out[4] ,
    \sb_1__1__22_chany_bottom_out[5] ,
    \sb_1__1__22_chany_bottom_out[6] ,
    \sb_1__1__22_chany_bottom_out[7] ,
    \sb_1__1__22_chany_bottom_out[8] ,
    \sb_1__1__22_chany_bottom_out[9] ,
    \sb_1__1__22_chany_bottom_out[10] ,
    \sb_1__1__22_chany_bottom_out[11] ,
    \sb_1__1__22_chany_bottom_out[12] ,
    \sb_1__1__22_chany_bottom_out[13] ,
    \sb_1__1__22_chany_bottom_out[14] ,
    \sb_1__1__22_chany_bottom_out[15] ,
    \sb_1__1__22_chany_bottom_out[16] ,
    \sb_1__1__22_chany_bottom_out[17] ,
    \sb_1__1__22_chany_bottom_out[18] ,
    \sb_1__1__22_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__25_chany_top_out[0] ,
    \cby_1__1__25_chany_top_out[1] ,
    \cby_1__1__25_chany_top_out[2] ,
    \cby_1__1__25_chany_top_out[3] ,
    \cby_1__1__25_chany_top_out[4] ,
    \cby_1__1__25_chany_top_out[5] ,
    \cby_1__1__25_chany_top_out[6] ,
    \cby_1__1__25_chany_top_out[7] ,
    \cby_1__1__25_chany_top_out[8] ,
    \cby_1__1__25_chany_top_out[9] ,
    \cby_1__1__25_chany_top_out[10] ,
    \cby_1__1__25_chany_top_out[11] ,
    \cby_1__1__25_chany_top_out[12] ,
    \cby_1__1__25_chany_top_out[13] ,
    \cby_1__1__25_chany_top_out[14] ,
    \cby_1__1__25_chany_top_out[15] ,
    \cby_1__1__25_chany_top_out[16] ,
    \cby_1__1__25_chany_top_out[17] ,
    \cby_1__1__25_chany_top_out[18] ,
    \cby_1__1__25_chany_top_out[19] }));
 cby_1__1_ cby_4__3_ (.Test_en_E_in(\Test_enWires[5] ),
    .Test_en_E_out(\Test_enWires[51] ),
    .Test_en_N_out(\Test_enWires[6] ),
    .Test_en_S_in(\Test_enWires[5] ),
    .Test_en_W_in(\Test_enWires[5] ),
    .Test_en_W_out(\Test_enWires[49] ),
    .ccff_head(grid_clb_26_ccff_tail),
    .ccff_tail(cby_1__1__26_ccff_tail),
    .clk_3_N_out(\clk_3_wires[31] ),
    .clk_3_S_in(\clk_3_wires[32] ),
    .left_grid_pin_16_(cby_1__1__26_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__26_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__26_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__26_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__26_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__26_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__26_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__26_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__26_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__26_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__26_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__26_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__26_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__26_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__26_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__26_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[103] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[102] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[31] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[32] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__22_chany_top_out[0] ,
    \sb_1__1__22_chany_top_out[1] ,
    \sb_1__1__22_chany_top_out[2] ,
    \sb_1__1__22_chany_top_out[3] ,
    \sb_1__1__22_chany_top_out[4] ,
    \sb_1__1__22_chany_top_out[5] ,
    \sb_1__1__22_chany_top_out[6] ,
    \sb_1__1__22_chany_top_out[7] ,
    \sb_1__1__22_chany_top_out[8] ,
    \sb_1__1__22_chany_top_out[9] ,
    \sb_1__1__22_chany_top_out[10] ,
    \sb_1__1__22_chany_top_out[11] ,
    \sb_1__1__22_chany_top_out[12] ,
    \sb_1__1__22_chany_top_out[13] ,
    \sb_1__1__22_chany_top_out[14] ,
    \sb_1__1__22_chany_top_out[15] ,
    \sb_1__1__22_chany_top_out[16] ,
    \sb_1__1__22_chany_top_out[17] ,
    \sb_1__1__22_chany_top_out[18] ,
    \sb_1__1__22_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__26_chany_bottom_out[0] ,
    \cby_1__1__26_chany_bottom_out[1] ,
    \cby_1__1__26_chany_bottom_out[2] ,
    \cby_1__1__26_chany_bottom_out[3] ,
    \cby_1__1__26_chany_bottom_out[4] ,
    \cby_1__1__26_chany_bottom_out[5] ,
    \cby_1__1__26_chany_bottom_out[6] ,
    \cby_1__1__26_chany_bottom_out[7] ,
    \cby_1__1__26_chany_bottom_out[8] ,
    \cby_1__1__26_chany_bottom_out[9] ,
    \cby_1__1__26_chany_bottom_out[10] ,
    \cby_1__1__26_chany_bottom_out[11] ,
    \cby_1__1__26_chany_bottom_out[12] ,
    \cby_1__1__26_chany_bottom_out[13] ,
    \cby_1__1__26_chany_bottom_out[14] ,
    \cby_1__1__26_chany_bottom_out[15] ,
    \cby_1__1__26_chany_bottom_out[16] ,
    \cby_1__1__26_chany_bottom_out[17] ,
    \cby_1__1__26_chany_bottom_out[18] ,
    \cby_1__1__26_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__23_chany_bottom_out[0] ,
    \sb_1__1__23_chany_bottom_out[1] ,
    \sb_1__1__23_chany_bottom_out[2] ,
    \sb_1__1__23_chany_bottom_out[3] ,
    \sb_1__1__23_chany_bottom_out[4] ,
    \sb_1__1__23_chany_bottom_out[5] ,
    \sb_1__1__23_chany_bottom_out[6] ,
    \sb_1__1__23_chany_bottom_out[7] ,
    \sb_1__1__23_chany_bottom_out[8] ,
    \sb_1__1__23_chany_bottom_out[9] ,
    \sb_1__1__23_chany_bottom_out[10] ,
    \sb_1__1__23_chany_bottom_out[11] ,
    \sb_1__1__23_chany_bottom_out[12] ,
    \sb_1__1__23_chany_bottom_out[13] ,
    \sb_1__1__23_chany_bottom_out[14] ,
    \sb_1__1__23_chany_bottom_out[15] ,
    \sb_1__1__23_chany_bottom_out[16] ,
    \sb_1__1__23_chany_bottom_out[17] ,
    \sb_1__1__23_chany_bottom_out[18] ,
    \sb_1__1__23_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__26_chany_top_out[0] ,
    \cby_1__1__26_chany_top_out[1] ,
    \cby_1__1__26_chany_top_out[2] ,
    \cby_1__1__26_chany_top_out[3] ,
    \cby_1__1__26_chany_top_out[4] ,
    \cby_1__1__26_chany_top_out[5] ,
    \cby_1__1__26_chany_top_out[6] ,
    \cby_1__1__26_chany_top_out[7] ,
    \cby_1__1__26_chany_top_out[8] ,
    \cby_1__1__26_chany_top_out[9] ,
    \cby_1__1__26_chany_top_out[10] ,
    \cby_1__1__26_chany_top_out[11] ,
    \cby_1__1__26_chany_top_out[12] ,
    \cby_1__1__26_chany_top_out[13] ,
    \cby_1__1__26_chany_top_out[14] ,
    \cby_1__1__26_chany_top_out[15] ,
    \cby_1__1__26_chany_top_out[16] ,
    \cby_1__1__26_chany_top_out[17] ,
    \cby_1__1__26_chany_top_out[18] ,
    \cby_1__1__26_chany_top_out[19] }));
 cby_1__1_ cby_4__4_ (.Test_en_E_in(\Test_enWires[7] ),
    .Test_en_E_out(\Test_enWires[65] ),
    .Test_en_N_out(\Test_enWires[8] ),
    .Test_en_S_in(\Test_enWires[7] ),
    .Test_en_W_in(\Test_enWires[7] ),
    .Test_en_W_out(\Test_enWires[63] ),
    .ccff_head(grid_clb_27_ccff_tail),
    .ccff_tail(cby_1__1__27_ccff_tail),
    .clk_3_N_out(\clk_3_wires[33] ),
    .clk_3_S_in(\clk_3_wires[34] ),
    .left_grid_pin_16_(cby_1__1__27_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__27_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__27_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__27_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__27_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__27_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__27_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__27_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__27_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__27_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__27_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__27_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__27_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__27_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__27_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__27_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[106] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[105] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[33] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[34] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__23_chany_top_out[0] ,
    \sb_1__1__23_chany_top_out[1] ,
    \sb_1__1__23_chany_top_out[2] ,
    \sb_1__1__23_chany_top_out[3] ,
    \sb_1__1__23_chany_top_out[4] ,
    \sb_1__1__23_chany_top_out[5] ,
    \sb_1__1__23_chany_top_out[6] ,
    \sb_1__1__23_chany_top_out[7] ,
    \sb_1__1__23_chany_top_out[8] ,
    \sb_1__1__23_chany_top_out[9] ,
    \sb_1__1__23_chany_top_out[10] ,
    \sb_1__1__23_chany_top_out[11] ,
    \sb_1__1__23_chany_top_out[12] ,
    \sb_1__1__23_chany_top_out[13] ,
    \sb_1__1__23_chany_top_out[14] ,
    \sb_1__1__23_chany_top_out[15] ,
    \sb_1__1__23_chany_top_out[16] ,
    \sb_1__1__23_chany_top_out[17] ,
    \sb_1__1__23_chany_top_out[18] ,
    \sb_1__1__23_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__27_chany_bottom_out[0] ,
    \cby_1__1__27_chany_bottom_out[1] ,
    \cby_1__1__27_chany_bottom_out[2] ,
    \cby_1__1__27_chany_bottom_out[3] ,
    \cby_1__1__27_chany_bottom_out[4] ,
    \cby_1__1__27_chany_bottom_out[5] ,
    \cby_1__1__27_chany_bottom_out[6] ,
    \cby_1__1__27_chany_bottom_out[7] ,
    \cby_1__1__27_chany_bottom_out[8] ,
    \cby_1__1__27_chany_bottom_out[9] ,
    \cby_1__1__27_chany_bottom_out[10] ,
    \cby_1__1__27_chany_bottom_out[11] ,
    \cby_1__1__27_chany_bottom_out[12] ,
    \cby_1__1__27_chany_bottom_out[13] ,
    \cby_1__1__27_chany_bottom_out[14] ,
    \cby_1__1__27_chany_bottom_out[15] ,
    \cby_1__1__27_chany_bottom_out[16] ,
    \cby_1__1__27_chany_bottom_out[17] ,
    \cby_1__1__27_chany_bottom_out[18] ,
    \cby_1__1__27_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__24_chany_bottom_out[0] ,
    \sb_1__1__24_chany_bottom_out[1] ,
    \sb_1__1__24_chany_bottom_out[2] ,
    \sb_1__1__24_chany_bottom_out[3] ,
    \sb_1__1__24_chany_bottom_out[4] ,
    \sb_1__1__24_chany_bottom_out[5] ,
    \sb_1__1__24_chany_bottom_out[6] ,
    \sb_1__1__24_chany_bottom_out[7] ,
    \sb_1__1__24_chany_bottom_out[8] ,
    \sb_1__1__24_chany_bottom_out[9] ,
    \sb_1__1__24_chany_bottom_out[10] ,
    \sb_1__1__24_chany_bottom_out[11] ,
    \sb_1__1__24_chany_bottom_out[12] ,
    \sb_1__1__24_chany_bottom_out[13] ,
    \sb_1__1__24_chany_bottom_out[14] ,
    \sb_1__1__24_chany_bottom_out[15] ,
    \sb_1__1__24_chany_bottom_out[16] ,
    \sb_1__1__24_chany_bottom_out[17] ,
    \sb_1__1__24_chany_bottom_out[18] ,
    \sb_1__1__24_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__27_chany_top_out[0] ,
    \cby_1__1__27_chany_top_out[1] ,
    \cby_1__1__27_chany_top_out[2] ,
    \cby_1__1__27_chany_top_out[3] ,
    \cby_1__1__27_chany_top_out[4] ,
    \cby_1__1__27_chany_top_out[5] ,
    \cby_1__1__27_chany_top_out[6] ,
    \cby_1__1__27_chany_top_out[7] ,
    \cby_1__1__27_chany_top_out[8] ,
    \cby_1__1__27_chany_top_out[9] ,
    \cby_1__1__27_chany_top_out[10] ,
    \cby_1__1__27_chany_top_out[11] ,
    \cby_1__1__27_chany_top_out[12] ,
    \cby_1__1__27_chany_top_out[13] ,
    \cby_1__1__27_chany_top_out[14] ,
    \cby_1__1__27_chany_top_out[15] ,
    \cby_1__1__27_chany_top_out[16] ,
    \cby_1__1__27_chany_top_out[17] ,
    \cby_1__1__27_chany_top_out[18] ,
    \cby_1__1__27_chany_top_out[19] }));
 cby_1__1_ cby_4__5_ (.Test_en_E_in(\Test_enWires[9] ),
    .Test_en_E_out(\Test_enWires[79] ),
    .Test_en_N_out(\Test_enWires[10] ),
    .Test_en_S_in(\Test_enWires[9] ),
    .Test_en_W_in(\Test_enWires[9] ),
    .Test_en_W_out(\Test_enWires[77] ),
    .ccff_head(grid_clb_28_ccff_tail),
    .ccff_tail(cby_1__1__28_ccff_tail),
    .left_grid_pin_16_(cby_1__1__28_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__28_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__28_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__28_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__28_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__28_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__28_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__28_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__28_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__28_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__28_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__28_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__28_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__28_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__28_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__28_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[109] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[108] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__24_chany_top_out[0] ,
    \sb_1__1__24_chany_top_out[1] ,
    \sb_1__1__24_chany_top_out[2] ,
    \sb_1__1__24_chany_top_out[3] ,
    \sb_1__1__24_chany_top_out[4] ,
    \sb_1__1__24_chany_top_out[5] ,
    \sb_1__1__24_chany_top_out[6] ,
    \sb_1__1__24_chany_top_out[7] ,
    \sb_1__1__24_chany_top_out[8] ,
    \sb_1__1__24_chany_top_out[9] ,
    \sb_1__1__24_chany_top_out[10] ,
    \sb_1__1__24_chany_top_out[11] ,
    \sb_1__1__24_chany_top_out[12] ,
    \sb_1__1__24_chany_top_out[13] ,
    \sb_1__1__24_chany_top_out[14] ,
    \sb_1__1__24_chany_top_out[15] ,
    \sb_1__1__24_chany_top_out[16] ,
    \sb_1__1__24_chany_top_out[17] ,
    \sb_1__1__24_chany_top_out[18] ,
    \sb_1__1__24_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__28_chany_bottom_out[0] ,
    \cby_1__1__28_chany_bottom_out[1] ,
    \cby_1__1__28_chany_bottom_out[2] ,
    \cby_1__1__28_chany_bottom_out[3] ,
    \cby_1__1__28_chany_bottom_out[4] ,
    \cby_1__1__28_chany_bottom_out[5] ,
    \cby_1__1__28_chany_bottom_out[6] ,
    \cby_1__1__28_chany_bottom_out[7] ,
    \cby_1__1__28_chany_bottom_out[8] ,
    \cby_1__1__28_chany_bottom_out[9] ,
    \cby_1__1__28_chany_bottom_out[10] ,
    \cby_1__1__28_chany_bottom_out[11] ,
    \cby_1__1__28_chany_bottom_out[12] ,
    \cby_1__1__28_chany_bottom_out[13] ,
    \cby_1__1__28_chany_bottom_out[14] ,
    \cby_1__1__28_chany_bottom_out[15] ,
    \cby_1__1__28_chany_bottom_out[16] ,
    \cby_1__1__28_chany_bottom_out[17] ,
    \cby_1__1__28_chany_bottom_out[18] ,
    \cby_1__1__28_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__25_chany_bottom_out[0] ,
    \sb_1__1__25_chany_bottom_out[1] ,
    \sb_1__1__25_chany_bottom_out[2] ,
    \sb_1__1__25_chany_bottom_out[3] ,
    \sb_1__1__25_chany_bottom_out[4] ,
    \sb_1__1__25_chany_bottom_out[5] ,
    \sb_1__1__25_chany_bottom_out[6] ,
    \sb_1__1__25_chany_bottom_out[7] ,
    \sb_1__1__25_chany_bottom_out[8] ,
    \sb_1__1__25_chany_bottom_out[9] ,
    \sb_1__1__25_chany_bottom_out[10] ,
    \sb_1__1__25_chany_bottom_out[11] ,
    \sb_1__1__25_chany_bottom_out[12] ,
    \sb_1__1__25_chany_bottom_out[13] ,
    \sb_1__1__25_chany_bottom_out[14] ,
    \sb_1__1__25_chany_bottom_out[15] ,
    \sb_1__1__25_chany_bottom_out[16] ,
    \sb_1__1__25_chany_bottom_out[17] ,
    \sb_1__1__25_chany_bottom_out[18] ,
    \sb_1__1__25_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__28_chany_top_out[0] ,
    \cby_1__1__28_chany_top_out[1] ,
    \cby_1__1__28_chany_top_out[2] ,
    \cby_1__1__28_chany_top_out[3] ,
    \cby_1__1__28_chany_top_out[4] ,
    \cby_1__1__28_chany_top_out[5] ,
    \cby_1__1__28_chany_top_out[6] ,
    \cby_1__1__28_chany_top_out[7] ,
    \cby_1__1__28_chany_top_out[8] ,
    \cby_1__1__28_chany_top_out[9] ,
    \cby_1__1__28_chany_top_out[10] ,
    \cby_1__1__28_chany_top_out[11] ,
    \cby_1__1__28_chany_top_out[12] ,
    \cby_1__1__28_chany_top_out[13] ,
    \cby_1__1__28_chany_top_out[14] ,
    \cby_1__1__28_chany_top_out[15] ,
    \cby_1__1__28_chany_top_out[16] ,
    \cby_1__1__28_chany_top_out[17] ,
    \cby_1__1__28_chany_top_out[18] ,
    \cby_1__1__28_chany_top_out[19] }));
 cby_1__1_ cby_4__6_ (.Test_en_E_in(\Test_enWires[11] ),
    .Test_en_E_out(\Test_enWires[93] ),
    .Test_en_N_out(\Test_enWires[12] ),
    .Test_en_S_in(\Test_enWires[11] ),
    .Test_en_W_in(\Test_enWires[11] ),
    .Test_en_W_out(\Test_enWires[91] ),
    .ccff_head(grid_clb_29_ccff_tail),
    .ccff_tail(cby_1__1__29_ccff_tail),
    .left_grid_pin_16_(cby_1__1__29_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__29_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__29_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__29_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__29_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__29_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__29_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__29_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__29_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__29_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__29_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__29_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__29_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__29_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__29_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__29_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[112] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[111] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__25_chany_top_out[0] ,
    \sb_1__1__25_chany_top_out[1] ,
    \sb_1__1__25_chany_top_out[2] ,
    \sb_1__1__25_chany_top_out[3] ,
    \sb_1__1__25_chany_top_out[4] ,
    \sb_1__1__25_chany_top_out[5] ,
    \sb_1__1__25_chany_top_out[6] ,
    \sb_1__1__25_chany_top_out[7] ,
    \sb_1__1__25_chany_top_out[8] ,
    \sb_1__1__25_chany_top_out[9] ,
    \sb_1__1__25_chany_top_out[10] ,
    \sb_1__1__25_chany_top_out[11] ,
    \sb_1__1__25_chany_top_out[12] ,
    \sb_1__1__25_chany_top_out[13] ,
    \sb_1__1__25_chany_top_out[14] ,
    \sb_1__1__25_chany_top_out[15] ,
    \sb_1__1__25_chany_top_out[16] ,
    \sb_1__1__25_chany_top_out[17] ,
    \sb_1__1__25_chany_top_out[18] ,
    \sb_1__1__25_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__29_chany_bottom_out[0] ,
    \cby_1__1__29_chany_bottom_out[1] ,
    \cby_1__1__29_chany_bottom_out[2] ,
    \cby_1__1__29_chany_bottom_out[3] ,
    \cby_1__1__29_chany_bottom_out[4] ,
    \cby_1__1__29_chany_bottom_out[5] ,
    \cby_1__1__29_chany_bottom_out[6] ,
    \cby_1__1__29_chany_bottom_out[7] ,
    \cby_1__1__29_chany_bottom_out[8] ,
    \cby_1__1__29_chany_bottom_out[9] ,
    \cby_1__1__29_chany_bottom_out[10] ,
    \cby_1__1__29_chany_bottom_out[11] ,
    \cby_1__1__29_chany_bottom_out[12] ,
    \cby_1__1__29_chany_bottom_out[13] ,
    \cby_1__1__29_chany_bottom_out[14] ,
    \cby_1__1__29_chany_bottom_out[15] ,
    \cby_1__1__29_chany_bottom_out[16] ,
    \cby_1__1__29_chany_bottom_out[17] ,
    \cby_1__1__29_chany_bottom_out[18] ,
    \cby_1__1__29_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__26_chany_bottom_out[0] ,
    \sb_1__1__26_chany_bottom_out[1] ,
    \sb_1__1__26_chany_bottom_out[2] ,
    \sb_1__1__26_chany_bottom_out[3] ,
    \sb_1__1__26_chany_bottom_out[4] ,
    \sb_1__1__26_chany_bottom_out[5] ,
    \sb_1__1__26_chany_bottom_out[6] ,
    \sb_1__1__26_chany_bottom_out[7] ,
    \sb_1__1__26_chany_bottom_out[8] ,
    \sb_1__1__26_chany_bottom_out[9] ,
    \sb_1__1__26_chany_bottom_out[10] ,
    \sb_1__1__26_chany_bottom_out[11] ,
    \sb_1__1__26_chany_bottom_out[12] ,
    \sb_1__1__26_chany_bottom_out[13] ,
    \sb_1__1__26_chany_bottom_out[14] ,
    \sb_1__1__26_chany_bottom_out[15] ,
    \sb_1__1__26_chany_bottom_out[16] ,
    \sb_1__1__26_chany_bottom_out[17] ,
    \sb_1__1__26_chany_bottom_out[18] ,
    \sb_1__1__26_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__29_chany_top_out[0] ,
    \cby_1__1__29_chany_top_out[1] ,
    \cby_1__1__29_chany_top_out[2] ,
    \cby_1__1__29_chany_top_out[3] ,
    \cby_1__1__29_chany_top_out[4] ,
    \cby_1__1__29_chany_top_out[5] ,
    \cby_1__1__29_chany_top_out[6] ,
    \cby_1__1__29_chany_top_out[7] ,
    \cby_1__1__29_chany_top_out[8] ,
    \cby_1__1__29_chany_top_out[9] ,
    \cby_1__1__29_chany_top_out[10] ,
    \cby_1__1__29_chany_top_out[11] ,
    \cby_1__1__29_chany_top_out[12] ,
    \cby_1__1__29_chany_top_out[13] ,
    \cby_1__1__29_chany_top_out[14] ,
    \cby_1__1__29_chany_top_out[15] ,
    \cby_1__1__29_chany_top_out[16] ,
    \cby_1__1__29_chany_top_out[17] ,
    \cby_1__1__29_chany_top_out[18] ,
    \cby_1__1__29_chany_top_out[19] }));
 cby_1__1_ cby_4__7_ (.Test_en_E_in(\Test_enWires[13] ),
    .Test_en_E_out(\Test_enWires[107] ),
    .Test_en_N_out(\Test_enWires[14] ),
    .Test_en_S_in(\Test_enWires[13] ),
    .Test_en_W_in(\Test_enWires[13] ),
    .Test_en_W_out(\Test_enWires[105] ),
    .ccff_head(grid_clb_30_ccff_tail),
    .ccff_tail(cby_1__1__30_ccff_tail),
    .left_grid_pin_16_(cby_1__1__30_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__30_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__30_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__30_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__30_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__30_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__30_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__30_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__30_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__30_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__30_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__30_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__30_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__30_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__30_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__30_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[115] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[114] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__26_chany_top_out[0] ,
    \sb_1__1__26_chany_top_out[1] ,
    \sb_1__1__26_chany_top_out[2] ,
    \sb_1__1__26_chany_top_out[3] ,
    \sb_1__1__26_chany_top_out[4] ,
    \sb_1__1__26_chany_top_out[5] ,
    \sb_1__1__26_chany_top_out[6] ,
    \sb_1__1__26_chany_top_out[7] ,
    \sb_1__1__26_chany_top_out[8] ,
    \sb_1__1__26_chany_top_out[9] ,
    \sb_1__1__26_chany_top_out[10] ,
    \sb_1__1__26_chany_top_out[11] ,
    \sb_1__1__26_chany_top_out[12] ,
    \sb_1__1__26_chany_top_out[13] ,
    \sb_1__1__26_chany_top_out[14] ,
    \sb_1__1__26_chany_top_out[15] ,
    \sb_1__1__26_chany_top_out[16] ,
    \sb_1__1__26_chany_top_out[17] ,
    \sb_1__1__26_chany_top_out[18] ,
    \sb_1__1__26_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__30_chany_bottom_out[0] ,
    \cby_1__1__30_chany_bottom_out[1] ,
    \cby_1__1__30_chany_bottom_out[2] ,
    \cby_1__1__30_chany_bottom_out[3] ,
    \cby_1__1__30_chany_bottom_out[4] ,
    \cby_1__1__30_chany_bottom_out[5] ,
    \cby_1__1__30_chany_bottom_out[6] ,
    \cby_1__1__30_chany_bottom_out[7] ,
    \cby_1__1__30_chany_bottom_out[8] ,
    \cby_1__1__30_chany_bottom_out[9] ,
    \cby_1__1__30_chany_bottom_out[10] ,
    \cby_1__1__30_chany_bottom_out[11] ,
    \cby_1__1__30_chany_bottom_out[12] ,
    \cby_1__1__30_chany_bottom_out[13] ,
    \cby_1__1__30_chany_bottom_out[14] ,
    \cby_1__1__30_chany_bottom_out[15] ,
    \cby_1__1__30_chany_bottom_out[16] ,
    \cby_1__1__30_chany_bottom_out[17] ,
    \cby_1__1__30_chany_bottom_out[18] ,
    \cby_1__1__30_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__27_chany_bottom_out[0] ,
    \sb_1__1__27_chany_bottom_out[1] ,
    \sb_1__1__27_chany_bottom_out[2] ,
    \sb_1__1__27_chany_bottom_out[3] ,
    \sb_1__1__27_chany_bottom_out[4] ,
    \sb_1__1__27_chany_bottom_out[5] ,
    \sb_1__1__27_chany_bottom_out[6] ,
    \sb_1__1__27_chany_bottom_out[7] ,
    \sb_1__1__27_chany_bottom_out[8] ,
    \sb_1__1__27_chany_bottom_out[9] ,
    \sb_1__1__27_chany_bottom_out[10] ,
    \sb_1__1__27_chany_bottom_out[11] ,
    \sb_1__1__27_chany_bottom_out[12] ,
    \sb_1__1__27_chany_bottom_out[13] ,
    \sb_1__1__27_chany_bottom_out[14] ,
    \sb_1__1__27_chany_bottom_out[15] ,
    \sb_1__1__27_chany_bottom_out[16] ,
    \sb_1__1__27_chany_bottom_out[17] ,
    \sb_1__1__27_chany_bottom_out[18] ,
    \sb_1__1__27_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__30_chany_top_out[0] ,
    \cby_1__1__30_chany_top_out[1] ,
    \cby_1__1__30_chany_top_out[2] ,
    \cby_1__1__30_chany_top_out[3] ,
    \cby_1__1__30_chany_top_out[4] ,
    \cby_1__1__30_chany_top_out[5] ,
    \cby_1__1__30_chany_top_out[6] ,
    \cby_1__1__30_chany_top_out[7] ,
    \cby_1__1__30_chany_top_out[8] ,
    \cby_1__1__30_chany_top_out[9] ,
    \cby_1__1__30_chany_top_out[10] ,
    \cby_1__1__30_chany_top_out[11] ,
    \cby_1__1__30_chany_top_out[12] ,
    \cby_1__1__30_chany_top_out[13] ,
    \cby_1__1__30_chany_top_out[14] ,
    \cby_1__1__30_chany_top_out[15] ,
    \cby_1__1__30_chany_top_out[16] ,
    \cby_1__1__30_chany_top_out[17] ,
    \cby_1__1__30_chany_top_out[18] ,
    \cby_1__1__30_chany_top_out[19] }));
 cby_1__1_ cby_4__8_ (.Test_en_E_in(\Test_enWires[15] ),
    .Test_en_E_out(\Test_enWires[121] ),
    .Test_en_S_in(\Test_enWires[15] ),
    .Test_en_W_in(\Test_enWires[15] ),
    .Test_en_W_out(\Test_enWires[119] ),
    .ccff_head(grid_clb_31_ccff_tail),
    .ccff_tail(cby_1__1__31_ccff_tail),
    .left_grid_pin_16_(cby_1__1__31_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__31_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__31_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__31_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__31_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__31_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__31_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__31_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__31_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__31_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__31_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__31_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__31_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__31_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__31_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__31_left_grid_pin_31_),
    .prog_clk_0_N_out(\prog_clk_0_wires[120] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[118] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[117] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__27_chany_top_out[0] ,
    \sb_1__1__27_chany_top_out[1] ,
    \sb_1__1__27_chany_top_out[2] ,
    \sb_1__1__27_chany_top_out[3] ,
    \sb_1__1__27_chany_top_out[4] ,
    \sb_1__1__27_chany_top_out[5] ,
    \sb_1__1__27_chany_top_out[6] ,
    \sb_1__1__27_chany_top_out[7] ,
    \sb_1__1__27_chany_top_out[8] ,
    \sb_1__1__27_chany_top_out[9] ,
    \sb_1__1__27_chany_top_out[10] ,
    \sb_1__1__27_chany_top_out[11] ,
    \sb_1__1__27_chany_top_out[12] ,
    \sb_1__1__27_chany_top_out[13] ,
    \sb_1__1__27_chany_top_out[14] ,
    \sb_1__1__27_chany_top_out[15] ,
    \sb_1__1__27_chany_top_out[16] ,
    \sb_1__1__27_chany_top_out[17] ,
    \sb_1__1__27_chany_top_out[18] ,
    \sb_1__1__27_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__31_chany_bottom_out[0] ,
    \cby_1__1__31_chany_bottom_out[1] ,
    \cby_1__1__31_chany_bottom_out[2] ,
    \cby_1__1__31_chany_bottom_out[3] ,
    \cby_1__1__31_chany_bottom_out[4] ,
    \cby_1__1__31_chany_bottom_out[5] ,
    \cby_1__1__31_chany_bottom_out[6] ,
    \cby_1__1__31_chany_bottom_out[7] ,
    \cby_1__1__31_chany_bottom_out[8] ,
    \cby_1__1__31_chany_bottom_out[9] ,
    \cby_1__1__31_chany_bottom_out[10] ,
    \cby_1__1__31_chany_bottom_out[11] ,
    \cby_1__1__31_chany_bottom_out[12] ,
    \cby_1__1__31_chany_bottom_out[13] ,
    \cby_1__1__31_chany_bottom_out[14] ,
    \cby_1__1__31_chany_bottom_out[15] ,
    \cby_1__1__31_chany_bottom_out[16] ,
    \cby_1__1__31_chany_bottom_out[17] ,
    \cby_1__1__31_chany_bottom_out[18] ,
    \cby_1__1__31_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__8__3_chany_bottom_out[0] ,
    \sb_1__8__3_chany_bottom_out[1] ,
    \sb_1__8__3_chany_bottom_out[2] ,
    \sb_1__8__3_chany_bottom_out[3] ,
    \sb_1__8__3_chany_bottom_out[4] ,
    \sb_1__8__3_chany_bottom_out[5] ,
    \sb_1__8__3_chany_bottom_out[6] ,
    \sb_1__8__3_chany_bottom_out[7] ,
    \sb_1__8__3_chany_bottom_out[8] ,
    \sb_1__8__3_chany_bottom_out[9] ,
    \sb_1__8__3_chany_bottom_out[10] ,
    \sb_1__8__3_chany_bottom_out[11] ,
    \sb_1__8__3_chany_bottom_out[12] ,
    \sb_1__8__3_chany_bottom_out[13] ,
    \sb_1__8__3_chany_bottom_out[14] ,
    \sb_1__8__3_chany_bottom_out[15] ,
    \sb_1__8__3_chany_bottom_out[16] ,
    \sb_1__8__3_chany_bottom_out[17] ,
    \sb_1__8__3_chany_bottom_out[18] ,
    \sb_1__8__3_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__31_chany_top_out[0] ,
    \cby_1__1__31_chany_top_out[1] ,
    \cby_1__1__31_chany_top_out[2] ,
    \cby_1__1__31_chany_top_out[3] ,
    \cby_1__1__31_chany_top_out[4] ,
    \cby_1__1__31_chany_top_out[5] ,
    \cby_1__1__31_chany_top_out[6] ,
    \cby_1__1__31_chany_top_out[7] ,
    \cby_1__1__31_chany_top_out[8] ,
    \cby_1__1__31_chany_top_out[9] ,
    \cby_1__1__31_chany_top_out[10] ,
    \cby_1__1__31_chany_top_out[11] ,
    \cby_1__1__31_chany_top_out[12] ,
    \cby_1__1__31_chany_top_out[13] ,
    \cby_1__1__31_chany_top_out[14] ,
    \cby_1__1__31_chany_top_out[15] ,
    \cby_1__1__31_chany_top_out[16] ,
    \cby_1__1__31_chany_top_out[17] ,
    \cby_1__1__31_chany_top_out[18] ,
    \cby_1__1__31_chany_top_out[19] }));
 cby_1__1_ cby_5__1_ (.Test_en_E_in(\Test_enWires[24] ),
    .Test_en_E_out(\Test_enWires[25] ),
    .Test_en_S_in(\Test_enWires[24] ),
    .Test_en_W_in(\Test_enWires[24] ),
    .ccff_head(grid_clb_32_ccff_tail),
    .ccff_tail(cby_1__1__32_ccff_tail),
    .left_grid_pin_16_(cby_1__1__32_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__32_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__32_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__32_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__32_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__32_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__32_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__32_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__32_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__32_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__32_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__32_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__32_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__32_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__32_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__32_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[123] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[122] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__0__4_chany_top_out[0] ,
    \sb_1__0__4_chany_top_out[1] ,
    \sb_1__0__4_chany_top_out[2] ,
    \sb_1__0__4_chany_top_out[3] ,
    \sb_1__0__4_chany_top_out[4] ,
    \sb_1__0__4_chany_top_out[5] ,
    \sb_1__0__4_chany_top_out[6] ,
    \sb_1__0__4_chany_top_out[7] ,
    \sb_1__0__4_chany_top_out[8] ,
    \sb_1__0__4_chany_top_out[9] ,
    \sb_1__0__4_chany_top_out[10] ,
    \sb_1__0__4_chany_top_out[11] ,
    \sb_1__0__4_chany_top_out[12] ,
    \sb_1__0__4_chany_top_out[13] ,
    \sb_1__0__4_chany_top_out[14] ,
    \sb_1__0__4_chany_top_out[15] ,
    \sb_1__0__4_chany_top_out[16] ,
    \sb_1__0__4_chany_top_out[17] ,
    \sb_1__0__4_chany_top_out[18] ,
    \sb_1__0__4_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__32_chany_bottom_out[0] ,
    \cby_1__1__32_chany_bottom_out[1] ,
    \cby_1__1__32_chany_bottom_out[2] ,
    \cby_1__1__32_chany_bottom_out[3] ,
    \cby_1__1__32_chany_bottom_out[4] ,
    \cby_1__1__32_chany_bottom_out[5] ,
    \cby_1__1__32_chany_bottom_out[6] ,
    \cby_1__1__32_chany_bottom_out[7] ,
    \cby_1__1__32_chany_bottom_out[8] ,
    \cby_1__1__32_chany_bottom_out[9] ,
    \cby_1__1__32_chany_bottom_out[10] ,
    \cby_1__1__32_chany_bottom_out[11] ,
    \cby_1__1__32_chany_bottom_out[12] ,
    \cby_1__1__32_chany_bottom_out[13] ,
    \cby_1__1__32_chany_bottom_out[14] ,
    \cby_1__1__32_chany_bottom_out[15] ,
    \cby_1__1__32_chany_bottom_out[16] ,
    \cby_1__1__32_chany_bottom_out[17] ,
    \cby_1__1__32_chany_bottom_out[18] ,
    \cby_1__1__32_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__28_chany_bottom_out[0] ,
    \sb_1__1__28_chany_bottom_out[1] ,
    \sb_1__1__28_chany_bottom_out[2] ,
    \sb_1__1__28_chany_bottom_out[3] ,
    \sb_1__1__28_chany_bottom_out[4] ,
    \sb_1__1__28_chany_bottom_out[5] ,
    \sb_1__1__28_chany_bottom_out[6] ,
    \sb_1__1__28_chany_bottom_out[7] ,
    \sb_1__1__28_chany_bottom_out[8] ,
    \sb_1__1__28_chany_bottom_out[9] ,
    \sb_1__1__28_chany_bottom_out[10] ,
    \sb_1__1__28_chany_bottom_out[11] ,
    \sb_1__1__28_chany_bottom_out[12] ,
    \sb_1__1__28_chany_bottom_out[13] ,
    \sb_1__1__28_chany_bottom_out[14] ,
    \sb_1__1__28_chany_bottom_out[15] ,
    \sb_1__1__28_chany_bottom_out[16] ,
    \sb_1__1__28_chany_bottom_out[17] ,
    \sb_1__1__28_chany_bottom_out[18] ,
    \sb_1__1__28_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__32_chany_top_out[0] ,
    \cby_1__1__32_chany_top_out[1] ,
    \cby_1__1__32_chany_top_out[2] ,
    \cby_1__1__32_chany_top_out[3] ,
    \cby_1__1__32_chany_top_out[4] ,
    \cby_1__1__32_chany_top_out[5] ,
    \cby_1__1__32_chany_top_out[6] ,
    \cby_1__1__32_chany_top_out[7] ,
    \cby_1__1__32_chany_top_out[8] ,
    \cby_1__1__32_chany_top_out[9] ,
    \cby_1__1__32_chany_top_out[10] ,
    \cby_1__1__32_chany_top_out[11] ,
    \cby_1__1__32_chany_top_out[12] ,
    \cby_1__1__32_chany_top_out[13] ,
    \cby_1__1__32_chany_top_out[14] ,
    \cby_1__1__32_chany_top_out[15] ,
    \cby_1__1__32_chany_top_out[16] ,
    \cby_1__1__32_chany_top_out[17] ,
    \cby_1__1__32_chany_top_out[18] ,
    \cby_1__1__32_chany_top_out[19] }));
 cby_1__1_ cby_5__2_ (.Test_en_E_in(\Test_enWires[38] ),
    .Test_en_E_out(\Test_enWires[39] ),
    .Test_en_S_in(\Test_enWires[38] ),
    .Test_en_W_in(\Test_enWires[38] ),
    .ccff_head(grid_clb_33_ccff_tail),
    .ccff_tail(cby_1__1__33_ccff_tail),
    .clk_2_S_in(\clk_2_wires[33] ),
    .clk_2_S_out(\clk_2_wires[34] ),
    .left_grid_pin_16_(cby_1__1__33_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__33_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__33_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__33_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__33_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__33_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__33_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__33_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__33_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__33_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__33_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__33_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__33_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__33_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__33_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__33_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[126] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[125] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[33] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[34] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__28_chany_top_out[0] ,
    \sb_1__1__28_chany_top_out[1] ,
    \sb_1__1__28_chany_top_out[2] ,
    \sb_1__1__28_chany_top_out[3] ,
    \sb_1__1__28_chany_top_out[4] ,
    \sb_1__1__28_chany_top_out[5] ,
    \sb_1__1__28_chany_top_out[6] ,
    \sb_1__1__28_chany_top_out[7] ,
    \sb_1__1__28_chany_top_out[8] ,
    \sb_1__1__28_chany_top_out[9] ,
    \sb_1__1__28_chany_top_out[10] ,
    \sb_1__1__28_chany_top_out[11] ,
    \sb_1__1__28_chany_top_out[12] ,
    \sb_1__1__28_chany_top_out[13] ,
    \sb_1__1__28_chany_top_out[14] ,
    \sb_1__1__28_chany_top_out[15] ,
    \sb_1__1__28_chany_top_out[16] ,
    \sb_1__1__28_chany_top_out[17] ,
    \sb_1__1__28_chany_top_out[18] ,
    \sb_1__1__28_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__33_chany_bottom_out[0] ,
    \cby_1__1__33_chany_bottom_out[1] ,
    \cby_1__1__33_chany_bottom_out[2] ,
    \cby_1__1__33_chany_bottom_out[3] ,
    \cby_1__1__33_chany_bottom_out[4] ,
    \cby_1__1__33_chany_bottom_out[5] ,
    \cby_1__1__33_chany_bottom_out[6] ,
    \cby_1__1__33_chany_bottom_out[7] ,
    \cby_1__1__33_chany_bottom_out[8] ,
    \cby_1__1__33_chany_bottom_out[9] ,
    \cby_1__1__33_chany_bottom_out[10] ,
    \cby_1__1__33_chany_bottom_out[11] ,
    \cby_1__1__33_chany_bottom_out[12] ,
    \cby_1__1__33_chany_bottom_out[13] ,
    \cby_1__1__33_chany_bottom_out[14] ,
    \cby_1__1__33_chany_bottom_out[15] ,
    \cby_1__1__33_chany_bottom_out[16] ,
    \cby_1__1__33_chany_bottom_out[17] ,
    \cby_1__1__33_chany_bottom_out[18] ,
    \cby_1__1__33_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__29_chany_bottom_out[0] ,
    \sb_1__1__29_chany_bottom_out[1] ,
    \sb_1__1__29_chany_bottom_out[2] ,
    \sb_1__1__29_chany_bottom_out[3] ,
    \sb_1__1__29_chany_bottom_out[4] ,
    \sb_1__1__29_chany_bottom_out[5] ,
    \sb_1__1__29_chany_bottom_out[6] ,
    \sb_1__1__29_chany_bottom_out[7] ,
    \sb_1__1__29_chany_bottom_out[8] ,
    \sb_1__1__29_chany_bottom_out[9] ,
    \sb_1__1__29_chany_bottom_out[10] ,
    \sb_1__1__29_chany_bottom_out[11] ,
    \sb_1__1__29_chany_bottom_out[12] ,
    \sb_1__1__29_chany_bottom_out[13] ,
    \sb_1__1__29_chany_bottom_out[14] ,
    \sb_1__1__29_chany_bottom_out[15] ,
    \sb_1__1__29_chany_bottom_out[16] ,
    \sb_1__1__29_chany_bottom_out[17] ,
    \sb_1__1__29_chany_bottom_out[18] ,
    \sb_1__1__29_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__33_chany_top_out[0] ,
    \cby_1__1__33_chany_top_out[1] ,
    \cby_1__1__33_chany_top_out[2] ,
    \cby_1__1__33_chany_top_out[3] ,
    \cby_1__1__33_chany_top_out[4] ,
    \cby_1__1__33_chany_top_out[5] ,
    \cby_1__1__33_chany_top_out[6] ,
    \cby_1__1__33_chany_top_out[7] ,
    \cby_1__1__33_chany_top_out[8] ,
    \cby_1__1__33_chany_top_out[9] ,
    \cby_1__1__33_chany_top_out[10] ,
    \cby_1__1__33_chany_top_out[11] ,
    \cby_1__1__33_chany_top_out[12] ,
    \cby_1__1__33_chany_top_out[13] ,
    \cby_1__1__33_chany_top_out[14] ,
    \cby_1__1__33_chany_top_out[15] ,
    \cby_1__1__33_chany_top_out[16] ,
    \cby_1__1__33_chany_top_out[17] ,
    \cby_1__1__33_chany_top_out[18] ,
    \cby_1__1__33_chany_top_out[19] }));
 cby_1__1_ cby_5__3_ (.Test_en_E_in(\Test_enWires[52] ),
    .Test_en_E_out(\Test_enWires[53] ),
    .Test_en_S_in(\Test_enWires[52] ),
    .Test_en_W_in(\Test_enWires[52] ),
    .ccff_head(grid_clb_34_ccff_tail),
    .ccff_tail(cby_1__1__34_ccff_tail),
    .clk_2_N_out(\clk_2_wires[32] ),
    .clk_2_S_in(\clk_2_wires[31] ),
    .left_grid_pin_16_(cby_1__1__34_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__34_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__34_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__34_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__34_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__34_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__34_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__34_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__34_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__34_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__34_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__34_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__34_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__34_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__34_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__34_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[129] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[128] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[32] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[31] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__29_chany_top_out[0] ,
    \sb_1__1__29_chany_top_out[1] ,
    \sb_1__1__29_chany_top_out[2] ,
    \sb_1__1__29_chany_top_out[3] ,
    \sb_1__1__29_chany_top_out[4] ,
    \sb_1__1__29_chany_top_out[5] ,
    \sb_1__1__29_chany_top_out[6] ,
    \sb_1__1__29_chany_top_out[7] ,
    \sb_1__1__29_chany_top_out[8] ,
    \sb_1__1__29_chany_top_out[9] ,
    \sb_1__1__29_chany_top_out[10] ,
    \sb_1__1__29_chany_top_out[11] ,
    \sb_1__1__29_chany_top_out[12] ,
    \sb_1__1__29_chany_top_out[13] ,
    \sb_1__1__29_chany_top_out[14] ,
    \sb_1__1__29_chany_top_out[15] ,
    \sb_1__1__29_chany_top_out[16] ,
    \sb_1__1__29_chany_top_out[17] ,
    \sb_1__1__29_chany_top_out[18] ,
    \sb_1__1__29_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__34_chany_bottom_out[0] ,
    \cby_1__1__34_chany_bottom_out[1] ,
    \cby_1__1__34_chany_bottom_out[2] ,
    \cby_1__1__34_chany_bottom_out[3] ,
    \cby_1__1__34_chany_bottom_out[4] ,
    \cby_1__1__34_chany_bottom_out[5] ,
    \cby_1__1__34_chany_bottom_out[6] ,
    \cby_1__1__34_chany_bottom_out[7] ,
    \cby_1__1__34_chany_bottom_out[8] ,
    \cby_1__1__34_chany_bottom_out[9] ,
    \cby_1__1__34_chany_bottom_out[10] ,
    \cby_1__1__34_chany_bottom_out[11] ,
    \cby_1__1__34_chany_bottom_out[12] ,
    \cby_1__1__34_chany_bottom_out[13] ,
    \cby_1__1__34_chany_bottom_out[14] ,
    \cby_1__1__34_chany_bottom_out[15] ,
    \cby_1__1__34_chany_bottom_out[16] ,
    \cby_1__1__34_chany_bottom_out[17] ,
    \cby_1__1__34_chany_bottom_out[18] ,
    \cby_1__1__34_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__30_chany_bottom_out[0] ,
    \sb_1__1__30_chany_bottom_out[1] ,
    \sb_1__1__30_chany_bottom_out[2] ,
    \sb_1__1__30_chany_bottom_out[3] ,
    \sb_1__1__30_chany_bottom_out[4] ,
    \sb_1__1__30_chany_bottom_out[5] ,
    \sb_1__1__30_chany_bottom_out[6] ,
    \sb_1__1__30_chany_bottom_out[7] ,
    \sb_1__1__30_chany_bottom_out[8] ,
    \sb_1__1__30_chany_bottom_out[9] ,
    \sb_1__1__30_chany_bottom_out[10] ,
    \sb_1__1__30_chany_bottom_out[11] ,
    \sb_1__1__30_chany_bottom_out[12] ,
    \sb_1__1__30_chany_bottom_out[13] ,
    \sb_1__1__30_chany_bottom_out[14] ,
    \sb_1__1__30_chany_bottom_out[15] ,
    \sb_1__1__30_chany_bottom_out[16] ,
    \sb_1__1__30_chany_bottom_out[17] ,
    \sb_1__1__30_chany_bottom_out[18] ,
    \sb_1__1__30_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__34_chany_top_out[0] ,
    \cby_1__1__34_chany_top_out[1] ,
    \cby_1__1__34_chany_top_out[2] ,
    \cby_1__1__34_chany_top_out[3] ,
    \cby_1__1__34_chany_top_out[4] ,
    \cby_1__1__34_chany_top_out[5] ,
    \cby_1__1__34_chany_top_out[6] ,
    \cby_1__1__34_chany_top_out[7] ,
    \cby_1__1__34_chany_top_out[8] ,
    \cby_1__1__34_chany_top_out[9] ,
    \cby_1__1__34_chany_top_out[10] ,
    \cby_1__1__34_chany_top_out[11] ,
    \cby_1__1__34_chany_top_out[12] ,
    \cby_1__1__34_chany_top_out[13] ,
    \cby_1__1__34_chany_top_out[14] ,
    \cby_1__1__34_chany_top_out[15] ,
    \cby_1__1__34_chany_top_out[16] ,
    \cby_1__1__34_chany_top_out[17] ,
    \cby_1__1__34_chany_top_out[18] ,
    \cby_1__1__34_chany_top_out[19] }));
 cby_1__1_ cby_5__4_ (.Test_en_E_in(\Test_enWires[66] ),
    .Test_en_E_out(\Test_enWires[67] ),
    .Test_en_S_in(\Test_enWires[66] ),
    .Test_en_W_in(\Test_enWires[66] ),
    .ccff_head(grid_clb_35_ccff_tail),
    .ccff_tail(cby_1__1__35_ccff_tail),
    .left_grid_pin_16_(cby_1__1__35_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__35_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__35_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__35_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__35_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__35_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__35_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__35_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__35_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__35_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__35_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__35_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__35_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__35_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__35_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__35_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[132] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[131] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__30_chany_top_out[0] ,
    \sb_1__1__30_chany_top_out[1] ,
    \sb_1__1__30_chany_top_out[2] ,
    \sb_1__1__30_chany_top_out[3] ,
    \sb_1__1__30_chany_top_out[4] ,
    \sb_1__1__30_chany_top_out[5] ,
    \sb_1__1__30_chany_top_out[6] ,
    \sb_1__1__30_chany_top_out[7] ,
    \sb_1__1__30_chany_top_out[8] ,
    \sb_1__1__30_chany_top_out[9] ,
    \sb_1__1__30_chany_top_out[10] ,
    \sb_1__1__30_chany_top_out[11] ,
    \sb_1__1__30_chany_top_out[12] ,
    \sb_1__1__30_chany_top_out[13] ,
    \sb_1__1__30_chany_top_out[14] ,
    \sb_1__1__30_chany_top_out[15] ,
    \sb_1__1__30_chany_top_out[16] ,
    \sb_1__1__30_chany_top_out[17] ,
    \sb_1__1__30_chany_top_out[18] ,
    \sb_1__1__30_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__35_chany_bottom_out[0] ,
    \cby_1__1__35_chany_bottom_out[1] ,
    \cby_1__1__35_chany_bottom_out[2] ,
    \cby_1__1__35_chany_bottom_out[3] ,
    \cby_1__1__35_chany_bottom_out[4] ,
    \cby_1__1__35_chany_bottom_out[5] ,
    \cby_1__1__35_chany_bottom_out[6] ,
    \cby_1__1__35_chany_bottom_out[7] ,
    \cby_1__1__35_chany_bottom_out[8] ,
    \cby_1__1__35_chany_bottom_out[9] ,
    \cby_1__1__35_chany_bottom_out[10] ,
    \cby_1__1__35_chany_bottom_out[11] ,
    \cby_1__1__35_chany_bottom_out[12] ,
    \cby_1__1__35_chany_bottom_out[13] ,
    \cby_1__1__35_chany_bottom_out[14] ,
    \cby_1__1__35_chany_bottom_out[15] ,
    \cby_1__1__35_chany_bottom_out[16] ,
    \cby_1__1__35_chany_bottom_out[17] ,
    \cby_1__1__35_chany_bottom_out[18] ,
    \cby_1__1__35_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__31_chany_bottom_out[0] ,
    \sb_1__1__31_chany_bottom_out[1] ,
    \sb_1__1__31_chany_bottom_out[2] ,
    \sb_1__1__31_chany_bottom_out[3] ,
    \sb_1__1__31_chany_bottom_out[4] ,
    \sb_1__1__31_chany_bottom_out[5] ,
    \sb_1__1__31_chany_bottom_out[6] ,
    \sb_1__1__31_chany_bottom_out[7] ,
    \sb_1__1__31_chany_bottom_out[8] ,
    \sb_1__1__31_chany_bottom_out[9] ,
    \sb_1__1__31_chany_bottom_out[10] ,
    \sb_1__1__31_chany_bottom_out[11] ,
    \sb_1__1__31_chany_bottom_out[12] ,
    \sb_1__1__31_chany_bottom_out[13] ,
    \sb_1__1__31_chany_bottom_out[14] ,
    \sb_1__1__31_chany_bottom_out[15] ,
    \sb_1__1__31_chany_bottom_out[16] ,
    \sb_1__1__31_chany_bottom_out[17] ,
    \sb_1__1__31_chany_bottom_out[18] ,
    \sb_1__1__31_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__35_chany_top_out[0] ,
    \cby_1__1__35_chany_top_out[1] ,
    \cby_1__1__35_chany_top_out[2] ,
    \cby_1__1__35_chany_top_out[3] ,
    \cby_1__1__35_chany_top_out[4] ,
    \cby_1__1__35_chany_top_out[5] ,
    \cby_1__1__35_chany_top_out[6] ,
    \cby_1__1__35_chany_top_out[7] ,
    \cby_1__1__35_chany_top_out[8] ,
    \cby_1__1__35_chany_top_out[9] ,
    \cby_1__1__35_chany_top_out[10] ,
    \cby_1__1__35_chany_top_out[11] ,
    \cby_1__1__35_chany_top_out[12] ,
    \cby_1__1__35_chany_top_out[13] ,
    \cby_1__1__35_chany_top_out[14] ,
    \cby_1__1__35_chany_top_out[15] ,
    \cby_1__1__35_chany_top_out[16] ,
    \cby_1__1__35_chany_top_out[17] ,
    \cby_1__1__35_chany_top_out[18] ,
    \cby_1__1__35_chany_top_out[19] }));
 cby_1__1_ cby_5__5_ (.Test_en_E_in(\Test_enWires[80] ),
    .Test_en_E_out(\Test_enWires[81] ),
    .Test_en_S_in(\Test_enWires[80] ),
    .Test_en_W_in(\Test_enWires[80] ),
    .ccff_head(grid_clb_36_ccff_tail),
    .ccff_tail(cby_1__1__36_ccff_tail),
    .left_grid_pin_16_(cby_1__1__36_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__36_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__36_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__36_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__36_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__36_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__36_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__36_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__36_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__36_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__36_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__36_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__36_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__36_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__36_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__36_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[135] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[134] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__31_chany_top_out[0] ,
    \sb_1__1__31_chany_top_out[1] ,
    \sb_1__1__31_chany_top_out[2] ,
    \sb_1__1__31_chany_top_out[3] ,
    \sb_1__1__31_chany_top_out[4] ,
    \sb_1__1__31_chany_top_out[5] ,
    \sb_1__1__31_chany_top_out[6] ,
    \sb_1__1__31_chany_top_out[7] ,
    \sb_1__1__31_chany_top_out[8] ,
    \sb_1__1__31_chany_top_out[9] ,
    \sb_1__1__31_chany_top_out[10] ,
    \sb_1__1__31_chany_top_out[11] ,
    \sb_1__1__31_chany_top_out[12] ,
    \sb_1__1__31_chany_top_out[13] ,
    \sb_1__1__31_chany_top_out[14] ,
    \sb_1__1__31_chany_top_out[15] ,
    \sb_1__1__31_chany_top_out[16] ,
    \sb_1__1__31_chany_top_out[17] ,
    \sb_1__1__31_chany_top_out[18] ,
    \sb_1__1__31_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__36_chany_bottom_out[0] ,
    \cby_1__1__36_chany_bottom_out[1] ,
    \cby_1__1__36_chany_bottom_out[2] ,
    \cby_1__1__36_chany_bottom_out[3] ,
    \cby_1__1__36_chany_bottom_out[4] ,
    \cby_1__1__36_chany_bottom_out[5] ,
    \cby_1__1__36_chany_bottom_out[6] ,
    \cby_1__1__36_chany_bottom_out[7] ,
    \cby_1__1__36_chany_bottom_out[8] ,
    \cby_1__1__36_chany_bottom_out[9] ,
    \cby_1__1__36_chany_bottom_out[10] ,
    \cby_1__1__36_chany_bottom_out[11] ,
    \cby_1__1__36_chany_bottom_out[12] ,
    \cby_1__1__36_chany_bottom_out[13] ,
    \cby_1__1__36_chany_bottom_out[14] ,
    \cby_1__1__36_chany_bottom_out[15] ,
    \cby_1__1__36_chany_bottom_out[16] ,
    \cby_1__1__36_chany_bottom_out[17] ,
    \cby_1__1__36_chany_bottom_out[18] ,
    \cby_1__1__36_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__32_chany_bottom_out[0] ,
    \sb_1__1__32_chany_bottom_out[1] ,
    \sb_1__1__32_chany_bottom_out[2] ,
    \sb_1__1__32_chany_bottom_out[3] ,
    \sb_1__1__32_chany_bottom_out[4] ,
    \sb_1__1__32_chany_bottom_out[5] ,
    \sb_1__1__32_chany_bottom_out[6] ,
    \sb_1__1__32_chany_bottom_out[7] ,
    \sb_1__1__32_chany_bottom_out[8] ,
    \sb_1__1__32_chany_bottom_out[9] ,
    \sb_1__1__32_chany_bottom_out[10] ,
    \sb_1__1__32_chany_bottom_out[11] ,
    \sb_1__1__32_chany_bottom_out[12] ,
    \sb_1__1__32_chany_bottom_out[13] ,
    \sb_1__1__32_chany_bottom_out[14] ,
    \sb_1__1__32_chany_bottom_out[15] ,
    \sb_1__1__32_chany_bottom_out[16] ,
    \sb_1__1__32_chany_bottom_out[17] ,
    \sb_1__1__32_chany_bottom_out[18] ,
    \sb_1__1__32_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__36_chany_top_out[0] ,
    \cby_1__1__36_chany_top_out[1] ,
    \cby_1__1__36_chany_top_out[2] ,
    \cby_1__1__36_chany_top_out[3] ,
    \cby_1__1__36_chany_top_out[4] ,
    \cby_1__1__36_chany_top_out[5] ,
    \cby_1__1__36_chany_top_out[6] ,
    \cby_1__1__36_chany_top_out[7] ,
    \cby_1__1__36_chany_top_out[8] ,
    \cby_1__1__36_chany_top_out[9] ,
    \cby_1__1__36_chany_top_out[10] ,
    \cby_1__1__36_chany_top_out[11] ,
    \cby_1__1__36_chany_top_out[12] ,
    \cby_1__1__36_chany_top_out[13] ,
    \cby_1__1__36_chany_top_out[14] ,
    \cby_1__1__36_chany_top_out[15] ,
    \cby_1__1__36_chany_top_out[16] ,
    \cby_1__1__36_chany_top_out[17] ,
    \cby_1__1__36_chany_top_out[18] ,
    \cby_1__1__36_chany_top_out[19] }));
 cby_1__1_ cby_5__6_ (.Test_en_E_in(\Test_enWires[94] ),
    .Test_en_E_out(\Test_enWires[95] ),
    .Test_en_S_in(\Test_enWires[94] ),
    .Test_en_W_in(\Test_enWires[94] ),
    .ccff_head(grid_clb_37_ccff_tail),
    .ccff_tail(cby_1__1__37_ccff_tail),
    .clk_2_S_in(\clk_2_wires[46] ),
    .clk_2_S_out(\clk_2_wires[47] ),
    .left_grid_pin_16_(cby_1__1__37_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__37_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__37_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__37_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__37_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__37_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__37_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__37_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__37_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__37_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__37_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__37_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__37_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__37_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__37_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__37_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[138] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[137] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[46] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[47] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__32_chany_top_out[0] ,
    \sb_1__1__32_chany_top_out[1] ,
    \sb_1__1__32_chany_top_out[2] ,
    \sb_1__1__32_chany_top_out[3] ,
    \sb_1__1__32_chany_top_out[4] ,
    \sb_1__1__32_chany_top_out[5] ,
    \sb_1__1__32_chany_top_out[6] ,
    \sb_1__1__32_chany_top_out[7] ,
    \sb_1__1__32_chany_top_out[8] ,
    \sb_1__1__32_chany_top_out[9] ,
    \sb_1__1__32_chany_top_out[10] ,
    \sb_1__1__32_chany_top_out[11] ,
    \sb_1__1__32_chany_top_out[12] ,
    \sb_1__1__32_chany_top_out[13] ,
    \sb_1__1__32_chany_top_out[14] ,
    \sb_1__1__32_chany_top_out[15] ,
    \sb_1__1__32_chany_top_out[16] ,
    \sb_1__1__32_chany_top_out[17] ,
    \sb_1__1__32_chany_top_out[18] ,
    \sb_1__1__32_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__37_chany_bottom_out[0] ,
    \cby_1__1__37_chany_bottom_out[1] ,
    \cby_1__1__37_chany_bottom_out[2] ,
    \cby_1__1__37_chany_bottom_out[3] ,
    \cby_1__1__37_chany_bottom_out[4] ,
    \cby_1__1__37_chany_bottom_out[5] ,
    \cby_1__1__37_chany_bottom_out[6] ,
    \cby_1__1__37_chany_bottom_out[7] ,
    \cby_1__1__37_chany_bottom_out[8] ,
    \cby_1__1__37_chany_bottom_out[9] ,
    \cby_1__1__37_chany_bottom_out[10] ,
    \cby_1__1__37_chany_bottom_out[11] ,
    \cby_1__1__37_chany_bottom_out[12] ,
    \cby_1__1__37_chany_bottom_out[13] ,
    \cby_1__1__37_chany_bottom_out[14] ,
    \cby_1__1__37_chany_bottom_out[15] ,
    \cby_1__1__37_chany_bottom_out[16] ,
    \cby_1__1__37_chany_bottom_out[17] ,
    \cby_1__1__37_chany_bottom_out[18] ,
    \cby_1__1__37_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__33_chany_bottom_out[0] ,
    \sb_1__1__33_chany_bottom_out[1] ,
    \sb_1__1__33_chany_bottom_out[2] ,
    \sb_1__1__33_chany_bottom_out[3] ,
    \sb_1__1__33_chany_bottom_out[4] ,
    \sb_1__1__33_chany_bottom_out[5] ,
    \sb_1__1__33_chany_bottom_out[6] ,
    \sb_1__1__33_chany_bottom_out[7] ,
    \sb_1__1__33_chany_bottom_out[8] ,
    \sb_1__1__33_chany_bottom_out[9] ,
    \sb_1__1__33_chany_bottom_out[10] ,
    \sb_1__1__33_chany_bottom_out[11] ,
    \sb_1__1__33_chany_bottom_out[12] ,
    \sb_1__1__33_chany_bottom_out[13] ,
    \sb_1__1__33_chany_bottom_out[14] ,
    \sb_1__1__33_chany_bottom_out[15] ,
    \sb_1__1__33_chany_bottom_out[16] ,
    \sb_1__1__33_chany_bottom_out[17] ,
    \sb_1__1__33_chany_bottom_out[18] ,
    \sb_1__1__33_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__37_chany_top_out[0] ,
    \cby_1__1__37_chany_top_out[1] ,
    \cby_1__1__37_chany_top_out[2] ,
    \cby_1__1__37_chany_top_out[3] ,
    \cby_1__1__37_chany_top_out[4] ,
    \cby_1__1__37_chany_top_out[5] ,
    \cby_1__1__37_chany_top_out[6] ,
    \cby_1__1__37_chany_top_out[7] ,
    \cby_1__1__37_chany_top_out[8] ,
    \cby_1__1__37_chany_top_out[9] ,
    \cby_1__1__37_chany_top_out[10] ,
    \cby_1__1__37_chany_top_out[11] ,
    \cby_1__1__37_chany_top_out[12] ,
    \cby_1__1__37_chany_top_out[13] ,
    \cby_1__1__37_chany_top_out[14] ,
    \cby_1__1__37_chany_top_out[15] ,
    \cby_1__1__37_chany_top_out[16] ,
    \cby_1__1__37_chany_top_out[17] ,
    \cby_1__1__37_chany_top_out[18] ,
    \cby_1__1__37_chany_top_out[19] }));
 cby_1__1_ cby_5__7_ (.Test_en_E_in(\Test_enWires[108] ),
    .Test_en_E_out(\Test_enWires[109] ),
    .Test_en_S_in(\Test_enWires[108] ),
    .Test_en_W_in(\Test_enWires[108] ),
    .ccff_head(grid_clb_38_ccff_tail),
    .ccff_tail(cby_1__1__38_ccff_tail),
    .clk_2_N_out(\clk_2_wires[45] ),
    .clk_2_S_in(\clk_2_wires[44] ),
    .left_grid_pin_16_(cby_1__1__38_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__38_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__38_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__38_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__38_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__38_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__38_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__38_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__38_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__38_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__38_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__38_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__38_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__38_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__38_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__38_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[141] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[140] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[45] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[44] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__33_chany_top_out[0] ,
    \sb_1__1__33_chany_top_out[1] ,
    \sb_1__1__33_chany_top_out[2] ,
    \sb_1__1__33_chany_top_out[3] ,
    \sb_1__1__33_chany_top_out[4] ,
    \sb_1__1__33_chany_top_out[5] ,
    \sb_1__1__33_chany_top_out[6] ,
    \sb_1__1__33_chany_top_out[7] ,
    \sb_1__1__33_chany_top_out[8] ,
    \sb_1__1__33_chany_top_out[9] ,
    \sb_1__1__33_chany_top_out[10] ,
    \sb_1__1__33_chany_top_out[11] ,
    \sb_1__1__33_chany_top_out[12] ,
    \sb_1__1__33_chany_top_out[13] ,
    \sb_1__1__33_chany_top_out[14] ,
    \sb_1__1__33_chany_top_out[15] ,
    \sb_1__1__33_chany_top_out[16] ,
    \sb_1__1__33_chany_top_out[17] ,
    \sb_1__1__33_chany_top_out[18] ,
    \sb_1__1__33_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__38_chany_bottom_out[0] ,
    \cby_1__1__38_chany_bottom_out[1] ,
    \cby_1__1__38_chany_bottom_out[2] ,
    \cby_1__1__38_chany_bottom_out[3] ,
    \cby_1__1__38_chany_bottom_out[4] ,
    \cby_1__1__38_chany_bottom_out[5] ,
    \cby_1__1__38_chany_bottom_out[6] ,
    \cby_1__1__38_chany_bottom_out[7] ,
    \cby_1__1__38_chany_bottom_out[8] ,
    \cby_1__1__38_chany_bottom_out[9] ,
    \cby_1__1__38_chany_bottom_out[10] ,
    \cby_1__1__38_chany_bottom_out[11] ,
    \cby_1__1__38_chany_bottom_out[12] ,
    \cby_1__1__38_chany_bottom_out[13] ,
    \cby_1__1__38_chany_bottom_out[14] ,
    \cby_1__1__38_chany_bottom_out[15] ,
    \cby_1__1__38_chany_bottom_out[16] ,
    \cby_1__1__38_chany_bottom_out[17] ,
    \cby_1__1__38_chany_bottom_out[18] ,
    \cby_1__1__38_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__34_chany_bottom_out[0] ,
    \sb_1__1__34_chany_bottom_out[1] ,
    \sb_1__1__34_chany_bottom_out[2] ,
    \sb_1__1__34_chany_bottom_out[3] ,
    \sb_1__1__34_chany_bottom_out[4] ,
    \sb_1__1__34_chany_bottom_out[5] ,
    \sb_1__1__34_chany_bottom_out[6] ,
    \sb_1__1__34_chany_bottom_out[7] ,
    \sb_1__1__34_chany_bottom_out[8] ,
    \sb_1__1__34_chany_bottom_out[9] ,
    \sb_1__1__34_chany_bottom_out[10] ,
    \sb_1__1__34_chany_bottom_out[11] ,
    \sb_1__1__34_chany_bottom_out[12] ,
    \sb_1__1__34_chany_bottom_out[13] ,
    \sb_1__1__34_chany_bottom_out[14] ,
    \sb_1__1__34_chany_bottom_out[15] ,
    \sb_1__1__34_chany_bottom_out[16] ,
    \sb_1__1__34_chany_bottom_out[17] ,
    \sb_1__1__34_chany_bottom_out[18] ,
    \sb_1__1__34_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__38_chany_top_out[0] ,
    \cby_1__1__38_chany_top_out[1] ,
    \cby_1__1__38_chany_top_out[2] ,
    \cby_1__1__38_chany_top_out[3] ,
    \cby_1__1__38_chany_top_out[4] ,
    \cby_1__1__38_chany_top_out[5] ,
    \cby_1__1__38_chany_top_out[6] ,
    \cby_1__1__38_chany_top_out[7] ,
    \cby_1__1__38_chany_top_out[8] ,
    \cby_1__1__38_chany_top_out[9] ,
    \cby_1__1__38_chany_top_out[10] ,
    \cby_1__1__38_chany_top_out[11] ,
    \cby_1__1__38_chany_top_out[12] ,
    \cby_1__1__38_chany_top_out[13] ,
    \cby_1__1__38_chany_top_out[14] ,
    \cby_1__1__38_chany_top_out[15] ,
    \cby_1__1__38_chany_top_out[16] ,
    \cby_1__1__38_chany_top_out[17] ,
    \cby_1__1__38_chany_top_out[18] ,
    \cby_1__1__38_chany_top_out[19] }));
 cby_1__1_ cby_5__8_ (.Test_en_E_in(\Test_enWires[122] ),
    .Test_en_E_out(\Test_enWires[123] ),
    .Test_en_S_in(\Test_enWires[122] ),
    .Test_en_W_in(\Test_enWires[122] ),
    .ccff_head(grid_clb_39_ccff_tail),
    .ccff_tail(cby_1__1__39_ccff_tail),
    .left_grid_pin_16_(cby_1__1__39_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__39_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__39_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__39_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__39_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__39_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__39_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__39_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__39_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__39_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__39_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__39_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__39_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__39_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__39_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__39_left_grid_pin_31_),
    .prog_clk_0_N_out(\prog_clk_0_wires[146] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[144] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[143] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__34_chany_top_out[0] ,
    \sb_1__1__34_chany_top_out[1] ,
    \sb_1__1__34_chany_top_out[2] ,
    \sb_1__1__34_chany_top_out[3] ,
    \sb_1__1__34_chany_top_out[4] ,
    \sb_1__1__34_chany_top_out[5] ,
    \sb_1__1__34_chany_top_out[6] ,
    \sb_1__1__34_chany_top_out[7] ,
    \sb_1__1__34_chany_top_out[8] ,
    \sb_1__1__34_chany_top_out[9] ,
    \sb_1__1__34_chany_top_out[10] ,
    \sb_1__1__34_chany_top_out[11] ,
    \sb_1__1__34_chany_top_out[12] ,
    \sb_1__1__34_chany_top_out[13] ,
    \sb_1__1__34_chany_top_out[14] ,
    \sb_1__1__34_chany_top_out[15] ,
    \sb_1__1__34_chany_top_out[16] ,
    \sb_1__1__34_chany_top_out[17] ,
    \sb_1__1__34_chany_top_out[18] ,
    \sb_1__1__34_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__39_chany_bottom_out[0] ,
    \cby_1__1__39_chany_bottom_out[1] ,
    \cby_1__1__39_chany_bottom_out[2] ,
    \cby_1__1__39_chany_bottom_out[3] ,
    \cby_1__1__39_chany_bottom_out[4] ,
    \cby_1__1__39_chany_bottom_out[5] ,
    \cby_1__1__39_chany_bottom_out[6] ,
    \cby_1__1__39_chany_bottom_out[7] ,
    \cby_1__1__39_chany_bottom_out[8] ,
    \cby_1__1__39_chany_bottom_out[9] ,
    \cby_1__1__39_chany_bottom_out[10] ,
    \cby_1__1__39_chany_bottom_out[11] ,
    \cby_1__1__39_chany_bottom_out[12] ,
    \cby_1__1__39_chany_bottom_out[13] ,
    \cby_1__1__39_chany_bottom_out[14] ,
    \cby_1__1__39_chany_bottom_out[15] ,
    \cby_1__1__39_chany_bottom_out[16] ,
    \cby_1__1__39_chany_bottom_out[17] ,
    \cby_1__1__39_chany_bottom_out[18] ,
    \cby_1__1__39_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__8__4_chany_bottom_out[0] ,
    \sb_1__8__4_chany_bottom_out[1] ,
    \sb_1__8__4_chany_bottom_out[2] ,
    \sb_1__8__4_chany_bottom_out[3] ,
    \sb_1__8__4_chany_bottom_out[4] ,
    \sb_1__8__4_chany_bottom_out[5] ,
    \sb_1__8__4_chany_bottom_out[6] ,
    \sb_1__8__4_chany_bottom_out[7] ,
    \sb_1__8__4_chany_bottom_out[8] ,
    \sb_1__8__4_chany_bottom_out[9] ,
    \sb_1__8__4_chany_bottom_out[10] ,
    \sb_1__8__4_chany_bottom_out[11] ,
    \sb_1__8__4_chany_bottom_out[12] ,
    \sb_1__8__4_chany_bottom_out[13] ,
    \sb_1__8__4_chany_bottom_out[14] ,
    \sb_1__8__4_chany_bottom_out[15] ,
    \sb_1__8__4_chany_bottom_out[16] ,
    \sb_1__8__4_chany_bottom_out[17] ,
    \sb_1__8__4_chany_bottom_out[18] ,
    \sb_1__8__4_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__39_chany_top_out[0] ,
    \cby_1__1__39_chany_top_out[1] ,
    \cby_1__1__39_chany_top_out[2] ,
    \cby_1__1__39_chany_top_out[3] ,
    \cby_1__1__39_chany_top_out[4] ,
    \cby_1__1__39_chany_top_out[5] ,
    \cby_1__1__39_chany_top_out[6] ,
    \cby_1__1__39_chany_top_out[7] ,
    \cby_1__1__39_chany_top_out[8] ,
    \cby_1__1__39_chany_top_out[9] ,
    \cby_1__1__39_chany_top_out[10] ,
    \cby_1__1__39_chany_top_out[11] ,
    \cby_1__1__39_chany_top_out[12] ,
    \cby_1__1__39_chany_top_out[13] ,
    \cby_1__1__39_chany_top_out[14] ,
    \cby_1__1__39_chany_top_out[15] ,
    \cby_1__1__39_chany_top_out[16] ,
    \cby_1__1__39_chany_top_out[17] ,
    \cby_1__1__39_chany_top_out[18] ,
    \cby_1__1__39_chany_top_out[19] }));
 cby_1__1_ cby_6__1_ (.Test_en_E_in(\Test_enWires[26] ),
    .Test_en_E_out(\Test_enWires[27] ),
    .Test_en_S_in(\Test_enWires[26] ),
    .Test_en_W_in(\Test_enWires[26] ),
    .ccff_head(grid_clb_40_ccff_tail),
    .ccff_tail(cby_1__1__40_ccff_tail),
    .left_grid_pin_16_(cby_1__1__40_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__40_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__40_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__40_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__40_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__40_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__40_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__40_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__40_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__40_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__40_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__40_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__40_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__40_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__40_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__40_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[149] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[148] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__0__5_chany_top_out[0] ,
    \sb_1__0__5_chany_top_out[1] ,
    \sb_1__0__5_chany_top_out[2] ,
    \sb_1__0__5_chany_top_out[3] ,
    \sb_1__0__5_chany_top_out[4] ,
    \sb_1__0__5_chany_top_out[5] ,
    \sb_1__0__5_chany_top_out[6] ,
    \sb_1__0__5_chany_top_out[7] ,
    \sb_1__0__5_chany_top_out[8] ,
    \sb_1__0__5_chany_top_out[9] ,
    \sb_1__0__5_chany_top_out[10] ,
    \sb_1__0__5_chany_top_out[11] ,
    \sb_1__0__5_chany_top_out[12] ,
    \sb_1__0__5_chany_top_out[13] ,
    \sb_1__0__5_chany_top_out[14] ,
    \sb_1__0__5_chany_top_out[15] ,
    \sb_1__0__5_chany_top_out[16] ,
    \sb_1__0__5_chany_top_out[17] ,
    \sb_1__0__5_chany_top_out[18] ,
    \sb_1__0__5_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__40_chany_bottom_out[0] ,
    \cby_1__1__40_chany_bottom_out[1] ,
    \cby_1__1__40_chany_bottom_out[2] ,
    \cby_1__1__40_chany_bottom_out[3] ,
    \cby_1__1__40_chany_bottom_out[4] ,
    \cby_1__1__40_chany_bottom_out[5] ,
    \cby_1__1__40_chany_bottom_out[6] ,
    \cby_1__1__40_chany_bottom_out[7] ,
    \cby_1__1__40_chany_bottom_out[8] ,
    \cby_1__1__40_chany_bottom_out[9] ,
    \cby_1__1__40_chany_bottom_out[10] ,
    \cby_1__1__40_chany_bottom_out[11] ,
    \cby_1__1__40_chany_bottom_out[12] ,
    \cby_1__1__40_chany_bottom_out[13] ,
    \cby_1__1__40_chany_bottom_out[14] ,
    \cby_1__1__40_chany_bottom_out[15] ,
    \cby_1__1__40_chany_bottom_out[16] ,
    \cby_1__1__40_chany_bottom_out[17] ,
    \cby_1__1__40_chany_bottom_out[18] ,
    \cby_1__1__40_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__35_chany_bottom_out[0] ,
    \sb_1__1__35_chany_bottom_out[1] ,
    \sb_1__1__35_chany_bottom_out[2] ,
    \sb_1__1__35_chany_bottom_out[3] ,
    \sb_1__1__35_chany_bottom_out[4] ,
    \sb_1__1__35_chany_bottom_out[5] ,
    \sb_1__1__35_chany_bottom_out[6] ,
    \sb_1__1__35_chany_bottom_out[7] ,
    \sb_1__1__35_chany_bottom_out[8] ,
    \sb_1__1__35_chany_bottom_out[9] ,
    \sb_1__1__35_chany_bottom_out[10] ,
    \sb_1__1__35_chany_bottom_out[11] ,
    \sb_1__1__35_chany_bottom_out[12] ,
    \sb_1__1__35_chany_bottom_out[13] ,
    \sb_1__1__35_chany_bottom_out[14] ,
    \sb_1__1__35_chany_bottom_out[15] ,
    \sb_1__1__35_chany_bottom_out[16] ,
    \sb_1__1__35_chany_bottom_out[17] ,
    \sb_1__1__35_chany_bottom_out[18] ,
    \sb_1__1__35_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__40_chany_top_out[0] ,
    \cby_1__1__40_chany_top_out[1] ,
    \cby_1__1__40_chany_top_out[2] ,
    \cby_1__1__40_chany_top_out[3] ,
    \cby_1__1__40_chany_top_out[4] ,
    \cby_1__1__40_chany_top_out[5] ,
    \cby_1__1__40_chany_top_out[6] ,
    \cby_1__1__40_chany_top_out[7] ,
    \cby_1__1__40_chany_top_out[8] ,
    \cby_1__1__40_chany_top_out[9] ,
    \cby_1__1__40_chany_top_out[10] ,
    \cby_1__1__40_chany_top_out[11] ,
    \cby_1__1__40_chany_top_out[12] ,
    \cby_1__1__40_chany_top_out[13] ,
    \cby_1__1__40_chany_top_out[14] ,
    \cby_1__1__40_chany_top_out[15] ,
    \cby_1__1__40_chany_top_out[16] ,
    \cby_1__1__40_chany_top_out[17] ,
    \cby_1__1__40_chany_top_out[18] ,
    \cby_1__1__40_chany_top_out[19] }));
 cby_1__1_ cby_6__2_ (.Test_en_E_in(\Test_enWires[40] ),
    .Test_en_E_out(\Test_enWires[41] ),
    .Test_en_S_in(\Test_enWires[40] ),
    .Test_en_W_in(\Test_enWires[40] ),
    .ccff_head(grid_clb_41_ccff_tail),
    .ccff_tail(cby_1__1__41_ccff_tail),
    .left_grid_pin_16_(cby_1__1__41_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__41_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__41_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__41_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__41_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__41_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__41_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__41_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__41_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__41_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__41_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__41_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__41_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__41_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__41_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__41_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[152] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[151] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__35_chany_top_out[0] ,
    \sb_1__1__35_chany_top_out[1] ,
    \sb_1__1__35_chany_top_out[2] ,
    \sb_1__1__35_chany_top_out[3] ,
    \sb_1__1__35_chany_top_out[4] ,
    \sb_1__1__35_chany_top_out[5] ,
    \sb_1__1__35_chany_top_out[6] ,
    \sb_1__1__35_chany_top_out[7] ,
    \sb_1__1__35_chany_top_out[8] ,
    \sb_1__1__35_chany_top_out[9] ,
    \sb_1__1__35_chany_top_out[10] ,
    \sb_1__1__35_chany_top_out[11] ,
    \sb_1__1__35_chany_top_out[12] ,
    \sb_1__1__35_chany_top_out[13] ,
    \sb_1__1__35_chany_top_out[14] ,
    \sb_1__1__35_chany_top_out[15] ,
    \sb_1__1__35_chany_top_out[16] ,
    \sb_1__1__35_chany_top_out[17] ,
    \sb_1__1__35_chany_top_out[18] ,
    \sb_1__1__35_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__41_chany_bottom_out[0] ,
    \cby_1__1__41_chany_bottom_out[1] ,
    \cby_1__1__41_chany_bottom_out[2] ,
    \cby_1__1__41_chany_bottom_out[3] ,
    \cby_1__1__41_chany_bottom_out[4] ,
    \cby_1__1__41_chany_bottom_out[5] ,
    \cby_1__1__41_chany_bottom_out[6] ,
    \cby_1__1__41_chany_bottom_out[7] ,
    \cby_1__1__41_chany_bottom_out[8] ,
    \cby_1__1__41_chany_bottom_out[9] ,
    \cby_1__1__41_chany_bottom_out[10] ,
    \cby_1__1__41_chany_bottom_out[11] ,
    \cby_1__1__41_chany_bottom_out[12] ,
    \cby_1__1__41_chany_bottom_out[13] ,
    \cby_1__1__41_chany_bottom_out[14] ,
    \cby_1__1__41_chany_bottom_out[15] ,
    \cby_1__1__41_chany_bottom_out[16] ,
    \cby_1__1__41_chany_bottom_out[17] ,
    \cby_1__1__41_chany_bottom_out[18] ,
    \cby_1__1__41_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__36_chany_bottom_out[0] ,
    \sb_1__1__36_chany_bottom_out[1] ,
    \sb_1__1__36_chany_bottom_out[2] ,
    \sb_1__1__36_chany_bottom_out[3] ,
    \sb_1__1__36_chany_bottom_out[4] ,
    \sb_1__1__36_chany_bottom_out[5] ,
    \sb_1__1__36_chany_bottom_out[6] ,
    \sb_1__1__36_chany_bottom_out[7] ,
    \sb_1__1__36_chany_bottom_out[8] ,
    \sb_1__1__36_chany_bottom_out[9] ,
    \sb_1__1__36_chany_bottom_out[10] ,
    \sb_1__1__36_chany_bottom_out[11] ,
    \sb_1__1__36_chany_bottom_out[12] ,
    \sb_1__1__36_chany_bottom_out[13] ,
    \sb_1__1__36_chany_bottom_out[14] ,
    \sb_1__1__36_chany_bottom_out[15] ,
    \sb_1__1__36_chany_bottom_out[16] ,
    \sb_1__1__36_chany_bottom_out[17] ,
    \sb_1__1__36_chany_bottom_out[18] ,
    \sb_1__1__36_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__41_chany_top_out[0] ,
    \cby_1__1__41_chany_top_out[1] ,
    \cby_1__1__41_chany_top_out[2] ,
    \cby_1__1__41_chany_top_out[3] ,
    \cby_1__1__41_chany_top_out[4] ,
    \cby_1__1__41_chany_top_out[5] ,
    \cby_1__1__41_chany_top_out[6] ,
    \cby_1__1__41_chany_top_out[7] ,
    \cby_1__1__41_chany_top_out[8] ,
    \cby_1__1__41_chany_top_out[9] ,
    \cby_1__1__41_chany_top_out[10] ,
    \cby_1__1__41_chany_top_out[11] ,
    \cby_1__1__41_chany_top_out[12] ,
    \cby_1__1__41_chany_top_out[13] ,
    \cby_1__1__41_chany_top_out[14] ,
    \cby_1__1__41_chany_top_out[15] ,
    \cby_1__1__41_chany_top_out[16] ,
    \cby_1__1__41_chany_top_out[17] ,
    \cby_1__1__41_chany_top_out[18] ,
    \cby_1__1__41_chany_top_out[19] }));
 cby_1__1_ cby_6__3_ (.Test_en_E_in(\Test_enWires[54] ),
    .Test_en_E_out(\Test_enWires[55] ),
    .Test_en_S_in(\Test_enWires[54] ),
    .Test_en_W_in(\Test_enWires[54] ),
    .ccff_head(grid_clb_42_ccff_tail),
    .ccff_tail(cby_1__1__42_ccff_tail),
    .clk_3_S_in(\clk_3_wires[24] ),
    .clk_3_S_out(\clk_3_wires[25] ),
    .left_grid_pin_16_(cby_1__1__42_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__42_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__42_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__42_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__42_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__42_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__42_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__42_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__42_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__42_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__42_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__42_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__42_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__42_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__42_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__42_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[155] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[154] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[24] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[25] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__36_chany_top_out[0] ,
    \sb_1__1__36_chany_top_out[1] ,
    \sb_1__1__36_chany_top_out[2] ,
    \sb_1__1__36_chany_top_out[3] ,
    \sb_1__1__36_chany_top_out[4] ,
    \sb_1__1__36_chany_top_out[5] ,
    \sb_1__1__36_chany_top_out[6] ,
    \sb_1__1__36_chany_top_out[7] ,
    \sb_1__1__36_chany_top_out[8] ,
    \sb_1__1__36_chany_top_out[9] ,
    \sb_1__1__36_chany_top_out[10] ,
    \sb_1__1__36_chany_top_out[11] ,
    \sb_1__1__36_chany_top_out[12] ,
    \sb_1__1__36_chany_top_out[13] ,
    \sb_1__1__36_chany_top_out[14] ,
    \sb_1__1__36_chany_top_out[15] ,
    \sb_1__1__36_chany_top_out[16] ,
    \sb_1__1__36_chany_top_out[17] ,
    \sb_1__1__36_chany_top_out[18] ,
    \sb_1__1__36_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__42_chany_bottom_out[0] ,
    \cby_1__1__42_chany_bottom_out[1] ,
    \cby_1__1__42_chany_bottom_out[2] ,
    \cby_1__1__42_chany_bottom_out[3] ,
    \cby_1__1__42_chany_bottom_out[4] ,
    \cby_1__1__42_chany_bottom_out[5] ,
    \cby_1__1__42_chany_bottom_out[6] ,
    \cby_1__1__42_chany_bottom_out[7] ,
    \cby_1__1__42_chany_bottom_out[8] ,
    \cby_1__1__42_chany_bottom_out[9] ,
    \cby_1__1__42_chany_bottom_out[10] ,
    \cby_1__1__42_chany_bottom_out[11] ,
    \cby_1__1__42_chany_bottom_out[12] ,
    \cby_1__1__42_chany_bottom_out[13] ,
    \cby_1__1__42_chany_bottom_out[14] ,
    \cby_1__1__42_chany_bottom_out[15] ,
    \cby_1__1__42_chany_bottom_out[16] ,
    \cby_1__1__42_chany_bottom_out[17] ,
    \cby_1__1__42_chany_bottom_out[18] ,
    \cby_1__1__42_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__37_chany_bottom_out[0] ,
    \sb_1__1__37_chany_bottom_out[1] ,
    \sb_1__1__37_chany_bottom_out[2] ,
    \sb_1__1__37_chany_bottom_out[3] ,
    \sb_1__1__37_chany_bottom_out[4] ,
    \sb_1__1__37_chany_bottom_out[5] ,
    \sb_1__1__37_chany_bottom_out[6] ,
    \sb_1__1__37_chany_bottom_out[7] ,
    \sb_1__1__37_chany_bottom_out[8] ,
    \sb_1__1__37_chany_bottom_out[9] ,
    \sb_1__1__37_chany_bottom_out[10] ,
    \sb_1__1__37_chany_bottom_out[11] ,
    \sb_1__1__37_chany_bottom_out[12] ,
    \sb_1__1__37_chany_bottom_out[13] ,
    \sb_1__1__37_chany_bottom_out[14] ,
    \sb_1__1__37_chany_bottom_out[15] ,
    \sb_1__1__37_chany_bottom_out[16] ,
    \sb_1__1__37_chany_bottom_out[17] ,
    \sb_1__1__37_chany_bottom_out[18] ,
    \sb_1__1__37_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__42_chany_top_out[0] ,
    \cby_1__1__42_chany_top_out[1] ,
    \cby_1__1__42_chany_top_out[2] ,
    \cby_1__1__42_chany_top_out[3] ,
    \cby_1__1__42_chany_top_out[4] ,
    \cby_1__1__42_chany_top_out[5] ,
    \cby_1__1__42_chany_top_out[6] ,
    \cby_1__1__42_chany_top_out[7] ,
    \cby_1__1__42_chany_top_out[8] ,
    \cby_1__1__42_chany_top_out[9] ,
    \cby_1__1__42_chany_top_out[10] ,
    \cby_1__1__42_chany_top_out[11] ,
    \cby_1__1__42_chany_top_out[12] ,
    \cby_1__1__42_chany_top_out[13] ,
    \cby_1__1__42_chany_top_out[14] ,
    \cby_1__1__42_chany_top_out[15] ,
    \cby_1__1__42_chany_top_out[16] ,
    \cby_1__1__42_chany_top_out[17] ,
    \cby_1__1__42_chany_top_out[18] ,
    \cby_1__1__42_chany_top_out[19] }));
 cby_1__1_ cby_6__4_ (.Test_en_E_in(\Test_enWires[68] ),
    .Test_en_E_out(\Test_enWires[69] ),
    .Test_en_S_in(\Test_enWires[68] ),
    .Test_en_W_in(\Test_enWires[68] ),
    .ccff_head(grid_clb_43_ccff_tail),
    .ccff_tail(cby_1__1__43_ccff_tail),
    .clk_3_S_in(\clk_3_wires[20] ),
    .clk_3_S_out(\clk_3_wires[21] ),
    .left_grid_pin_16_(cby_1__1__43_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__43_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__43_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__43_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__43_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__43_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__43_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__43_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__43_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__43_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__43_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__43_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__43_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__43_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__43_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__43_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[158] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[157] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[20] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[21] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__37_chany_top_out[0] ,
    \sb_1__1__37_chany_top_out[1] ,
    \sb_1__1__37_chany_top_out[2] ,
    \sb_1__1__37_chany_top_out[3] ,
    \sb_1__1__37_chany_top_out[4] ,
    \sb_1__1__37_chany_top_out[5] ,
    \sb_1__1__37_chany_top_out[6] ,
    \sb_1__1__37_chany_top_out[7] ,
    \sb_1__1__37_chany_top_out[8] ,
    \sb_1__1__37_chany_top_out[9] ,
    \sb_1__1__37_chany_top_out[10] ,
    \sb_1__1__37_chany_top_out[11] ,
    \sb_1__1__37_chany_top_out[12] ,
    \sb_1__1__37_chany_top_out[13] ,
    \sb_1__1__37_chany_top_out[14] ,
    \sb_1__1__37_chany_top_out[15] ,
    \sb_1__1__37_chany_top_out[16] ,
    \sb_1__1__37_chany_top_out[17] ,
    \sb_1__1__37_chany_top_out[18] ,
    \sb_1__1__37_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__43_chany_bottom_out[0] ,
    \cby_1__1__43_chany_bottom_out[1] ,
    \cby_1__1__43_chany_bottom_out[2] ,
    \cby_1__1__43_chany_bottom_out[3] ,
    \cby_1__1__43_chany_bottom_out[4] ,
    \cby_1__1__43_chany_bottom_out[5] ,
    \cby_1__1__43_chany_bottom_out[6] ,
    \cby_1__1__43_chany_bottom_out[7] ,
    \cby_1__1__43_chany_bottom_out[8] ,
    \cby_1__1__43_chany_bottom_out[9] ,
    \cby_1__1__43_chany_bottom_out[10] ,
    \cby_1__1__43_chany_bottom_out[11] ,
    \cby_1__1__43_chany_bottom_out[12] ,
    \cby_1__1__43_chany_bottom_out[13] ,
    \cby_1__1__43_chany_bottom_out[14] ,
    \cby_1__1__43_chany_bottom_out[15] ,
    \cby_1__1__43_chany_bottom_out[16] ,
    \cby_1__1__43_chany_bottom_out[17] ,
    \cby_1__1__43_chany_bottom_out[18] ,
    \cby_1__1__43_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__38_chany_bottom_out[0] ,
    \sb_1__1__38_chany_bottom_out[1] ,
    \sb_1__1__38_chany_bottom_out[2] ,
    \sb_1__1__38_chany_bottom_out[3] ,
    \sb_1__1__38_chany_bottom_out[4] ,
    \sb_1__1__38_chany_bottom_out[5] ,
    \sb_1__1__38_chany_bottom_out[6] ,
    \sb_1__1__38_chany_bottom_out[7] ,
    \sb_1__1__38_chany_bottom_out[8] ,
    \sb_1__1__38_chany_bottom_out[9] ,
    \sb_1__1__38_chany_bottom_out[10] ,
    \sb_1__1__38_chany_bottom_out[11] ,
    \sb_1__1__38_chany_bottom_out[12] ,
    \sb_1__1__38_chany_bottom_out[13] ,
    \sb_1__1__38_chany_bottom_out[14] ,
    \sb_1__1__38_chany_bottom_out[15] ,
    \sb_1__1__38_chany_bottom_out[16] ,
    \sb_1__1__38_chany_bottom_out[17] ,
    \sb_1__1__38_chany_bottom_out[18] ,
    \sb_1__1__38_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__43_chany_top_out[0] ,
    \cby_1__1__43_chany_top_out[1] ,
    \cby_1__1__43_chany_top_out[2] ,
    \cby_1__1__43_chany_top_out[3] ,
    \cby_1__1__43_chany_top_out[4] ,
    \cby_1__1__43_chany_top_out[5] ,
    \cby_1__1__43_chany_top_out[6] ,
    \cby_1__1__43_chany_top_out[7] ,
    \cby_1__1__43_chany_top_out[8] ,
    \cby_1__1__43_chany_top_out[9] ,
    \cby_1__1__43_chany_top_out[10] ,
    \cby_1__1__43_chany_top_out[11] ,
    \cby_1__1__43_chany_top_out[12] ,
    \cby_1__1__43_chany_top_out[13] ,
    \cby_1__1__43_chany_top_out[14] ,
    \cby_1__1__43_chany_top_out[15] ,
    \cby_1__1__43_chany_top_out[16] ,
    \cby_1__1__43_chany_top_out[17] ,
    \cby_1__1__43_chany_top_out[18] ,
    \cby_1__1__43_chany_top_out[19] }));
 cby_1__1_ cby_6__5_ (.Test_en_E_in(\Test_enWires[82] ),
    .Test_en_E_out(\Test_enWires[83] ),
    .Test_en_S_in(\Test_enWires[82] ),
    .Test_en_W_in(\Test_enWires[82] ),
    .ccff_head(grid_clb_44_ccff_tail),
    .ccff_tail(cby_1__1__44_ccff_tail),
    .clk_3_N_out(\clk_3_wires[19] ),
    .clk_3_S_in(\clk_3_wires[18] ),
    .left_grid_pin_16_(cby_1__1__44_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__44_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__44_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__44_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__44_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__44_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__44_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__44_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__44_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__44_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__44_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__44_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__44_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__44_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__44_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__44_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[161] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[160] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[19] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[18] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__38_chany_top_out[0] ,
    \sb_1__1__38_chany_top_out[1] ,
    \sb_1__1__38_chany_top_out[2] ,
    \sb_1__1__38_chany_top_out[3] ,
    \sb_1__1__38_chany_top_out[4] ,
    \sb_1__1__38_chany_top_out[5] ,
    \sb_1__1__38_chany_top_out[6] ,
    \sb_1__1__38_chany_top_out[7] ,
    \sb_1__1__38_chany_top_out[8] ,
    \sb_1__1__38_chany_top_out[9] ,
    \sb_1__1__38_chany_top_out[10] ,
    \sb_1__1__38_chany_top_out[11] ,
    \sb_1__1__38_chany_top_out[12] ,
    \sb_1__1__38_chany_top_out[13] ,
    \sb_1__1__38_chany_top_out[14] ,
    \sb_1__1__38_chany_top_out[15] ,
    \sb_1__1__38_chany_top_out[16] ,
    \sb_1__1__38_chany_top_out[17] ,
    \sb_1__1__38_chany_top_out[18] ,
    \sb_1__1__38_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__44_chany_bottom_out[0] ,
    \cby_1__1__44_chany_bottom_out[1] ,
    \cby_1__1__44_chany_bottom_out[2] ,
    \cby_1__1__44_chany_bottom_out[3] ,
    \cby_1__1__44_chany_bottom_out[4] ,
    \cby_1__1__44_chany_bottom_out[5] ,
    \cby_1__1__44_chany_bottom_out[6] ,
    \cby_1__1__44_chany_bottom_out[7] ,
    \cby_1__1__44_chany_bottom_out[8] ,
    \cby_1__1__44_chany_bottom_out[9] ,
    \cby_1__1__44_chany_bottom_out[10] ,
    \cby_1__1__44_chany_bottom_out[11] ,
    \cby_1__1__44_chany_bottom_out[12] ,
    \cby_1__1__44_chany_bottom_out[13] ,
    \cby_1__1__44_chany_bottom_out[14] ,
    \cby_1__1__44_chany_bottom_out[15] ,
    \cby_1__1__44_chany_bottom_out[16] ,
    \cby_1__1__44_chany_bottom_out[17] ,
    \cby_1__1__44_chany_bottom_out[18] ,
    \cby_1__1__44_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__39_chany_bottom_out[0] ,
    \sb_1__1__39_chany_bottom_out[1] ,
    \sb_1__1__39_chany_bottom_out[2] ,
    \sb_1__1__39_chany_bottom_out[3] ,
    \sb_1__1__39_chany_bottom_out[4] ,
    \sb_1__1__39_chany_bottom_out[5] ,
    \sb_1__1__39_chany_bottom_out[6] ,
    \sb_1__1__39_chany_bottom_out[7] ,
    \sb_1__1__39_chany_bottom_out[8] ,
    \sb_1__1__39_chany_bottom_out[9] ,
    \sb_1__1__39_chany_bottom_out[10] ,
    \sb_1__1__39_chany_bottom_out[11] ,
    \sb_1__1__39_chany_bottom_out[12] ,
    \sb_1__1__39_chany_bottom_out[13] ,
    \sb_1__1__39_chany_bottom_out[14] ,
    \sb_1__1__39_chany_bottom_out[15] ,
    \sb_1__1__39_chany_bottom_out[16] ,
    \sb_1__1__39_chany_bottom_out[17] ,
    \sb_1__1__39_chany_bottom_out[18] ,
    \sb_1__1__39_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__44_chany_top_out[0] ,
    \cby_1__1__44_chany_top_out[1] ,
    \cby_1__1__44_chany_top_out[2] ,
    \cby_1__1__44_chany_top_out[3] ,
    \cby_1__1__44_chany_top_out[4] ,
    \cby_1__1__44_chany_top_out[5] ,
    \cby_1__1__44_chany_top_out[6] ,
    \cby_1__1__44_chany_top_out[7] ,
    \cby_1__1__44_chany_top_out[8] ,
    \cby_1__1__44_chany_top_out[9] ,
    \cby_1__1__44_chany_top_out[10] ,
    \cby_1__1__44_chany_top_out[11] ,
    \cby_1__1__44_chany_top_out[12] ,
    \cby_1__1__44_chany_top_out[13] ,
    \cby_1__1__44_chany_top_out[14] ,
    \cby_1__1__44_chany_top_out[15] ,
    \cby_1__1__44_chany_top_out[16] ,
    \cby_1__1__44_chany_top_out[17] ,
    \cby_1__1__44_chany_top_out[18] ,
    \cby_1__1__44_chany_top_out[19] }));
 cby_1__1_ cby_6__6_ (.Test_en_E_in(\Test_enWires[96] ),
    .Test_en_E_out(\Test_enWires[97] ),
    .Test_en_S_in(\Test_enWires[96] ),
    .Test_en_W_in(\Test_enWires[96] ),
    .ccff_head(grid_clb_45_ccff_tail),
    .ccff_tail(cby_1__1__45_ccff_tail),
    .clk_3_N_out(\clk_3_wires[23] ),
    .clk_3_S_in(\clk_3_wires[22] ),
    .left_grid_pin_16_(cby_1__1__45_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__45_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__45_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__45_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__45_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__45_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__45_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__45_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__45_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__45_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__45_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__45_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__45_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__45_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__45_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__45_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[164] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[163] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[23] ),
    .prog_clk_3_S_in(\prog_clk_3_wires[22] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__39_chany_top_out[0] ,
    \sb_1__1__39_chany_top_out[1] ,
    \sb_1__1__39_chany_top_out[2] ,
    \sb_1__1__39_chany_top_out[3] ,
    \sb_1__1__39_chany_top_out[4] ,
    \sb_1__1__39_chany_top_out[5] ,
    \sb_1__1__39_chany_top_out[6] ,
    \sb_1__1__39_chany_top_out[7] ,
    \sb_1__1__39_chany_top_out[8] ,
    \sb_1__1__39_chany_top_out[9] ,
    \sb_1__1__39_chany_top_out[10] ,
    \sb_1__1__39_chany_top_out[11] ,
    \sb_1__1__39_chany_top_out[12] ,
    \sb_1__1__39_chany_top_out[13] ,
    \sb_1__1__39_chany_top_out[14] ,
    \sb_1__1__39_chany_top_out[15] ,
    \sb_1__1__39_chany_top_out[16] ,
    \sb_1__1__39_chany_top_out[17] ,
    \sb_1__1__39_chany_top_out[18] ,
    \sb_1__1__39_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__45_chany_bottom_out[0] ,
    \cby_1__1__45_chany_bottom_out[1] ,
    \cby_1__1__45_chany_bottom_out[2] ,
    \cby_1__1__45_chany_bottom_out[3] ,
    \cby_1__1__45_chany_bottom_out[4] ,
    \cby_1__1__45_chany_bottom_out[5] ,
    \cby_1__1__45_chany_bottom_out[6] ,
    \cby_1__1__45_chany_bottom_out[7] ,
    \cby_1__1__45_chany_bottom_out[8] ,
    \cby_1__1__45_chany_bottom_out[9] ,
    \cby_1__1__45_chany_bottom_out[10] ,
    \cby_1__1__45_chany_bottom_out[11] ,
    \cby_1__1__45_chany_bottom_out[12] ,
    \cby_1__1__45_chany_bottom_out[13] ,
    \cby_1__1__45_chany_bottom_out[14] ,
    \cby_1__1__45_chany_bottom_out[15] ,
    \cby_1__1__45_chany_bottom_out[16] ,
    \cby_1__1__45_chany_bottom_out[17] ,
    \cby_1__1__45_chany_bottom_out[18] ,
    \cby_1__1__45_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__40_chany_bottom_out[0] ,
    \sb_1__1__40_chany_bottom_out[1] ,
    \sb_1__1__40_chany_bottom_out[2] ,
    \sb_1__1__40_chany_bottom_out[3] ,
    \sb_1__1__40_chany_bottom_out[4] ,
    \sb_1__1__40_chany_bottom_out[5] ,
    \sb_1__1__40_chany_bottom_out[6] ,
    \sb_1__1__40_chany_bottom_out[7] ,
    \sb_1__1__40_chany_bottom_out[8] ,
    \sb_1__1__40_chany_bottom_out[9] ,
    \sb_1__1__40_chany_bottom_out[10] ,
    \sb_1__1__40_chany_bottom_out[11] ,
    \sb_1__1__40_chany_bottom_out[12] ,
    \sb_1__1__40_chany_bottom_out[13] ,
    \sb_1__1__40_chany_bottom_out[14] ,
    \sb_1__1__40_chany_bottom_out[15] ,
    \sb_1__1__40_chany_bottom_out[16] ,
    \sb_1__1__40_chany_bottom_out[17] ,
    \sb_1__1__40_chany_bottom_out[18] ,
    \sb_1__1__40_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__45_chany_top_out[0] ,
    \cby_1__1__45_chany_top_out[1] ,
    \cby_1__1__45_chany_top_out[2] ,
    \cby_1__1__45_chany_top_out[3] ,
    \cby_1__1__45_chany_top_out[4] ,
    \cby_1__1__45_chany_top_out[5] ,
    \cby_1__1__45_chany_top_out[6] ,
    \cby_1__1__45_chany_top_out[7] ,
    \cby_1__1__45_chany_top_out[8] ,
    \cby_1__1__45_chany_top_out[9] ,
    \cby_1__1__45_chany_top_out[10] ,
    \cby_1__1__45_chany_top_out[11] ,
    \cby_1__1__45_chany_top_out[12] ,
    \cby_1__1__45_chany_top_out[13] ,
    \cby_1__1__45_chany_top_out[14] ,
    \cby_1__1__45_chany_top_out[15] ,
    \cby_1__1__45_chany_top_out[16] ,
    \cby_1__1__45_chany_top_out[17] ,
    \cby_1__1__45_chany_top_out[18] ,
    \cby_1__1__45_chany_top_out[19] }));
 cby_1__1_ cby_6__7_ (.Test_en_E_in(\Test_enWires[110] ),
    .Test_en_E_out(\Test_enWires[111] ),
    .Test_en_S_in(\Test_enWires[110] ),
    .Test_en_W_in(\Test_enWires[110] ),
    .ccff_head(grid_clb_46_ccff_tail),
    .ccff_tail(cby_1__1__46_ccff_tail),
    .left_grid_pin_16_(cby_1__1__46_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__46_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__46_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__46_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__46_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__46_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__46_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__46_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__46_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__46_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__46_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__46_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__46_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__46_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__46_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__46_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[167] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[166] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__40_chany_top_out[0] ,
    \sb_1__1__40_chany_top_out[1] ,
    \sb_1__1__40_chany_top_out[2] ,
    \sb_1__1__40_chany_top_out[3] ,
    \sb_1__1__40_chany_top_out[4] ,
    \sb_1__1__40_chany_top_out[5] ,
    \sb_1__1__40_chany_top_out[6] ,
    \sb_1__1__40_chany_top_out[7] ,
    \sb_1__1__40_chany_top_out[8] ,
    \sb_1__1__40_chany_top_out[9] ,
    \sb_1__1__40_chany_top_out[10] ,
    \sb_1__1__40_chany_top_out[11] ,
    \sb_1__1__40_chany_top_out[12] ,
    \sb_1__1__40_chany_top_out[13] ,
    \sb_1__1__40_chany_top_out[14] ,
    \sb_1__1__40_chany_top_out[15] ,
    \sb_1__1__40_chany_top_out[16] ,
    \sb_1__1__40_chany_top_out[17] ,
    \sb_1__1__40_chany_top_out[18] ,
    \sb_1__1__40_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__46_chany_bottom_out[0] ,
    \cby_1__1__46_chany_bottom_out[1] ,
    \cby_1__1__46_chany_bottom_out[2] ,
    \cby_1__1__46_chany_bottom_out[3] ,
    \cby_1__1__46_chany_bottom_out[4] ,
    \cby_1__1__46_chany_bottom_out[5] ,
    \cby_1__1__46_chany_bottom_out[6] ,
    \cby_1__1__46_chany_bottom_out[7] ,
    \cby_1__1__46_chany_bottom_out[8] ,
    \cby_1__1__46_chany_bottom_out[9] ,
    \cby_1__1__46_chany_bottom_out[10] ,
    \cby_1__1__46_chany_bottom_out[11] ,
    \cby_1__1__46_chany_bottom_out[12] ,
    \cby_1__1__46_chany_bottom_out[13] ,
    \cby_1__1__46_chany_bottom_out[14] ,
    \cby_1__1__46_chany_bottom_out[15] ,
    \cby_1__1__46_chany_bottom_out[16] ,
    \cby_1__1__46_chany_bottom_out[17] ,
    \cby_1__1__46_chany_bottom_out[18] ,
    \cby_1__1__46_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__41_chany_bottom_out[0] ,
    \sb_1__1__41_chany_bottom_out[1] ,
    \sb_1__1__41_chany_bottom_out[2] ,
    \sb_1__1__41_chany_bottom_out[3] ,
    \sb_1__1__41_chany_bottom_out[4] ,
    \sb_1__1__41_chany_bottom_out[5] ,
    \sb_1__1__41_chany_bottom_out[6] ,
    \sb_1__1__41_chany_bottom_out[7] ,
    \sb_1__1__41_chany_bottom_out[8] ,
    \sb_1__1__41_chany_bottom_out[9] ,
    \sb_1__1__41_chany_bottom_out[10] ,
    \sb_1__1__41_chany_bottom_out[11] ,
    \sb_1__1__41_chany_bottom_out[12] ,
    \sb_1__1__41_chany_bottom_out[13] ,
    \sb_1__1__41_chany_bottom_out[14] ,
    \sb_1__1__41_chany_bottom_out[15] ,
    \sb_1__1__41_chany_bottom_out[16] ,
    \sb_1__1__41_chany_bottom_out[17] ,
    \sb_1__1__41_chany_bottom_out[18] ,
    \sb_1__1__41_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__46_chany_top_out[0] ,
    \cby_1__1__46_chany_top_out[1] ,
    \cby_1__1__46_chany_top_out[2] ,
    \cby_1__1__46_chany_top_out[3] ,
    \cby_1__1__46_chany_top_out[4] ,
    \cby_1__1__46_chany_top_out[5] ,
    \cby_1__1__46_chany_top_out[6] ,
    \cby_1__1__46_chany_top_out[7] ,
    \cby_1__1__46_chany_top_out[8] ,
    \cby_1__1__46_chany_top_out[9] ,
    \cby_1__1__46_chany_top_out[10] ,
    \cby_1__1__46_chany_top_out[11] ,
    \cby_1__1__46_chany_top_out[12] ,
    \cby_1__1__46_chany_top_out[13] ,
    \cby_1__1__46_chany_top_out[14] ,
    \cby_1__1__46_chany_top_out[15] ,
    \cby_1__1__46_chany_top_out[16] ,
    \cby_1__1__46_chany_top_out[17] ,
    \cby_1__1__46_chany_top_out[18] ,
    \cby_1__1__46_chany_top_out[19] }));
 cby_1__1_ cby_6__8_ (.Test_en_E_in(\Test_enWires[124] ),
    .Test_en_E_out(\Test_enWires[125] ),
    .Test_en_S_in(\Test_enWires[124] ),
    .Test_en_W_in(\Test_enWires[124] ),
    .ccff_head(grid_clb_47_ccff_tail),
    .ccff_tail(cby_1__1__47_ccff_tail),
    .left_grid_pin_16_(cby_1__1__47_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__47_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__47_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__47_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__47_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__47_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__47_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__47_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__47_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__47_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__47_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__47_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__47_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__47_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__47_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__47_left_grid_pin_31_),
    .prog_clk_0_N_out(\prog_clk_0_wires[172] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[170] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[169] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__41_chany_top_out[0] ,
    \sb_1__1__41_chany_top_out[1] ,
    \sb_1__1__41_chany_top_out[2] ,
    \sb_1__1__41_chany_top_out[3] ,
    \sb_1__1__41_chany_top_out[4] ,
    \sb_1__1__41_chany_top_out[5] ,
    \sb_1__1__41_chany_top_out[6] ,
    \sb_1__1__41_chany_top_out[7] ,
    \sb_1__1__41_chany_top_out[8] ,
    \sb_1__1__41_chany_top_out[9] ,
    \sb_1__1__41_chany_top_out[10] ,
    \sb_1__1__41_chany_top_out[11] ,
    \sb_1__1__41_chany_top_out[12] ,
    \sb_1__1__41_chany_top_out[13] ,
    \sb_1__1__41_chany_top_out[14] ,
    \sb_1__1__41_chany_top_out[15] ,
    \sb_1__1__41_chany_top_out[16] ,
    \sb_1__1__41_chany_top_out[17] ,
    \sb_1__1__41_chany_top_out[18] ,
    \sb_1__1__41_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__47_chany_bottom_out[0] ,
    \cby_1__1__47_chany_bottom_out[1] ,
    \cby_1__1__47_chany_bottom_out[2] ,
    \cby_1__1__47_chany_bottom_out[3] ,
    \cby_1__1__47_chany_bottom_out[4] ,
    \cby_1__1__47_chany_bottom_out[5] ,
    \cby_1__1__47_chany_bottom_out[6] ,
    \cby_1__1__47_chany_bottom_out[7] ,
    \cby_1__1__47_chany_bottom_out[8] ,
    \cby_1__1__47_chany_bottom_out[9] ,
    \cby_1__1__47_chany_bottom_out[10] ,
    \cby_1__1__47_chany_bottom_out[11] ,
    \cby_1__1__47_chany_bottom_out[12] ,
    \cby_1__1__47_chany_bottom_out[13] ,
    \cby_1__1__47_chany_bottom_out[14] ,
    \cby_1__1__47_chany_bottom_out[15] ,
    \cby_1__1__47_chany_bottom_out[16] ,
    \cby_1__1__47_chany_bottom_out[17] ,
    \cby_1__1__47_chany_bottom_out[18] ,
    \cby_1__1__47_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__8__5_chany_bottom_out[0] ,
    \sb_1__8__5_chany_bottom_out[1] ,
    \sb_1__8__5_chany_bottom_out[2] ,
    \sb_1__8__5_chany_bottom_out[3] ,
    \sb_1__8__5_chany_bottom_out[4] ,
    \sb_1__8__5_chany_bottom_out[5] ,
    \sb_1__8__5_chany_bottom_out[6] ,
    \sb_1__8__5_chany_bottom_out[7] ,
    \sb_1__8__5_chany_bottom_out[8] ,
    \sb_1__8__5_chany_bottom_out[9] ,
    \sb_1__8__5_chany_bottom_out[10] ,
    \sb_1__8__5_chany_bottom_out[11] ,
    \sb_1__8__5_chany_bottom_out[12] ,
    \sb_1__8__5_chany_bottom_out[13] ,
    \sb_1__8__5_chany_bottom_out[14] ,
    \sb_1__8__5_chany_bottom_out[15] ,
    \sb_1__8__5_chany_bottom_out[16] ,
    \sb_1__8__5_chany_bottom_out[17] ,
    \sb_1__8__5_chany_bottom_out[18] ,
    \sb_1__8__5_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__47_chany_top_out[0] ,
    \cby_1__1__47_chany_top_out[1] ,
    \cby_1__1__47_chany_top_out[2] ,
    \cby_1__1__47_chany_top_out[3] ,
    \cby_1__1__47_chany_top_out[4] ,
    \cby_1__1__47_chany_top_out[5] ,
    \cby_1__1__47_chany_top_out[6] ,
    \cby_1__1__47_chany_top_out[7] ,
    \cby_1__1__47_chany_top_out[8] ,
    \cby_1__1__47_chany_top_out[9] ,
    \cby_1__1__47_chany_top_out[10] ,
    \cby_1__1__47_chany_top_out[11] ,
    \cby_1__1__47_chany_top_out[12] ,
    \cby_1__1__47_chany_top_out[13] ,
    \cby_1__1__47_chany_top_out[14] ,
    \cby_1__1__47_chany_top_out[15] ,
    \cby_1__1__47_chany_top_out[16] ,
    \cby_1__1__47_chany_top_out[17] ,
    \cby_1__1__47_chany_top_out[18] ,
    \cby_1__1__47_chany_top_out[19] }));
 cby_1__1_ cby_7__1_ (.Test_en_E_in(\Test_enWires[28] ),
    .Test_en_E_out(\Test_enWires[29] ),
    .Test_en_S_in(\Test_enWires[28] ),
    .Test_en_W_in(\Test_enWires[28] ),
    .ccff_head(grid_clb_48_ccff_tail),
    .ccff_tail(cby_1__1__48_ccff_tail),
    .left_grid_pin_16_(cby_1__1__48_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__48_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__48_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__48_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__48_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__48_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__48_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__48_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__48_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__48_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__48_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__48_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__48_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__48_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__48_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__48_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[175] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[174] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__0__6_chany_top_out[0] ,
    \sb_1__0__6_chany_top_out[1] ,
    \sb_1__0__6_chany_top_out[2] ,
    \sb_1__0__6_chany_top_out[3] ,
    \sb_1__0__6_chany_top_out[4] ,
    \sb_1__0__6_chany_top_out[5] ,
    \sb_1__0__6_chany_top_out[6] ,
    \sb_1__0__6_chany_top_out[7] ,
    \sb_1__0__6_chany_top_out[8] ,
    \sb_1__0__6_chany_top_out[9] ,
    \sb_1__0__6_chany_top_out[10] ,
    \sb_1__0__6_chany_top_out[11] ,
    \sb_1__0__6_chany_top_out[12] ,
    \sb_1__0__6_chany_top_out[13] ,
    \sb_1__0__6_chany_top_out[14] ,
    \sb_1__0__6_chany_top_out[15] ,
    \sb_1__0__6_chany_top_out[16] ,
    \sb_1__0__6_chany_top_out[17] ,
    \sb_1__0__6_chany_top_out[18] ,
    \sb_1__0__6_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__48_chany_bottom_out[0] ,
    \cby_1__1__48_chany_bottom_out[1] ,
    \cby_1__1__48_chany_bottom_out[2] ,
    \cby_1__1__48_chany_bottom_out[3] ,
    \cby_1__1__48_chany_bottom_out[4] ,
    \cby_1__1__48_chany_bottom_out[5] ,
    \cby_1__1__48_chany_bottom_out[6] ,
    \cby_1__1__48_chany_bottom_out[7] ,
    \cby_1__1__48_chany_bottom_out[8] ,
    \cby_1__1__48_chany_bottom_out[9] ,
    \cby_1__1__48_chany_bottom_out[10] ,
    \cby_1__1__48_chany_bottom_out[11] ,
    \cby_1__1__48_chany_bottom_out[12] ,
    \cby_1__1__48_chany_bottom_out[13] ,
    \cby_1__1__48_chany_bottom_out[14] ,
    \cby_1__1__48_chany_bottom_out[15] ,
    \cby_1__1__48_chany_bottom_out[16] ,
    \cby_1__1__48_chany_bottom_out[17] ,
    \cby_1__1__48_chany_bottom_out[18] ,
    \cby_1__1__48_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__42_chany_bottom_out[0] ,
    \sb_1__1__42_chany_bottom_out[1] ,
    \sb_1__1__42_chany_bottom_out[2] ,
    \sb_1__1__42_chany_bottom_out[3] ,
    \sb_1__1__42_chany_bottom_out[4] ,
    \sb_1__1__42_chany_bottom_out[5] ,
    \sb_1__1__42_chany_bottom_out[6] ,
    \sb_1__1__42_chany_bottom_out[7] ,
    \sb_1__1__42_chany_bottom_out[8] ,
    \sb_1__1__42_chany_bottom_out[9] ,
    \sb_1__1__42_chany_bottom_out[10] ,
    \sb_1__1__42_chany_bottom_out[11] ,
    \sb_1__1__42_chany_bottom_out[12] ,
    \sb_1__1__42_chany_bottom_out[13] ,
    \sb_1__1__42_chany_bottom_out[14] ,
    \sb_1__1__42_chany_bottom_out[15] ,
    \sb_1__1__42_chany_bottom_out[16] ,
    \sb_1__1__42_chany_bottom_out[17] ,
    \sb_1__1__42_chany_bottom_out[18] ,
    \sb_1__1__42_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__48_chany_top_out[0] ,
    \cby_1__1__48_chany_top_out[1] ,
    \cby_1__1__48_chany_top_out[2] ,
    \cby_1__1__48_chany_top_out[3] ,
    \cby_1__1__48_chany_top_out[4] ,
    \cby_1__1__48_chany_top_out[5] ,
    \cby_1__1__48_chany_top_out[6] ,
    \cby_1__1__48_chany_top_out[7] ,
    \cby_1__1__48_chany_top_out[8] ,
    \cby_1__1__48_chany_top_out[9] ,
    \cby_1__1__48_chany_top_out[10] ,
    \cby_1__1__48_chany_top_out[11] ,
    \cby_1__1__48_chany_top_out[12] ,
    \cby_1__1__48_chany_top_out[13] ,
    \cby_1__1__48_chany_top_out[14] ,
    \cby_1__1__48_chany_top_out[15] ,
    \cby_1__1__48_chany_top_out[16] ,
    \cby_1__1__48_chany_top_out[17] ,
    \cby_1__1__48_chany_top_out[18] ,
    \cby_1__1__48_chany_top_out[19] }));
 cby_1__1_ cby_7__2_ (.Test_en_E_in(\Test_enWires[42] ),
    .Test_en_E_out(\Test_enWires[43] ),
    .Test_en_S_in(\Test_enWires[42] ),
    .Test_en_W_in(\Test_enWires[42] ),
    .ccff_head(grid_clb_49_ccff_tail),
    .ccff_tail(cby_1__1__49_ccff_tail),
    .clk_2_S_in(\clk_2_wires[37] ),
    .clk_2_S_out(\clk_2_wires[38] ),
    .left_grid_pin_16_(cby_1__1__49_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__49_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__49_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__49_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__49_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__49_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__49_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__49_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__49_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__49_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__49_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__49_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__49_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__49_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__49_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__49_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[178] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[177] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[37] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[38] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__42_chany_top_out[0] ,
    \sb_1__1__42_chany_top_out[1] ,
    \sb_1__1__42_chany_top_out[2] ,
    \sb_1__1__42_chany_top_out[3] ,
    \sb_1__1__42_chany_top_out[4] ,
    \sb_1__1__42_chany_top_out[5] ,
    \sb_1__1__42_chany_top_out[6] ,
    \sb_1__1__42_chany_top_out[7] ,
    \sb_1__1__42_chany_top_out[8] ,
    \sb_1__1__42_chany_top_out[9] ,
    \sb_1__1__42_chany_top_out[10] ,
    \sb_1__1__42_chany_top_out[11] ,
    \sb_1__1__42_chany_top_out[12] ,
    \sb_1__1__42_chany_top_out[13] ,
    \sb_1__1__42_chany_top_out[14] ,
    \sb_1__1__42_chany_top_out[15] ,
    \sb_1__1__42_chany_top_out[16] ,
    \sb_1__1__42_chany_top_out[17] ,
    \sb_1__1__42_chany_top_out[18] ,
    \sb_1__1__42_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__49_chany_bottom_out[0] ,
    \cby_1__1__49_chany_bottom_out[1] ,
    \cby_1__1__49_chany_bottom_out[2] ,
    \cby_1__1__49_chany_bottom_out[3] ,
    \cby_1__1__49_chany_bottom_out[4] ,
    \cby_1__1__49_chany_bottom_out[5] ,
    \cby_1__1__49_chany_bottom_out[6] ,
    \cby_1__1__49_chany_bottom_out[7] ,
    \cby_1__1__49_chany_bottom_out[8] ,
    \cby_1__1__49_chany_bottom_out[9] ,
    \cby_1__1__49_chany_bottom_out[10] ,
    \cby_1__1__49_chany_bottom_out[11] ,
    \cby_1__1__49_chany_bottom_out[12] ,
    \cby_1__1__49_chany_bottom_out[13] ,
    \cby_1__1__49_chany_bottom_out[14] ,
    \cby_1__1__49_chany_bottom_out[15] ,
    \cby_1__1__49_chany_bottom_out[16] ,
    \cby_1__1__49_chany_bottom_out[17] ,
    \cby_1__1__49_chany_bottom_out[18] ,
    \cby_1__1__49_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__43_chany_bottom_out[0] ,
    \sb_1__1__43_chany_bottom_out[1] ,
    \sb_1__1__43_chany_bottom_out[2] ,
    \sb_1__1__43_chany_bottom_out[3] ,
    \sb_1__1__43_chany_bottom_out[4] ,
    \sb_1__1__43_chany_bottom_out[5] ,
    \sb_1__1__43_chany_bottom_out[6] ,
    \sb_1__1__43_chany_bottom_out[7] ,
    \sb_1__1__43_chany_bottom_out[8] ,
    \sb_1__1__43_chany_bottom_out[9] ,
    \sb_1__1__43_chany_bottom_out[10] ,
    \sb_1__1__43_chany_bottom_out[11] ,
    \sb_1__1__43_chany_bottom_out[12] ,
    \sb_1__1__43_chany_bottom_out[13] ,
    \sb_1__1__43_chany_bottom_out[14] ,
    \sb_1__1__43_chany_bottom_out[15] ,
    \sb_1__1__43_chany_bottom_out[16] ,
    \sb_1__1__43_chany_bottom_out[17] ,
    \sb_1__1__43_chany_bottom_out[18] ,
    \sb_1__1__43_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__49_chany_top_out[0] ,
    \cby_1__1__49_chany_top_out[1] ,
    \cby_1__1__49_chany_top_out[2] ,
    \cby_1__1__49_chany_top_out[3] ,
    \cby_1__1__49_chany_top_out[4] ,
    \cby_1__1__49_chany_top_out[5] ,
    \cby_1__1__49_chany_top_out[6] ,
    \cby_1__1__49_chany_top_out[7] ,
    \cby_1__1__49_chany_top_out[8] ,
    \cby_1__1__49_chany_top_out[9] ,
    \cby_1__1__49_chany_top_out[10] ,
    \cby_1__1__49_chany_top_out[11] ,
    \cby_1__1__49_chany_top_out[12] ,
    \cby_1__1__49_chany_top_out[13] ,
    \cby_1__1__49_chany_top_out[14] ,
    \cby_1__1__49_chany_top_out[15] ,
    \cby_1__1__49_chany_top_out[16] ,
    \cby_1__1__49_chany_top_out[17] ,
    \cby_1__1__49_chany_top_out[18] ,
    \cby_1__1__49_chany_top_out[19] }));
 cby_1__1_ cby_7__3_ (.Test_en_E_in(\Test_enWires[56] ),
    .Test_en_E_out(\Test_enWires[57] ),
    .Test_en_S_in(\Test_enWires[56] ),
    .Test_en_W_in(\Test_enWires[56] ),
    .ccff_head(grid_clb_50_ccff_tail),
    .ccff_tail(cby_1__1__50_ccff_tail),
    .clk_2_N_out(\clk_2_wires[36] ),
    .clk_2_S_in(\clk_2_wires[35] ),
    .left_grid_pin_16_(cby_1__1__50_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__50_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__50_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__50_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__50_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__50_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__50_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__50_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__50_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__50_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__50_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__50_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__50_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__50_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__50_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__50_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[181] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[180] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[36] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[35] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__43_chany_top_out[0] ,
    \sb_1__1__43_chany_top_out[1] ,
    \sb_1__1__43_chany_top_out[2] ,
    \sb_1__1__43_chany_top_out[3] ,
    \sb_1__1__43_chany_top_out[4] ,
    \sb_1__1__43_chany_top_out[5] ,
    \sb_1__1__43_chany_top_out[6] ,
    \sb_1__1__43_chany_top_out[7] ,
    \sb_1__1__43_chany_top_out[8] ,
    \sb_1__1__43_chany_top_out[9] ,
    \sb_1__1__43_chany_top_out[10] ,
    \sb_1__1__43_chany_top_out[11] ,
    \sb_1__1__43_chany_top_out[12] ,
    \sb_1__1__43_chany_top_out[13] ,
    \sb_1__1__43_chany_top_out[14] ,
    \sb_1__1__43_chany_top_out[15] ,
    \sb_1__1__43_chany_top_out[16] ,
    \sb_1__1__43_chany_top_out[17] ,
    \sb_1__1__43_chany_top_out[18] ,
    \sb_1__1__43_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__50_chany_bottom_out[0] ,
    \cby_1__1__50_chany_bottom_out[1] ,
    \cby_1__1__50_chany_bottom_out[2] ,
    \cby_1__1__50_chany_bottom_out[3] ,
    \cby_1__1__50_chany_bottom_out[4] ,
    \cby_1__1__50_chany_bottom_out[5] ,
    \cby_1__1__50_chany_bottom_out[6] ,
    \cby_1__1__50_chany_bottom_out[7] ,
    \cby_1__1__50_chany_bottom_out[8] ,
    \cby_1__1__50_chany_bottom_out[9] ,
    \cby_1__1__50_chany_bottom_out[10] ,
    \cby_1__1__50_chany_bottom_out[11] ,
    \cby_1__1__50_chany_bottom_out[12] ,
    \cby_1__1__50_chany_bottom_out[13] ,
    \cby_1__1__50_chany_bottom_out[14] ,
    \cby_1__1__50_chany_bottom_out[15] ,
    \cby_1__1__50_chany_bottom_out[16] ,
    \cby_1__1__50_chany_bottom_out[17] ,
    \cby_1__1__50_chany_bottom_out[18] ,
    \cby_1__1__50_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__44_chany_bottom_out[0] ,
    \sb_1__1__44_chany_bottom_out[1] ,
    \sb_1__1__44_chany_bottom_out[2] ,
    \sb_1__1__44_chany_bottom_out[3] ,
    \sb_1__1__44_chany_bottom_out[4] ,
    \sb_1__1__44_chany_bottom_out[5] ,
    \sb_1__1__44_chany_bottom_out[6] ,
    \sb_1__1__44_chany_bottom_out[7] ,
    \sb_1__1__44_chany_bottom_out[8] ,
    \sb_1__1__44_chany_bottom_out[9] ,
    \sb_1__1__44_chany_bottom_out[10] ,
    \sb_1__1__44_chany_bottom_out[11] ,
    \sb_1__1__44_chany_bottom_out[12] ,
    \sb_1__1__44_chany_bottom_out[13] ,
    \sb_1__1__44_chany_bottom_out[14] ,
    \sb_1__1__44_chany_bottom_out[15] ,
    \sb_1__1__44_chany_bottom_out[16] ,
    \sb_1__1__44_chany_bottom_out[17] ,
    \sb_1__1__44_chany_bottom_out[18] ,
    \sb_1__1__44_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__50_chany_top_out[0] ,
    \cby_1__1__50_chany_top_out[1] ,
    \cby_1__1__50_chany_top_out[2] ,
    \cby_1__1__50_chany_top_out[3] ,
    \cby_1__1__50_chany_top_out[4] ,
    \cby_1__1__50_chany_top_out[5] ,
    \cby_1__1__50_chany_top_out[6] ,
    \cby_1__1__50_chany_top_out[7] ,
    \cby_1__1__50_chany_top_out[8] ,
    \cby_1__1__50_chany_top_out[9] ,
    \cby_1__1__50_chany_top_out[10] ,
    \cby_1__1__50_chany_top_out[11] ,
    \cby_1__1__50_chany_top_out[12] ,
    \cby_1__1__50_chany_top_out[13] ,
    \cby_1__1__50_chany_top_out[14] ,
    \cby_1__1__50_chany_top_out[15] ,
    \cby_1__1__50_chany_top_out[16] ,
    \cby_1__1__50_chany_top_out[17] ,
    \cby_1__1__50_chany_top_out[18] ,
    \cby_1__1__50_chany_top_out[19] }));
 cby_1__1_ cby_7__4_ (.Test_en_E_in(\Test_enWires[70] ),
    .Test_en_E_out(\Test_enWires[71] ),
    .Test_en_S_in(\Test_enWires[70] ),
    .Test_en_W_in(\Test_enWires[70] ),
    .ccff_head(grid_clb_51_ccff_tail),
    .ccff_tail(cby_1__1__51_ccff_tail),
    .left_grid_pin_16_(cby_1__1__51_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__51_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__51_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__51_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__51_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__51_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__51_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__51_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__51_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__51_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__51_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__51_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__51_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__51_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__51_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__51_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[184] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[183] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__44_chany_top_out[0] ,
    \sb_1__1__44_chany_top_out[1] ,
    \sb_1__1__44_chany_top_out[2] ,
    \sb_1__1__44_chany_top_out[3] ,
    \sb_1__1__44_chany_top_out[4] ,
    \sb_1__1__44_chany_top_out[5] ,
    \sb_1__1__44_chany_top_out[6] ,
    \sb_1__1__44_chany_top_out[7] ,
    \sb_1__1__44_chany_top_out[8] ,
    \sb_1__1__44_chany_top_out[9] ,
    \sb_1__1__44_chany_top_out[10] ,
    \sb_1__1__44_chany_top_out[11] ,
    \sb_1__1__44_chany_top_out[12] ,
    \sb_1__1__44_chany_top_out[13] ,
    \sb_1__1__44_chany_top_out[14] ,
    \sb_1__1__44_chany_top_out[15] ,
    \sb_1__1__44_chany_top_out[16] ,
    \sb_1__1__44_chany_top_out[17] ,
    \sb_1__1__44_chany_top_out[18] ,
    \sb_1__1__44_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__51_chany_bottom_out[0] ,
    \cby_1__1__51_chany_bottom_out[1] ,
    \cby_1__1__51_chany_bottom_out[2] ,
    \cby_1__1__51_chany_bottom_out[3] ,
    \cby_1__1__51_chany_bottom_out[4] ,
    \cby_1__1__51_chany_bottom_out[5] ,
    \cby_1__1__51_chany_bottom_out[6] ,
    \cby_1__1__51_chany_bottom_out[7] ,
    \cby_1__1__51_chany_bottom_out[8] ,
    \cby_1__1__51_chany_bottom_out[9] ,
    \cby_1__1__51_chany_bottom_out[10] ,
    \cby_1__1__51_chany_bottom_out[11] ,
    \cby_1__1__51_chany_bottom_out[12] ,
    \cby_1__1__51_chany_bottom_out[13] ,
    \cby_1__1__51_chany_bottom_out[14] ,
    \cby_1__1__51_chany_bottom_out[15] ,
    \cby_1__1__51_chany_bottom_out[16] ,
    \cby_1__1__51_chany_bottom_out[17] ,
    \cby_1__1__51_chany_bottom_out[18] ,
    \cby_1__1__51_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__45_chany_bottom_out[0] ,
    \sb_1__1__45_chany_bottom_out[1] ,
    \sb_1__1__45_chany_bottom_out[2] ,
    \sb_1__1__45_chany_bottom_out[3] ,
    \sb_1__1__45_chany_bottom_out[4] ,
    \sb_1__1__45_chany_bottom_out[5] ,
    \sb_1__1__45_chany_bottom_out[6] ,
    \sb_1__1__45_chany_bottom_out[7] ,
    \sb_1__1__45_chany_bottom_out[8] ,
    \sb_1__1__45_chany_bottom_out[9] ,
    \sb_1__1__45_chany_bottom_out[10] ,
    \sb_1__1__45_chany_bottom_out[11] ,
    \sb_1__1__45_chany_bottom_out[12] ,
    \sb_1__1__45_chany_bottom_out[13] ,
    \sb_1__1__45_chany_bottom_out[14] ,
    \sb_1__1__45_chany_bottom_out[15] ,
    \sb_1__1__45_chany_bottom_out[16] ,
    \sb_1__1__45_chany_bottom_out[17] ,
    \sb_1__1__45_chany_bottom_out[18] ,
    \sb_1__1__45_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__51_chany_top_out[0] ,
    \cby_1__1__51_chany_top_out[1] ,
    \cby_1__1__51_chany_top_out[2] ,
    \cby_1__1__51_chany_top_out[3] ,
    \cby_1__1__51_chany_top_out[4] ,
    \cby_1__1__51_chany_top_out[5] ,
    \cby_1__1__51_chany_top_out[6] ,
    \cby_1__1__51_chany_top_out[7] ,
    \cby_1__1__51_chany_top_out[8] ,
    \cby_1__1__51_chany_top_out[9] ,
    \cby_1__1__51_chany_top_out[10] ,
    \cby_1__1__51_chany_top_out[11] ,
    \cby_1__1__51_chany_top_out[12] ,
    \cby_1__1__51_chany_top_out[13] ,
    \cby_1__1__51_chany_top_out[14] ,
    \cby_1__1__51_chany_top_out[15] ,
    \cby_1__1__51_chany_top_out[16] ,
    \cby_1__1__51_chany_top_out[17] ,
    \cby_1__1__51_chany_top_out[18] ,
    \cby_1__1__51_chany_top_out[19] }));
 cby_1__1_ cby_7__5_ (.Test_en_E_in(\Test_enWires[84] ),
    .Test_en_E_out(\Test_enWires[85] ),
    .Test_en_S_in(\Test_enWires[84] ),
    .Test_en_W_in(\Test_enWires[84] ),
    .ccff_head(grid_clb_52_ccff_tail),
    .ccff_tail(cby_1__1__52_ccff_tail),
    .left_grid_pin_16_(cby_1__1__52_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__52_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__52_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__52_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__52_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__52_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__52_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__52_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__52_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__52_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__52_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__52_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__52_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__52_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__52_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__52_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[187] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[186] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__45_chany_top_out[0] ,
    \sb_1__1__45_chany_top_out[1] ,
    \sb_1__1__45_chany_top_out[2] ,
    \sb_1__1__45_chany_top_out[3] ,
    \sb_1__1__45_chany_top_out[4] ,
    \sb_1__1__45_chany_top_out[5] ,
    \sb_1__1__45_chany_top_out[6] ,
    \sb_1__1__45_chany_top_out[7] ,
    \sb_1__1__45_chany_top_out[8] ,
    \sb_1__1__45_chany_top_out[9] ,
    \sb_1__1__45_chany_top_out[10] ,
    \sb_1__1__45_chany_top_out[11] ,
    \sb_1__1__45_chany_top_out[12] ,
    \sb_1__1__45_chany_top_out[13] ,
    \sb_1__1__45_chany_top_out[14] ,
    \sb_1__1__45_chany_top_out[15] ,
    \sb_1__1__45_chany_top_out[16] ,
    \sb_1__1__45_chany_top_out[17] ,
    \sb_1__1__45_chany_top_out[18] ,
    \sb_1__1__45_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__52_chany_bottom_out[0] ,
    \cby_1__1__52_chany_bottom_out[1] ,
    \cby_1__1__52_chany_bottom_out[2] ,
    \cby_1__1__52_chany_bottom_out[3] ,
    \cby_1__1__52_chany_bottom_out[4] ,
    \cby_1__1__52_chany_bottom_out[5] ,
    \cby_1__1__52_chany_bottom_out[6] ,
    \cby_1__1__52_chany_bottom_out[7] ,
    \cby_1__1__52_chany_bottom_out[8] ,
    \cby_1__1__52_chany_bottom_out[9] ,
    \cby_1__1__52_chany_bottom_out[10] ,
    \cby_1__1__52_chany_bottom_out[11] ,
    \cby_1__1__52_chany_bottom_out[12] ,
    \cby_1__1__52_chany_bottom_out[13] ,
    \cby_1__1__52_chany_bottom_out[14] ,
    \cby_1__1__52_chany_bottom_out[15] ,
    \cby_1__1__52_chany_bottom_out[16] ,
    \cby_1__1__52_chany_bottom_out[17] ,
    \cby_1__1__52_chany_bottom_out[18] ,
    \cby_1__1__52_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__46_chany_bottom_out[0] ,
    \sb_1__1__46_chany_bottom_out[1] ,
    \sb_1__1__46_chany_bottom_out[2] ,
    \sb_1__1__46_chany_bottom_out[3] ,
    \sb_1__1__46_chany_bottom_out[4] ,
    \sb_1__1__46_chany_bottom_out[5] ,
    \sb_1__1__46_chany_bottom_out[6] ,
    \sb_1__1__46_chany_bottom_out[7] ,
    \sb_1__1__46_chany_bottom_out[8] ,
    \sb_1__1__46_chany_bottom_out[9] ,
    \sb_1__1__46_chany_bottom_out[10] ,
    \sb_1__1__46_chany_bottom_out[11] ,
    \sb_1__1__46_chany_bottom_out[12] ,
    \sb_1__1__46_chany_bottom_out[13] ,
    \sb_1__1__46_chany_bottom_out[14] ,
    \sb_1__1__46_chany_bottom_out[15] ,
    \sb_1__1__46_chany_bottom_out[16] ,
    \sb_1__1__46_chany_bottom_out[17] ,
    \sb_1__1__46_chany_bottom_out[18] ,
    \sb_1__1__46_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__52_chany_top_out[0] ,
    \cby_1__1__52_chany_top_out[1] ,
    \cby_1__1__52_chany_top_out[2] ,
    \cby_1__1__52_chany_top_out[3] ,
    \cby_1__1__52_chany_top_out[4] ,
    \cby_1__1__52_chany_top_out[5] ,
    \cby_1__1__52_chany_top_out[6] ,
    \cby_1__1__52_chany_top_out[7] ,
    \cby_1__1__52_chany_top_out[8] ,
    \cby_1__1__52_chany_top_out[9] ,
    \cby_1__1__52_chany_top_out[10] ,
    \cby_1__1__52_chany_top_out[11] ,
    \cby_1__1__52_chany_top_out[12] ,
    \cby_1__1__52_chany_top_out[13] ,
    \cby_1__1__52_chany_top_out[14] ,
    \cby_1__1__52_chany_top_out[15] ,
    \cby_1__1__52_chany_top_out[16] ,
    \cby_1__1__52_chany_top_out[17] ,
    \cby_1__1__52_chany_top_out[18] ,
    \cby_1__1__52_chany_top_out[19] }));
 cby_1__1_ cby_7__6_ (.Test_en_E_in(\Test_enWires[98] ),
    .Test_en_E_out(\Test_enWires[99] ),
    .Test_en_S_in(\Test_enWires[98] ),
    .Test_en_W_in(\Test_enWires[98] ),
    .ccff_head(grid_clb_53_ccff_tail),
    .ccff_tail(cby_1__1__53_ccff_tail),
    .clk_2_S_in(\clk_2_wires[50] ),
    .clk_2_S_out(\clk_2_wires[51] ),
    .left_grid_pin_16_(cby_1__1__53_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__53_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__53_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__53_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__53_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__53_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__53_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__53_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__53_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__53_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__53_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__53_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__53_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__53_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__53_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__53_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[190] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[189] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[50] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[51] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__46_chany_top_out[0] ,
    \sb_1__1__46_chany_top_out[1] ,
    \sb_1__1__46_chany_top_out[2] ,
    \sb_1__1__46_chany_top_out[3] ,
    \sb_1__1__46_chany_top_out[4] ,
    \sb_1__1__46_chany_top_out[5] ,
    \sb_1__1__46_chany_top_out[6] ,
    \sb_1__1__46_chany_top_out[7] ,
    \sb_1__1__46_chany_top_out[8] ,
    \sb_1__1__46_chany_top_out[9] ,
    \sb_1__1__46_chany_top_out[10] ,
    \sb_1__1__46_chany_top_out[11] ,
    \sb_1__1__46_chany_top_out[12] ,
    \sb_1__1__46_chany_top_out[13] ,
    \sb_1__1__46_chany_top_out[14] ,
    \sb_1__1__46_chany_top_out[15] ,
    \sb_1__1__46_chany_top_out[16] ,
    \sb_1__1__46_chany_top_out[17] ,
    \sb_1__1__46_chany_top_out[18] ,
    \sb_1__1__46_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__53_chany_bottom_out[0] ,
    \cby_1__1__53_chany_bottom_out[1] ,
    \cby_1__1__53_chany_bottom_out[2] ,
    \cby_1__1__53_chany_bottom_out[3] ,
    \cby_1__1__53_chany_bottom_out[4] ,
    \cby_1__1__53_chany_bottom_out[5] ,
    \cby_1__1__53_chany_bottom_out[6] ,
    \cby_1__1__53_chany_bottom_out[7] ,
    \cby_1__1__53_chany_bottom_out[8] ,
    \cby_1__1__53_chany_bottom_out[9] ,
    \cby_1__1__53_chany_bottom_out[10] ,
    \cby_1__1__53_chany_bottom_out[11] ,
    \cby_1__1__53_chany_bottom_out[12] ,
    \cby_1__1__53_chany_bottom_out[13] ,
    \cby_1__1__53_chany_bottom_out[14] ,
    \cby_1__1__53_chany_bottom_out[15] ,
    \cby_1__1__53_chany_bottom_out[16] ,
    \cby_1__1__53_chany_bottom_out[17] ,
    \cby_1__1__53_chany_bottom_out[18] ,
    \cby_1__1__53_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__47_chany_bottom_out[0] ,
    \sb_1__1__47_chany_bottom_out[1] ,
    \sb_1__1__47_chany_bottom_out[2] ,
    \sb_1__1__47_chany_bottom_out[3] ,
    \sb_1__1__47_chany_bottom_out[4] ,
    \sb_1__1__47_chany_bottom_out[5] ,
    \sb_1__1__47_chany_bottom_out[6] ,
    \sb_1__1__47_chany_bottom_out[7] ,
    \sb_1__1__47_chany_bottom_out[8] ,
    \sb_1__1__47_chany_bottom_out[9] ,
    \sb_1__1__47_chany_bottom_out[10] ,
    \sb_1__1__47_chany_bottom_out[11] ,
    \sb_1__1__47_chany_bottom_out[12] ,
    \sb_1__1__47_chany_bottom_out[13] ,
    \sb_1__1__47_chany_bottom_out[14] ,
    \sb_1__1__47_chany_bottom_out[15] ,
    \sb_1__1__47_chany_bottom_out[16] ,
    \sb_1__1__47_chany_bottom_out[17] ,
    \sb_1__1__47_chany_bottom_out[18] ,
    \sb_1__1__47_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__53_chany_top_out[0] ,
    \cby_1__1__53_chany_top_out[1] ,
    \cby_1__1__53_chany_top_out[2] ,
    \cby_1__1__53_chany_top_out[3] ,
    \cby_1__1__53_chany_top_out[4] ,
    \cby_1__1__53_chany_top_out[5] ,
    \cby_1__1__53_chany_top_out[6] ,
    \cby_1__1__53_chany_top_out[7] ,
    \cby_1__1__53_chany_top_out[8] ,
    \cby_1__1__53_chany_top_out[9] ,
    \cby_1__1__53_chany_top_out[10] ,
    \cby_1__1__53_chany_top_out[11] ,
    \cby_1__1__53_chany_top_out[12] ,
    \cby_1__1__53_chany_top_out[13] ,
    \cby_1__1__53_chany_top_out[14] ,
    \cby_1__1__53_chany_top_out[15] ,
    \cby_1__1__53_chany_top_out[16] ,
    \cby_1__1__53_chany_top_out[17] ,
    \cby_1__1__53_chany_top_out[18] ,
    \cby_1__1__53_chany_top_out[19] }));
 cby_1__1_ cby_7__7_ (.Test_en_E_in(\Test_enWires[112] ),
    .Test_en_E_out(\Test_enWires[113] ),
    .Test_en_S_in(\Test_enWires[112] ),
    .Test_en_W_in(\Test_enWires[112] ),
    .ccff_head(grid_clb_54_ccff_tail),
    .ccff_tail(cby_1__1__54_ccff_tail),
    .clk_2_N_out(\clk_2_wires[49] ),
    .clk_2_S_in(\clk_2_wires[48] ),
    .left_grid_pin_16_(cby_1__1__54_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__54_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__54_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__54_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__54_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__54_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__54_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__54_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__54_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__54_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__54_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__54_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__54_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__54_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__54_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__54_left_grid_pin_31_),
    .prog_clk_0_S_out(\prog_clk_0_wires[193] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[192] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[49] ),
    .prog_clk_2_S_in(\prog_clk_2_wires[48] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__47_chany_top_out[0] ,
    \sb_1__1__47_chany_top_out[1] ,
    \sb_1__1__47_chany_top_out[2] ,
    \sb_1__1__47_chany_top_out[3] ,
    \sb_1__1__47_chany_top_out[4] ,
    \sb_1__1__47_chany_top_out[5] ,
    \sb_1__1__47_chany_top_out[6] ,
    \sb_1__1__47_chany_top_out[7] ,
    \sb_1__1__47_chany_top_out[8] ,
    \sb_1__1__47_chany_top_out[9] ,
    \sb_1__1__47_chany_top_out[10] ,
    \sb_1__1__47_chany_top_out[11] ,
    \sb_1__1__47_chany_top_out[12] ,
    \sb_1__1__47_chany_top_out[13] ,
    \sb_1__1__47_chany_top_out[14] ,
    \sb_1__1__47_chany_top_out[15] ,
    \sb_1__1__47_chany_top_out[16] ,
    \sb_1__1__47_chany_top_out[17] ,
    \sb_1__1__47_chany_top_out[18] ,
    \sb_1__1__47_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__54_chany_bottom_out[0] ,
    \cby_1__1__54_chany_bottom_out[1] ,
    \cby_1__1__54_chany_bottom_out[2] ,
    \cby_1__1__54_chany_bottom_out[3] ,
    \cby_1__1__54_chany_bottom_out[4] ,
    \cby_1__1__54_chany_bottom_out[5] ,
    \cby_1__1__54_chany_bottom_out[6] ,
    \cby_1__1__54_chany_bottom_out[7] ,
    \cby_1__1__54_chany_bottom_out[8] ,
    \cby_1__1__54_chany_bottom_out[9] ,
    \cby_1__1__54_chany_bottom_out[10] ,
    \cby_1__1__54_chany_bottom_out[11] ,
    \cby_1__1__54_chany_bottom_out[12] ,
    \cby_1__1__54_chany_bottom_out[13] ,
    \cby_1__1__54_chany_bottom_out[14] ,
    \cby_1__1__54_chany_bottom_out[15] ,
    \cby_1__1__54_chany_bottom_out[16] ,
    \cby_1__1__54_chany_bottom_out[17] ,
    \cby_1__1__54_chany_bottom_out[18] ,
    \cby_1__1__54_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__1__48_chany_bottom_out[0] ,
    \sb_1__1__48_chany_bottom_out[1] ,
    \sb_1__1__48_chany_bottom_out[2] ,
    \sb_1__1__48_chany_bottom_out[3] ,
    \sb_1__1__48_chany_bottom_out[4] ,
    \sb_1__1__48_chany_bottom_out[5] ,
    \sb_1__1__48_chany_bottom_out[6] ,
    \sb_1__1__48_chany_bottom_out[7] ,
    \sb_1__1__48_chany_bottom_out[8] ,
    \sb_1__1__48_chany_bottom_out[9] ,
    \sb_1__1__48_chany_bottom_out[10] ,
    \sb_1__1__48_chany_bottom_out[11] ,
    \sb_1__1__48_chany_bottom_out[12] ,
    \sb_1__1__48_chany_bottom_out[13] ,
    \sb_1__1__48_chany_bottom_out[14] ,
    \sb_1__1__48_chany_bottom_out[15] ,
    \sb_1__1__48_chany_bottom_out[16] ,
    \sb_1__1__48_chany_bottom_out[17] ,
    \sb_1__1__48_chany_bottom_out[18] ,
    \sb_1__1__48_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__54_chany_top_out[0] ,
    \cby_1__1__54_chany_top_out[1] ,
    \cby_1__1__54_chany_top_out[2] ,
    \cby_1__1__54_chany_top_out[3] ,
    \cby_1__1__54_chany_top_out[4] ,
    \cby_1__1__54_chany_top_out[5] ,
    \cby_1__1__54_chany_top_out[6] ,
    \cby_1__1__54_chany_top_out[7] ,
    \cby_1__1__54_chany_top_out[8] ,
    \cby_1__1__54_chany_top_out[9] ,
    \cby_1__1__54_chany_top_out[10] ,
    \cby_1__1__54_chany_top_out[11] ,
    \cby_1__1__54_chany_top_out[12] ,
    \cby_1__1__54_chany_top_out[13] ,
    \cby_1__1__54_chany_top_out[14] ,
    \cby_1__1__54_chany_top_out[15] ,
    \cby_1__1__54_chany_top_out[16] ,
    \cby_1__1__54_chany_top_out[17] ,
    \cby_1__1__54_chany_top_out[18] ,
    \cby_1__1__54_chany_top_out[19] }));
 cby_1__1_ cby_7__8_ (.Test_en_E_in(\Test_enWires[126] ),
    .Test_en_E_out(\Test_enWires[127] ),
    .Test_en_S_in(\Test_enWires[126] ),
    .Test_en_W_in(\Test_enWires[126] ),
    .ccff_head(grid_clb_55_ccff_tail),
    .ccff_tail(cby_1__1__55_ccff_tail),
    .left_grid_pin_16_(cby_1__1__55_left_grid_pin_16_),
    .left_grid_pin_17_(cby_1__1__55_left_grid_pin_17_),
    .left_grid_pin_18_(cby_1__1__55_left_grid_pin_18_),
    .left_grid_pin_19_(cby_1__1__55_left_grid_pin_19_),
    .left_grid_pin_20_(cby_1__1__55_left_grid_pin_20_),
    .left_grid_pin_21_(cby_1__1__55_left_grid_pin_21_),
    .left_grid_pin_22_(cby_1__1__55_left_grid_pin_22_),
    .left_grid_pin_23_(cby_1__1__55_left_grid_pin_23_),
    .left_grid_pin_24_(cby_1__1__55_left_grid_pin_24_),
    .left_grid_pin_25_(cby_1__1__55_left_grid_pin_25_),
    .left_grid_pin_26_(cby_1__1__55_left_grid_pin_26_),
    .left_grid_pin_27_(cby_1__1__55_left_grid_pin_27_),
    .left_grid_pin_28_(cby_1__1__55_left_grid_pin_28_),
    .left_grid_pin_29_(cby_1__1__55_left_grid_pin_29_),
    .left_grid_pin_30_(cby_1__1__55_left_grid_pin_30_),
    .left_grid_pin_31_(cby_1__1__55_left_grid_pin_31_),
    .prog_clk_0_N_out(\prog_clk_0_wires[198] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[196] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[195] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_1__1__48_chany_top_out[0] ,
    \sb_1__1__48_chany_top_out[1] ,
    \sb_1__1__48_chany_top_out[2] ,
    \sb_1__1__48_chany_top_out[3] ,
    \sb_1__1__48_chany_top_out[4] ,
    \sb_1__1__48_chany_top_out[5] ,
    \sb_1__1__48_chany_top_out[6] ,
    \sb_1__1__48_chany_top_out[7] ,
    \sb_1__1__48_chany_top_out[8] ,
    \sb_1__1__48_chany_top_out[9] ,
    \sb_1__1__48_chany_top_out[10] ,
    \sb_1__1__48_chany_top_out[11] ,
    \sb_1__1__48_chany_top_out[12] ,
    \sb_1__1__48_chany_top_out[13] ,
    \sb_1__1__48_chany_top_out[14] ,
    \sb_1__1__48_chany_top_out[15] ,
    \sb_1__1__48_chany_top_out[16] ,
    \sb_1__1__48_chany_top_out[17] ,
    \sb_1__1__48_chany_top_out[18] ,
    \sb_1__1__48_chany_top_out[19] }),
    .chany_bottom_out({\cby_1__1__55_chany_bottom_out[0] ,
    \cby_1__1__55_chany_bottom_out[1] ,
    \cby_1__1__55_chany_bottom_out[2] ,
    \cby_1__1__55_chany_bottom_out[3] ,
    \cby_1__1__55_chany_bottom_out[4] ,
    \cby_1__1__55_chany_bottom_out[5] ,
    \cby_1__1__55_chany_bottom_out[6] ,
    \cby_1__1__55_chany_bottom_out[7] ,
    \cby_1__1__55_chany_bottom_out[8] ,
    \cby_1__1__55_chany_bottom_out[9] ,
    \cby_1__1__55_chany_bottom_out[10] ,
    \cby_1__1__55_chany_bottom_out[11] ,
    \cby_1__1__55_chany_bottom_out[12] ,
    \cby_1__1__55_chany_bottom_out[13] ,
    \cby_1__1__55_chany_bottom_out[14] ,
    \cby_1__1__55_chany_bottom_out[15] ,
    \cby_1__1__55_chany_bottom_out[16] ,
    \cby_1__1__55_chany_bottom_out[17] ,
    \cby_1__1__55_chany_bottom_out[18] ,
    \cby_1__1__55_chany_bottom_out[19] }),
    .chany_top_in({\sb_1__8__6_chany_bottom_out[0] ,
    \sb_1__8__6_chany_bottom_out[1] ,
    \sb_1__8__6_chany_bottom_out[2] ,
    \sb_1__8__6_chany_bottom_out[3] ,
    \sb_1__8__6_chany_bottom_out[4] ,
    \sb_1__8__6_chany_bottom_out[5] ,
    \sb_1__8__6_chany_bottom_out[6] ,
    \sb_1__8__6_chany_bottom_out[7] ,
    \sb_1__8__6_chany_bottom_out[8] ,
    \sb_1__8__6_chany_bottom_out[9] ,
    \sb_1__8__6_chany_bottom_out[10] ,
    \sb_1__8__6_chany_bottom_out[11] ,
    \sb_1__8__6_chany_bottom_out[12] ,
    \sb_1__8__6_chany_bottom_out[13] ,
    \sb_1__8__6_chany_bottom_out[14] ,
    \sb_1__8__6_chany_bottom_out[15] ,
    \sb_1__8__6_chany_bottom_out[16] ,
    \sb_1__8__6_chany_bottom_out[17] ,
    \sb_1__8__6_chany_bottom_out[18] ,
    \sb_1__8__6_chany_bottom_out[19] }),
    .chany_top_out({\cby_1__1__55_chany_top_out[0] ,
    \cby_1__1__55_chany_top_out[1] ,
    \cby_1__1__55_chany_top_out[2] ,
    \cby_1__1__55_chany_top_out[3] ,
    \cby_1__1__55_chany_top_out[4] ,
    \cby_1__1__55_chany_top_out[5] ,
    \cby_1__1__55_chany_top_out[6] ,
    \cby_1__1__55_chany_top_out[7] ,
    \cby_1__1__55_chany_top_out[8] ,
    \cby_1__1__55_chany_top_out[9] ,
    \cby_1__1__55_chany_top_out[10] ,
    \cby_1__1__55_chany_top_out[11] ,
    \cby_1__1__55_chany_top_out[12] ,
    \cby_1__1__55_chany_top_out[13] ,
    \cby_1__1__55_chany_top_out[14] ,
    \cby_1__1__55_chany_top_out[15] ,
    \cby_1__1__55_chany_top_out[16] ,
    \cby_1__1__55_chany_top_out[17] ,
    \cby_1__1__55_chany_top_out[18] ,
    \cby_1__1__55_chany_top_out[19] }));
 cby_2__1_ cby_8__1_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_56_ccff_tail),
    .ccff_tail(grid_io_right_7_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]),
    .left_grid_pin_16_(cby_8__1__0_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__0_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__0_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__0_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__0_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__0_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__0_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__0_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__0_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__0_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__0_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__0_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__0_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__0_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__0_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__0_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__0_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_7_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_7_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_S_out(\prog_clk_0_wires[201] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[200] ),
    .right_grid_pin_0_(cby_8__1__0_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__0__0_chany_top_out[0] ,
    \sb_8__0__0_chany_top_out[1] ,
    \sb_8__0__0_chany_top_out[2] ,
    \sb_8__0__0_chany_top_out[3] ,
    \sb_8__0__0_chany_top_out[4] ,
    \sb_8__0__0_chany_top_out[5] ,
    \sb_8__0__0_chany_top_out[6] ,
    \sb_8__0__0_chany_top_out[7] ,
    \sb_8__0__0_chany_top_out[8] ,
    \sb_8__0__0_chany_top_out[9] ,
    \sb_8__0__0_chany_top_out[10] ,
    \sb_8__0__0_chany_top_out[11] ,
    \sb_8__0__0_chany_top_out[12] ,
    \sb_8__0__0_chany_top_out[13] ,
    \sb_8__0__0_chany_top_out[14] ,
    \sb_8__0__0_chany_top_out[15] ,
    \sb_8__0__0_chany_top_out[16] ,
    \sb_8__0__0_chany_top_out[17] ,
    \sb_8__0__0_chany_top_out[18] ,
    \sb_8__0__0_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__0_chany_bottom_out[0] ,
    \cby_8__1__0_chany_bottom_out[1] ,
    \cby_8__1__0_chany_bottom_out[2] ,
    \cby_8__1__0_chany_bottom_out[3] ,
    \cby_8__1__0_chany_bottom_out[4] ,
    \cby_8__1__0_chany_bottom_out[5] ,
    \cby_8__1__0_chany_bottom_out[6] ,
    \cby_8__1__0_chany_bottom_out[7] ,
    \cby_8__1__0_chany_bottom_out[8] ,
    \cby_8__1__0_chany_bottom_out[9] ,
    \cby_8__1__0_chany_bottom_out[10] ,
    \cby_8__1__0_chany_bottom_out[11] ,
    \cby_8__1__0_chany_bottom_out[12] ,
    \cby_8__1__0_chany_bottom_out[13] ,
    \cby_8__1__0_chany_bottom_out[14] ,
    \cby_8__1__0_chany_bottom_out[15] ,
    \cby_8__1__0_chany_bottom_out[16] ,
    \cby_8__1__0_chany_bottom_out[17] ,
    \cby_8__1__0_chany_bottom_out[18] ,
    \cby_8__1__0_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__1__0_chany_bottom_out[0] ,
    \sb_8__1__0_chany_bottom_out[1] ,
    \sb_8__1__0_chany_bottom_out[2] ,
    \sb_8__1__0_chany_bottom_out[3] ,
    \sb_8__1__0_chany_bottom_out[4] ,
    \sb_8__1__0_chany_bottom_out[5] ,
    \sb_8__1__0_chany_bottom_out[6] ,
    \sb_8__1__0_chany_bottom_out[7] ,
    \sb_8__1__0_chany_bottom_out[8] ,
    \sb_8__1__0_chany_bottom_out[9] ,
    \sb_8__1__0_chany_bottom_out[10] ,
    \sb_8__1__0_chany_bottom_out[11] ,
    \sb_8__1__0_chany_bottom_out[12] ,
    \sb_8__1__0_chany_bottom_out[13] ,
    \sb_8__1__0_chany_bottom_out[14] ,
    \sb_8__1__0_chany_bottom_out[15] ,
    \sb_8__1__0_chany_bottom_out[16] ,
    \sb_8__1__0_chany_bottom_out[17] ,
    \sb_8__1__0_chany_bottom_out[18] ,
    \sb_8__1__0_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__0_chany_top_out[0] ,
    \cby_8__1__0_chany_top_out[1] ,
    \cby_8__1__0_chany_top_out[2] ,
    \cby_8__1__0_chany_top_out[3] ,
    \cby_8__1__0_chany_top_out[4] ,
    \cby_8__1__0_chany_top_out[5] ,
    \cby_8__1__0_chany_top_out[6] ,
    \cby_8__1__0_chany_top_out[7] ,
    \cby_8__1__0_chany_top_out[8] ,
    \cby_8__1__0_chany_top_out[9] ,
    \cby_8__1__0_chany_top_out[10] ,
    \cby_8__1__0_chany_top_out[11] ,
    \cby_8__1__0_chany_top_out[12] ,
    \cby_8__1__0_chany_top_out[13] ,
    \cby_8__1__0_chany_top_out[14] ,
    \cby_8__1__0_chany_top_out[15] ,
    \cby_8__1__0_chany_top_out[16] ,
    \cby_8__1__0_chany_top_out[17] ,
    \cby_8__1__0_chany_top_out[18] ,
    \cby_8__1__0_chany_top_out[19] }));
 cby_2__1_ cby_8__2_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_57_ccff_tail),
    .ccff_tail(grid_io_right_6_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]),
    .left_grid_pin_16_(cby_8__1__1_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__1_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__1_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__1_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__1_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__1_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__1_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__1_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__1_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__1_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__1_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__1_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__1_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__1_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__1_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__1_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__1_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_6_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_6_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_S_out(\prog_clk_0_wires[204] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[203] ),
    .right_grid_pin_0_(cby_8__1__1_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__1__0_chany_top_out[0] ,
    \sb_8__1__0_chany_top_out[1] ,
    \sb_8__1__0_chany_top_out[2] ,
    \sb_8__1__0_chany_top_out[3] ,
    \sb_8__1__0_chany_top_out[4] ,
    \sb_8__1__0_chany_top_out[5] ,
    \sb_8__1__0_chany_top_out[6] ,
    \sb_8__1__0_chany_top_out[7] ,
    \sb_8__1__0_chany_top_out[8] ,
    \sb_8__1__0_chany_top_out[9] ,
    \sb_8__1__0_chany_top_out[10] ,
    \sb_8__1__0_chany_top_out[11] ,
    \sb_8__1__0_chany_top_out[12] ,
    \sb_8__1__0_chany_top_out[13] ,
    \sb_8__1__0_chany_top_out[14] ,
    \sb_8__1__0_chany_top_out[15] ,
    \sb_8__1__0_chany_top_out[16] ,
    \sb_8__1__0_chany_top_out[17] ,
    \sb_8__1__0_chany_top_out[18] ,
    \sb_8__1__0_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__1_chany_bottom_out[0] ,
    \cby_8__1__1_chany_bottom_out[1] ,
    \cby_8__1__1_chany_bottom_out[2] ,
    \cby_8__1__1_chany_bottom_out[3] ,
    \cby_8__1__1_chany_bottom_out[4] ,
    \cby_8__1__1_chany_bottom_out[5] ,
    \cby_8__1__1_chany_bottom_out[6] ,
    \cby_8__1__1_chany_bottom_out[7] ,
    \cby_8__1__1_chany_bottom_out[8] ,
    \cby_8__1__1_chany_bottom_out[9] ,
    \cby_8__1__1_chany_bottom_out[10] ,
    \cby_8__1__1_chany_bottom_out[11] ,
    \cby_8__1__1_chany_bottom_out[12] ,
    \cby_8__1__1_chany_bottom_out[13] ,
    \cby_8__1__1_chany_bottom_out[14] ,
    \cby_8__1__1_chany_bottom_out[15] ,
    \cby_8__1__1_chany_bottom_out[16] ,
    \cby_8__1__1_chany_bottom_out[17] ,
    \cby_8__1__1_chany_bottom_out[18] ,
    \cby_8__1__1_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__1__1_chany_bottom_out[0] ,
    \sb_8__1__1_chany_bottom_out[1] ,
    \sb_8__1__1_chany_bottom_out[2] ,
    \sb_8__1__1_chany_bottom_out[3] ,
    \sb_8__1__1_chany_bottom_out[4] ,
    \sb_8__1__1_chany_bottom_out[5] ,
    \sb_8__1__1_chany_bottom_out[6] ,
    \sb_8__1__1_chany_bottom_out[7] ,
    \sb_8__1__1_chany_bottom_out[8] ,
    \sb_8__1__1_chany_bottom_out[9] ,
    \sb_8__1__1_chany_bottom_out[10] ,
    \sb_8__1__1_chany_bottom_out[11] ,
    \sb_8__1__1_chany_bottom_out[12] ,
    \sb_8__1__1_chany_bottom_out[13] ,
    \sb_8__1__1_chany_bottom_out[14] ,
    \sb_8__1__1_chany_bottom_out[15] ,
    \sb_8__1__1_chany_bottom_out[16] ,
    \sb_8__1__1_chany_bottom_out[17] ,
    \sb_8__1__1_chany_bottom_out[18] ,
    \sb_8__1__1_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__1_chany_top_out[0] ,
    \cby_8__1__1_chany_top_out[1] ,
    \cby_8__1__1_chany_top_out[2] ,
    \cby_8__1__1_chany_top_out[3] ,
    \cby_8__1__1_chany_top_out[4] ,
    \cby_8__1__1_chany_top_out[5] ,
    \cby_8__1__1_chany_top_out[6] ,
    \cby_8__1__1_chany_top_out[7] ,
    \cby_8__1__1_chany_top_out[8] ,
    \cby_8__1__1_chany_top_out[9] ,
    \cby_8__1__1_chany_top_out[10] ,
    \cby_8__1__1_chany_top_out[11] ,
    \cby_8__1__1_chany_top_out[12] ,
    \cby_8__1__1_chany_top_out[13] ,
    \cby_8__1__1_chany_top_out[14] ,
    \cby_8__1__1_chany_top_out[15] ,
    \cby_8__1__1_chany_top_out[16] ,
    \cby_8__1__1_chany_top_out[17] ,
    \cby_8__1__1_chany_top_out[18] ,
    \cby_8__1__1_chany_top_out[19] }));
 cby_2__1_ cby_8__3_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_58_ccff_tail),
    .ccff_tail(grid_io_right_5_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]),
    .left_grid_pin_16_(cby_8__1__2_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__2_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__2_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__2_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__2_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__2_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__2_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__2_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__2_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__2_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__2_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__2_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__2_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__2_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__2_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__2_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__2_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_5_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_5_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_S_out(\prog_clk_0_wires[207] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[206] ),
    .right_grid_pin_0_(cby_8__1__2_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__1__1_chany_top_out[0] ,
    \sb_8__1__1_chany_top_out[1] ,
    \sb_8__1__1_chany_top_out[2] ,
    \sb_8__1__1_chany_top_out[3] ,
    \sb_8__1__1_chany_top_out[4] ,
    \sb_8__1__1_chany_top_out[5] ,
    \sb_8__1__1_chany_top_out[6] ,
    \sb_8__1__1_chany_top_out[7] ,
    \sb_8__1__1_chany_top_out[8] ,
    \sb_8__1__1_chany_top_out[9] ,
    \sb_8__1__1_chany_top_out[10] ,
    \sb_8__1__1_chany_top_out[11] ,
    \sb_8__1__1_chany_top_out[12] ,
    \sb_8__1__1_chany_top_out[13] ,
    \sb_8__1__1_chany_top_out[14] ,
    \sb_8__1__1_chany_top_out[15] ,
    \sb_8__1__1_chany_top_out[16] ,
    \sb_8__1__1_chany_top_out[17] ,
    \sb_8__1__1_chany_top_out[18] ,
    \sb_8__1__1_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__2_chany_bottom_out[0] ,
    \cby_8__1__2_chany_bottom_out[1] ,
    \cby_8__1__2_chany_bottom_out[2] ,
    \cby_8__1__2_chany_bottom_out[3] ,
    \cby_8__1__2_chany_bottom_out[4] ,
    \cby_8__1__2_chany_bottom_out[5] ,
    \cby_8__1__2_chany_bottom_out[6] ,
    \cby_8__1__2_chany_bottom_out[7] ,
    \cby_8__1__2_chany_bottom_out[8] ,
    \cby_8__1__2_chany_bottom_out[9] ,
    \cby_8__1__2_chany_bottom_out[10] ,
    \cby_8__1__2_chany_bottom_out[11] ,
    \cby_8__1__2_chany_bottom_out[12] ,
    \cby_8__1__2_chany_bottom_out[13] ,
    \cby_8__1__2_chany_bottom_out[14] ,
    \cby_8__1__2_chany_bottom_out[15] ,
    \cby_8__1__2_chany_bottom_out[16] ,
    \cby_8__1__2_chany_bottom_out[17] ,
    \cby_8__1__2_chany_bottom_out[18] ,
    \cby_8__1__2_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__1__2_chany_bottom_out[0] ,
    \sb_8__1__2_chany_bottom_out[1] ,
    \sb_8__1__2_chany_bottom_out[2] ,
    \sb_8__1__2_chany_bottom_out[3] ,
    \sb_8__1__2_chany_bottom_out[4] ,
    \sb_8__1__2_chany_bottom_out[5] ,
    \sb_8__1__2_chany_bottom_out[6] ,
    \sb_8__1__2_chany_bottom_out[7] ,
    \sb_8__1__2_chany_bottom_out[8] ,
    \sb_8__1__2_chany_bottom_out[9] ,
    \sb_8__1__2_chany_bottom_out[10] ,
    \sb_8__1__2_chany_bottom_out[11] ,
    \sb_8__1__2_chany_bottom_out[12] ,
    \sb_8__1__2_chany_bottom_out[13] ,
    \sb_8__1__2_chany_bottom_out[14] ,
    \sb_8__1__2_chany_bottom_out[15] ,
    \sb_8__1__2_chany_bottom_out[16] ,
    \sb_8__1__2_chany_bottom_out[17] ,
    \sb_8__1__2_chany_bottom_out[18] ,
    \sb_8__1__2_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__2_chany_top_out[0] ,
    \cby_8__1__2_chany_top_out[1] ,
    \cby_8__1__2_chany_top_out[2] ,
    \cby_8__1__2_chany_top_out[3] ,
    \cby_8__1__2_chany_top_out[4] ,
    \cby_8__1__2_chany_top_out[5] ,
    \cby_8__1__2_chany_top_out[6] ,
    \cby_8__1__2_chany_top_out[7] ,
    \cby_8__1__2_chany_top_out[8] ,
    \cby_8__1__2_chany_top_out[9] ,
    \cby_8__1__2_chany_top_out[10] ,
    \cby_8__1__2_chany_top_out[11] ,
    \cby_8__1__2_chany_top_out[12] ,
    \cby_8__1__2_chany_top_out[13] ,
    \cby_8__1__2_chany_top_out[14] ,
    \cby_8__1__2_chany_top_out[15] ,
    \cby_8__1__2_chany_top_out[16] ,
    \cby_8__1__2_chany_top_out[17] ,
    \cby_8__1__2_chany_top_out[18] ,
    \cby_8__1__2_chany_top_out[19] }));
 cby_2__1_ cby_8__4_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_59_ccff_tail),
    .ccff_tail(grid_io_right_4_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]),
    .left_grid_pin_16_(cby_8__1__3_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__3_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__3_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__3_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__3_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__3_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__3_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__3_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__3_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__3_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__3_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__3_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__3_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__3_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__3_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__3_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__3_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_4_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_4_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_S_out(\prog_clk_0_wires[210] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[209] ),
    .right_grid_pin_0_(cby_8__1__3_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__1__2_chany_top_out[0] ,
    \sb_8__1__2_chany_top_out[1] ,
    \sb_8__1__2_chany_top_out[2] ,
    \sb_8__1__2_chany_top_out[3] ,
    \sb_8__1__2_chany_top_out[4] ,
    \sb_8__1__2_chany_top_out[5] ,
    \sb_8__1__2_chany_top_out[6] ,
    \sb_8__1__2_chany_top_out[7] ,
    \sb_8__1__2_chany_top_out[8] ,
    \sb_8__1__2_chany_top_out[9] ,
    \sb_8__1__2_chany_top_out[10] ,
    \sb_8__1__2_chany_top_out[11] ,
    \sb_8__1__2_chany_top_out[12] ,
    \sb_8__1__2_chany_top_out[13] ,
    \sb_8__1__2_chany_top_out[14] ,
    \sb_8__1__2_chany_top_out[15] ,
    \sb_8__1__2_chany_top_out[16] ,
    \sb_8__1__2_chany_top_out[17] ,
    \sb_8__1__2_chany_top_out[18] ,
    \sb_8__1__2_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__3_chany_bottom_out[0] ,
    \cby_8__1__3_chany_bottom_out[1] ,
    \cby_8__1__3_chany_bottom_out[2] ,
    \cby_8__1__3_chany_bottom_out[3] ,
    \cby_8__1__3_chany_bottom_out[4] ,
    \cby_8__1__3_chany_bottom_out[5] ,
    \cby_8__1__3_chany_bottom_out[6] ,
    \cby_8__1__3_chany_bottom_out[7] ,
    \cby_8__1__3_chany_bottom_out[8] ,
    \cby_8__1__3_chany_bottom_out[9] ,
    \cby_8__1__3_chany_bottom_out[10] ,
    \cby_8__1__3_chany_bottom_out[11] ,
    \cby_8__1__3_chany_bottom_out[12] ,
    \cby_8__1__3_chany_bottom_out[13] ,
    \cby_8__1__3_chany_bottom_out[14] ,
    \cby_8__1__3_chany_bottom_out[15] ,
    \cby_8__1__3_chany_bottom_out[16] ,
    \cby_8__1__3_chany_bottom_out[17] ,
    \cby_8__1__3_chany_bottom_out[18] ,
    \cby_8__1__3_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__1__3_chany_bottom_out[0] ,
    \sb_8__1__3_chany_bottom_out[1] ,
    \sb_8__1__3_chany_bottom_out[2] ,
    \sb_8__1__3_chany_bottom_out[3] ,
    \sb_8__1__3_chany_bottom_out[4] ,
    \sb_8__1__3_chany_bottom_out[5] ,
    \sb_8__1__3_chany_bottom_out[6] ,
    \sb_8__1__3_chany_bottom_out[7] ,
    \sb_8__1__3_chany_bottom_out[8] ,
    \sb_8__1__3_chany_bottom_out[9] ,
    \sb_8__1__3_chany_bottom_out[10] ,
    \sb_8__1__3_chany_bottom_out[11] ,
    \sb_8__1__3_chany_bottom_out[12] ,
    \sb_8__1__3_chany_bottom_out[13] ,
    \sb_8__1__3_chany_bottom_out[14] ,
    \sb_8__1__3_chany_bottom_out[15] ,
    \sb_8__1__3_chany_bottom_out[16] ,
    \sb_8__1__3_chany_bottom_out[17] ,
    \sb_8__1__3_chany_bottom_out[18] ,
    \sb_8__1__3_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__3_chany_top_out[0] ,
    \cby_8__1__3_chany_top_out[1] ,
    \cby_8__1__3_chany_top_out[2] ,
    \cby_8__1__3_chany_top_out[3] ,
    \cby_8__1__3_chany_top_out[4] ,
    \cby_8__1__3_chany_top_out[5] ,
    \cby_8__1__3_chany_top_out[6] ,
    \cby_8__1__3_chany_top_out[7] ,
    \cby_8__1__3_chany_top_out[8] ,
    \cby_8__1__3_chany_top_out[9] ,
    \cby_8__1__3_chany_top_out[10] ,
    \cby_8__1__3_chany_top_out[11] ,
    \cby_8__1__3_chany_top_out[12] ,
    \cby_8__1__3_chany_top_out[13] ,
    \cby_8__1__3_chany_top_out[14] ,
    \cby_8__1__3_chany_top_out[15] ,
    \cby_8__1__3_chany_top_out[16] ,
    \cby_8__1__3_chany_top_out[17] ,
    \cby_8__1__3_chany_top_out[18] ,
    \cby_8__1__3_chany_top_out[19] }));
 cby_2__1_ cby_8__5_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_60_ccff_tail),
    .ccff_tail(grid_io_right_3_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]),
    .left_grid_pin_16_(cby_8__1__4_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__4_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__4_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__4_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__4_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__4_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__4_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__4_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__4_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__4_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__4_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__4_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__4_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__4_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__4_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__4_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__4_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_3_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_3_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_S_out(\prog_clk_0_wires[213] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[212] ),
    .right_grid_pin_0_(cby_8__1__4_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__1__3_chany_top_out[0] ,
    \sb_8__1__3_chany_top_out[1] ,
    \sb_8__1__3_chany_top_out[2] ,
    \sb_8__1__3_chany_top_out[3] ,
    \sb_8__1__3_chany_top_out[4] ,
    \sb_8__1__3_chany_top_out[5] ,
    \sb_8__1__3_chany_top_out[6] ,
    \sb_8__1__3_chany_top_out[7] ,
    \sb_8__1__3_chany_top_out[8] ,
    \sb_8__1__3_chany_top_out[9] ,
    \sb_8__1__3_chany_top_out[10] ,
    \sb_8__1__3_chany_top_out[11] ,
    \sb_8__1__3_chany_top_out[12] ,
    \sb_8__1__3_chany_top_out[13] ,
    \sb_8__1__3_chany_top_out[14] ,
    \sb_8__1__3_chany_top_out[15] ,
    \sb_8__1__3_chany_top_out[16] ,
    \sb_8__1__3_chany_top_out[17] ,
    \sb_8__1__3_chany_top_out[18] ,
    \sb_8__1__3_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__4_chany_bottom_out[0] ,
    \cby_8__1__4_chany_bottom_out[1] ,
    \cby_8__1__4_chany_bottom_out[2] ,
    \cby_8__1__4_chany_bottom_out[3] ,
    \cby_8__1__4_chany_bottom_out[4] ,
    \cby_8__1__4_chany_bottom_out[5] ,
    \cby_8__1__4_chany_bottom_out[6] ,
    \cby_8__1__4_chany_bottom_out[7] ,
    \cby_8__1__4_chany_bottom_out[8] ,
    \cby_8__1__4_chany_bottom_out[9] ,
    \cby_8__1__4_chany_bottom_out[10] ,
    \cby_8__1__4_chany_bottom_out[11] ,
    \cby_8__1__4_chany_bottom_out[12] ,
    \cby_8__1__4_chany_bottom_out[13] ,
    \cby_8__1__4_chany_bottom_out[14] ,
    \cby_8__1__4_chany_bottom_out[15] ,
    \cby_8__1__4_chany_bottom_out[16] ,
    \cby_8__1__4_chany_bottom_out[17] ,
    \cby_8__1__4_chany_bottom_out[18] ,
    \cby_8__1__4_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__1__4_chany_bottom_out[0] ,
    \sb_8__1__4_chany_bottom_out[1] ,
    \sb_8__1__4_chany_bottom_out[2] ,
    \sb_8__1__4_chany_bottom_out[3] ,
    \sb_8__1__4_chany_bottom_out[4] ,
    \sb_8__1__4_chany_bottom_out[5] ,
    \sb_8__1__4_chany_bottom_out[6] ,
    \sb_8__1__4_chany_bottom_out[7] ,
    \sb_8__1__4_chany_bottom_out[8] ,
    \sb_8__1__4_chany_bottom_out[9] ,
    \sb_8__1__4_chany_bottom_out[10] ,
    \sb_8__1__4_chany_bottom_out[11] ,
    \sb_8__1__4_chany_bottom_out[12] ,
    \sb_8__1__4_chany_bottom_out[13] ,
    \sb_8__1__4_chany_bottom_out[14] ,
    \sb_8__1__4_chany_bottom_out[15] ,
    \sb_8__1__4_chany_bottom_out[16] ,
    \sb_8__1__4_chany_bottom_out[17] ,
    \sb_8__1__4_chany_bottom_out[18] ,
    \sb_8__1__4_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__4_chany_top_out[0] ,
    \cby_8__1__4_chany_top_out[1] ,
    \cby_8__1__4_chany_top_out[2] ,
    \cby_8__1__4_chany_top_out[3] ,
    \cby_8__1__4_chany_top_out[4] ,
    \cby_8__1__4_chany_top_out[5] ,
    \cby_8__1__4_chany_top_out[6] ,
    \cby_8__1__4_chany_top_out[7] ,
    \cby_8__1__4_chany_top_out[8] ,
    \cby_8__1__4_chany_top_out[9] ,
    \cby_8__1__4_chany_top_out[10] ,
    \cby_8__1__4_chany_top_out[11] ,
    \cby_8__1__4_chany_top_out[12] ,
    \cby_8__1__4_chany_top_out[13] ,
    \cby_8__1__4_chany_top_out[14] ,
    \cby_8__1__4_chany_top_out[15] ,
    \cby_8__1__4_chany_top_out[16] ,
    \cby_8__1__4_chany_top_out[17] ,
    \cby_8__1__4_chany_top_out[18] ,
    \cby_8__1__4_chany_top_out[19] }));
 cby_2__1_ cby_8__6_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_61_ccff_tail),
    .ccff_tail(grid_io_right_2_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]),
    .left_grid_pin_16_(cby_8__1__5_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__5_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__5_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__5_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__5_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__5_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__5_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__5_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__5_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__5_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__5_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__5_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__5_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__5_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__5_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__5_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__5_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_2_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_2_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_S_out(\prog_clk_0_wires[216] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[215] ),
    .right_grid_pin_0_(cby_8__1__5_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__1__4_chany_top_out[0] ,
    \sb_8__1__4_chany_top_out[1] ,
    \sb_8__1__4_chany_top_out[2] ,
    \sb_8__1__4_chany_top_out[3] ,
    \sb_8__1__4_chany_top_out[4] ,
    \sb_8__1__4_chany_top_out[5] ,
    \sb_8__1__4_chany_top_out[6] ,
    \sb_8__1__4_chany_top_out[7] ,
    \sb_8__1__4_chany_top_out[8] ,
    \sb_8__1__4_chany_top_out[9] ,
    \sb_8__1__4_chany_top_out[10] ,
    \sb_8__1__4_chany_top_out[11] ,
    \sb_8__1__4_chany_top_out[12] ,
    \sb_8__1__4_chany_top_out[13] ,
    \sb_8__1__4_chany_top_out[14] ,
    \sb_8__1__4_chany_top_out[15] ,
    \sb_8__1__4_chany_top_out[16] ,
    \sb_8__1__4_chany_top_out[17] ,
    \sb_8__1__4_chany_top_out[18] ,
    \sb_8__1__4_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__5_chany_bottom_out[0] ,
    \cby_8__1__5_chany_bottom_out[1] ,
    \cby_8__1__5_chany_bottom_out[2] ,
    \cby_8__1__5_chany_bottom_out[3] ,
    \cby_8__1__5_chany_bottom_out[4] ,
    \cby_8__1__5_chany_bottom_out[5] ,
    \cby_8__1__5_chany_bottom_out[6] ,
    \cby_8__1__5_chany_bottom_out[7] ,
    \cby_8__1__5_chany_bottom_out[8] ,
    \cby_8__1__5_chany_bottom_out[9] ,
    \cby_8__1__5_chany_bottom_out[10] ,
    \cby_8__1__5_chany_bottom_out[11] ,
    \cby_8__1__5_chany_bottom_out[12] ,
    \cby_8__1__5_chany_bottom_out[13] ,
    \cby_8__1__5_chany_bottom_out[14] ,
    \cby_8__1__5_chany_bottom_out[15] ,
    \cby_8__1__5_chany_bottom_out[16] ,
    \cby_8__1__5_chany_bottom_out[17] ,
    \cby_8__1__5_chany_bottom_out[18] ,
    \cby_8__1__5_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__1__5_chany_bottom_out[0] ,
    \sb_8__1__5_chany_bottom_out[1] ,
    \sb_8__1__5_chany_bottom_out[2] ,
    \sb_8__1__5_chany_bottom_out[3] ,
    \sb_8__1__5_chany_bottom_out[4] ,
    \sb_8__1__5_chany_bottom_out[5] ,
    \sb_8__1__5_chany_bottom_out[6] ,
    \sb_8__1__5_chany_bottom_out[7] ,
    \sb_8__1__5_chany_bottom_out[8] ,
    \sb_8__1__5_chany_bottom_out[9] ,
    \sb_8__1__5_chany_bottom_out[10] ,
    \sb_8__1__5_chany_bottom_out[11] ,
    \sb_8__1__5_chany_bottom_out[12] ,
    \sb_8__1__5_chany_bottom_out[13] ,
    \sb_8__1__5_chany_bottom_out[14] ,
    \sb_8__1__5_chany_bottom_out[15] ,
    \sb_8__1__5_chany_bottom_out[16] ,
    \sb_8__1__5_chany_bottom_out[17] ,
    \sb_8__1__5_chany_bottom_out[18] ,
    \sb_8__1__5_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__5_chany_top_out[0] ,
    \cby_8__1__5_chany_top_out[1] ,
    \cby_8__1__5_chany_top_out[2] ,
    \cby_8__1__5_chany_top_out[3] ,
    \cby_8__1__5_chany_top_out[4] ,
    \cby_8__1__5_chany_top_out[5] ,
    \cby_8__1__5_chany_top_out[6] ,
    \cby_8__1__5_chany_top_out[7] ,
    \cby_8__1__5_chany_top_out[8] ,
    \cby_8__1__5_chany_top_out[9] ,
    \cby_8__1__5_chany_top_out[10] ,
    \cby_8__1__5_chany_top_out[11] ,
    \cby_8__1__5_chany_top_out[12] ,
    \cby_8__1__5_chany_top_out[13] ,
    \cby_8__1__5_chany_top_out[14] ,
    \cby_8__1__5_chany_top_out[15] ,
    \cby_8__1__5_chany_top_out[16] ,
    \cby_8__1__5_chany_top_out[17] ,
    \cby_8__1__5_chany_top_out[18] ,
    \cby_8__1__5_chany_top_out[19] }));
 cby_2__1_ cby_8__7_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_62_ccff_tail),
    .ccff_tail(grid_io_right_1_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]),
    .left_grid_pin_16_(cby_8__1__6_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__6_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__6_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__6_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__6_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__6_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__6_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__6_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__6_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__6_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__6_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__6_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__6_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__6_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__6_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__6_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__6_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_1_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_1_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_S_out(\prog_clk_0_wires[219] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[218] ),
    .right_grid_pin_0_(cby_8__1__6_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__1__5_chany_top_out[0] ,
    \sb_8__1__5_chany_top_out[1] ,
    \sb_8__1__5_chany_top_out[2] ,
    \sb_8__1__5_chany_top_out[3] ,
    \sb_8__1__5_chany_top_out[4] ,
    \sb_8__1__5_chany_top_out[5] ,
    \sb_8__1__5_chany_top_out[6] ,
    \sb_8__1__5_chany_top_out[7] ,
    \sb_8__1__5_chany_top_out[8] ,
    \sb_8__1__5_chany_top_out[9] ,
    \sb_8__1__5_chany_top_out[10] ,
    \sb_8__1__5_chany_top_out[11] ,
    \sb_8__1__5_chany_top_out[12] ,
    \sb_8__1__5_chany_top_out[13] ,
    \sb_8__1__5_chany_top_out[14] ,
    \sb_8__1__5_chany_top_out[15] ,
    \sb_8__1__5_chany_top_out[16] ,
    \sb_8__1__5_chany_top_out[17] ,
    \sb_8__1__5_chany_top_out[18] ,
    \sb_8__1__5_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__6_chany_bottom_out[0] ,
    \cby_8__1__6_chany_bottom_out[1] ,
    \cby_8__1__6_chany_bottom_out[2] ,
    \cby_8__1__6_chany_bottom_out[3] ,
    \cby_8__1__6_chany_bottom_out[4] ,
    \cby_8__1__6_chany_bottom_out[5] ,
    \cby_8__1__6_chany_bottom_out[6] ,
    \cby_8__1__6_chany_bottom_out[7] ,
    \cby_8__1__6_chany_bottom_out[8] ,
    \cby_8__1__6_chany_bottom_out[9] ,
    \cby_8__1__6_chany_bottom_out[10] ,
    \cby_8__1__6_chany_bottom_out[11] ,
    \cby_8__1__6_chany_bottom_out[12] ,
    \cby_8__1__6_chany_bottom_out[13] ,
    \cby_8__1__6_chany_bottom_out[14] ,
    \cby_8__1__6_chany_bottom_out[15] ,
    \cby_8__1__6_chany_bottom_out[16] ,
    \cby_8__1__6_chany_bottom_out[17] ,
    \cby_8__1__6_chany_bottom_out[18] ,
    \cby_8__1__6_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__1__6_chany_bottom_out[0] ,
    \sb_8__1__6_chany_bottom_out[1] ,
    \sb_8__1__6_chany_bottom_out[2] ,
    \sb_8__1__6_chany_bottom_out[3] ,
    \sb_8__1__6_chany_bottom_out[4] ,
    \sb_8__1__6_chany_bottom_out[5] ,
    \sb_8__1__6_chany_bottom_out[6] ,
    \sb_8__1__6_chany_bottom_out[7] ,
    \sb_8__1__6_chany_bottom_out[8] ,
    \sb_8__1__6_chany_bottom_out[9] ,
    \sb_8__1__6_chany_bottom_out[10] ,
    \sb_8__1__6_chany_bottom_out[11] ,
    \sb_8__1__6_chany_bottom_out[12] ,
    \sb_8__1__6_chany_bottom_out[13] ,
    \sb_8__1__6_chany_bottom_out[14] ,
    \sb_8__1__6_chany_bottom_out[15] ,
    \sb_8__1__6_chany_bottom_out[16] ,
    \sb_8__1__6_chany_bottom_out[17] ,
    \sb_8__1__6_chany_bottom_out[18] ,
    \sb_8__1__6_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__6_chany_top_out[0] ,
    \cby_8__1__6_chany_top_out[1] ,
    \cby_8__1__6_chany_top_out[2] ,
    \cby_8__1__6_chany_top_out[3] ,
    \cby_8__1__6_chany_top_out[4] ,
    \cby_8__1__6_chany_top_out[5] ,
    \cby_8__1__6_chany_top_out[6] ,
    \cby_8__1__6_chany_top_out[7] ,
    \cby_8__1__6_chany_top_out[8] ,
    \cby_8__1__6_chany_top_out[9] ,
    \cby_8__1__6_chany_top_out[10] ,
    \cby_8__1__6_chany_top_out[11] ,
    \cby_8__1__6_chany_top_out[12] ,
    \cby_8__1__6_chany_top_out[13] ,
    \cby_8__1__6_chany_top_out[14] ,
    \cby_8__1__6_chany_top_out[15] ,
    \cby_8__1__6_chany_top_out[16] ,
    \cby_8__1__6_chany_top_out[17] ,
    \cby_8__1__6_chany_top_out[18] ,
    \cby_8__1__6_chany_top_out[19] }));
 cby_2__1_ cby_8__8_ (.IO_ISOL_N(IO_ISOL_N),
    .ccff_head(grid_clb_63_ccff_tail),
    .ccff_tail(grid_io_right_0_ccff_tail),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]),
    .left_grid_pin_16_(cby_8__1__7_left_grid_pin_16_),
    .left_grid_pin_17_(cby_8__1__7_left_grid_pin_17_),
    .left_grid_pin_18_(cby_8__1__7_left_grid_pin_18_),
    .left_grid_pin_19_(cby_8__1__7_left_grid_pin_19_),
    .left_grid_pin_20_(cby_8__1__7_left_grid_pin_20_),
    .left_grid_pin_21_(cby_8__1__7_left_grid_pin_21_),
    .left_grid_pin_22_(cby_8__1__7_left_grid_pin_22_),
    .left_grid_pin_23_(cby_8__1__7_left_grid_pin_23_),
    .left_grid_pin_24_(cby_8__1__7_left_grid_pin_24_),
    .left_grid_pin_25_(cby_8__1__7_left_grid_pin_25_),
    .left_grid_pin_26_(cby_8__1__7_left_grid_pin_26_),
    .left_grid_pin_27_(cby_8__1__7_left_grid_pin_27_),
    .left_grid_pin_28_(cby_8__1__7_left_grid_pin_28_),
    .left_grid_pin_29_(cby_8__1__7_left_grid_pin_29_),
    .left_grid_pin_30_(cby_8__1__7_left_grid_pin_30_),
    .left_grid_pin_31_(cby_8__1__7_left_grid_pin_31_),
    .left_width_0_height_0__pin_0_(cby_8__1__7_right_grid_pin_0_),
    .left_width_0_height_0__pin_1_lower(grid_io_right_0_left_width_0_height_0__pin_1_lower),
    .left_width_0_height_0__pin_1_upper(grid_io_right_0_left_width_0_height_0__pin_1_upper),
    .prog_clk_0_N_out(\prog_clk_0_wires[224] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[222] ),
    .prog_clk_0_W_in(\prog_clk_0_wires[221] ),
    .right_grid_pin_0_(cby_8__1__7_right_grid_pin_0_),
    .VPWR(VPWR),
    .VGND(VGND),
    .chany_bottom_in({\sb_8__1__6_chany_top_out[0] ,
    \sb_8__1__6_chany_top_out[1] ,
    \sb_8__1__6_chany_top_out[2] ,
    \sb_8__1__6_chany_top_out[3] ,
    \sb_8__1__6_chany_top_out[4] ,
    \sb_8__1__6_chany_top_out[5] ,
    \sb_8__1__6_chany_top_out[6] ,
    \sb_8__1__6_chany_top_out[7] ,
    \sb_8__1__6_chany_top_out[8] ,
    \sb_8__1__6_chany_top_out[9] ,
    \sb_8__1__6_chany_top_out[10] ,
    \sb_8__1__6_chany_top_out[11] ,
    \sb_8__1__6_chany_top_out[12] ,
    \sb_8__1__6_chany_top_out[13] ,
    \sb_8__1__6_chany_top_out[14] ,
    \sb_8__1__6_chany_top_out[15] ,
    \sb_8__1__6_chany_top_out[16] ,
    \sb_8__1__6_chany_top_out[17] ,
    \sb_8__1__6_chany_top_out[18] ,
    \sb_8__1__6_chany_top_out[19] }),
    .chany_bottom_out({\cby_8__1__7_chany_bottom_out[0] ,
    \cby_8__1__7_chany_bottom_out[1] ,
    \cby_8__1__7_chany_bottom_out[2] ,
    \cby_8__1__7_chany_bottom_out[3] ,
    \cby_8__1__7_chany_bottom_out[4] ,
    \cby_8__1__7_chany_bottom_out[5] ,
    \cby_8__1__7_chany_bottom_out[6] ,
    \cby_8__1__7_chany_bottom_out[7] ,
    \cby_8__1__7_chany_bottom_out[8] ,
    \cby_8__1__7_chany_bottom_out[9] ,
    \cby_8__1__7_chany_bottom_out[10] ,
    \cby_8__1__7_chany_bottom_out[11] ,
    \cby_8__1__7_chany_bottom_out[12] ,
    \cby_8__1__7_chany_bottom_out[13] ,
    \cby_8__1__7_chany_bottom_out[14] ,
    \cby_8__1__7_chany_bottom_out[15] ,
    \cby_8__1__7_chany_bottom_out[16] ,
    \cby_8__1__7_chany_bottom_out[17] ,
    \cby_8__1__7_chany_bottom_out[18] ,
    \cby_8__1__7_chany_bottom_out[19] }),
    .chany_top_in({\sb_8__8__0_chany_bottom_out[0] ,
    \sb_8__8__0_chany_bottom_out[1] ,
    \sb_8__8__0_chany_bottom_out[2] ,
    \sb_8__8__0_chany_bottom_out[3] ,
    \sb_8__8__0_chany_bottom_out[4] ,
    \sb_8__8__0_chany_bottom_out[5] ,
    \sb_8__8__0_chany_bottom_out[6] ,
    \sb_8__8__0_chany_bottom_out[7] ,
    \sb_8__8__0_chany_bottom_out[8] ,
    \sb_8__8__0_chany_bottom_out[9] ,
    \sb_8__8__0_chany_bottom_out[10] ,
    \sb_8__8__0_chany_bottom_out[11] ,
    \sb_8__8__0_chany_bottom_out[12] ,
    \sb_8__8__0_chany_bottom_out[13] ,
    \sb_8__8__0_chany_bottom_out[14] ,
    \sb_8__8__0_chany_bottom_out[15] ,
    \sb_8__8__0_chany_bottom_out[16] ,
    \sb_8__8__0_chany_bottom_out[17] ,
    \sb_8__8__0_chany_bottom_out[18] ,
    \sb_8__8__0_chany_bottom_out[19] }),
    .chany_top_out({\cby_8__1__7_chany_top_out[0] ,
    \cby_8__1__7_chany_top_out[1] ,
    \cby_8__1__7_chany_top_out[2] ,
    \cby_8__1__7_chany_top_out[3] ,
    \cby_8__1__7_chany_top_out[4] ,
    \cby_8__1__7_chany_top_out[5] ,
    \cby_8__1__7_chany_top_out[6] ,
    \cby_8__1__7_chany_top_out[7] ,
    \cby_8__1__7_chany_top_out[8] ,
    \cby_8__1__7_chany_top_out[9] ,
    \cby_8__1__7_chany_top_out[10] ,
    \cby_8__1__7_chany_top_out[11] ,
    \cby_8__1__7_chany_top_out[12] ,
    \cby_8__1__7_chany_top_out[13] ,
    \cby_8__1__7_chany_top_out[14] ,
    \cby_8__1__7_chany_top_out[15] ,
    \cby_8__1__7_chany_top_out[16] ,
    \cby_8__1__7_chany_top_out[17] ,
    \cby_8__1__7_chany_top_out[18] ,
    \cby_8__1__7_chany_top_out[19] }));
 grid_clb grid_clb_1__1_ (.SC_IN_TOP(\scff_Wires[15] ),
    .SC_OUT_BOT(\scff_Wires[17] ),
    .Test_en_E_in(\Test_enWires[16] ),
    .Test_en_W_in(\Test_enWires[16] ),
    .ccff_head(grid_io_left_0_ccff_tail),
    .ccff_tail(grid_clb_0_ccff_tail),
    .clk_0_N_in(\clk_1_wires[4] ),
    .clk_0_S_in(\clk_1_wires[4] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[1] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[4] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[4] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[0] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[3] ),
    .right_width_0_height_0__pin_16_(cby_1__1__0_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__0_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__0_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__0_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__0_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__0_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__0_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__0_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__0_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__0_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__0_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__0_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__0_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__0_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__0_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__0_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_0_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_0_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_0_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_0_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_0_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_0_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_0_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_0_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_0_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_0_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_0_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_0_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_0_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_0_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_0_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_0_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__0_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__0_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__0_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__0_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__0_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__0_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__0_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__0_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__0_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[0] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_0_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_0_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_0_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_0_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_0_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_0_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_0_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_0_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_0_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_0_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_0_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_0_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__0_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_0_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_0_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_0_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_0_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__0_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__0_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__0_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__0_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__0_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__0_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_1__2_ (.SC_IN_TOP(\scff_Wires[13] ),
    .SC_OUT_BOT(\scff_Wires[14] ),
    .Test_en_E_in(\Test_enWires[30] ),
    .Test_en_W_in(\Test_enWires[30] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[0] ),
    .ccff_head(grid_io_left_1_ccff_tail),
    .ccff_tail(grid_clb_1_ccff_tail),
    .clk_0_N_in(\clk_1_wires[3] ),
    .clk_0_S_in(\clk_1_wires[3] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[7] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[3] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[3] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[6] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[9] ),
    .right_width_0_height_0__pin_16_(cby_1__1__1_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__1_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__1_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__1_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__1_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__1_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__1_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__1_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__1_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__1_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__1_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__1_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__1_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__1_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__1_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__1_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_1_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_1_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_1_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_1_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_1_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_1_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_1_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_1_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_1_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_1_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_1_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_1_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_1_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_1_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_1_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_1_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__1_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__1_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__1_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__1_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__1_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__1_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__1_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__1_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__1_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[1] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_1_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_1_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_1_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_1_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_1_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_1_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_1_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_1_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_1_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_1_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_1_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_1_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__1_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_1_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_1_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_1_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_1_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__1_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__1_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__1_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__1_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__1_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__1_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_1__3_ (.SC_IN_TOP(\scff_Wires[11] ),
    .SC_OUT_BOT(\scff_Wires[12] ),
    .Test_en_E_in(\Test_enWires[44] ),
    .Test_en_W_in(\Test_enWires[44] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[1] ),
    .ccff_head(grid_io_left_2_ccff_tail),
    .ccff_tail(grid_clb_2_ccff_tail),
    .clk_0_N_in(\clk_1_wires[11] ),
    .clk_0_S_in(\clk_1_wires[11] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[12] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[11] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[11] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[11] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[14] ),
    .right_width_0_height_0__pin_16_(cby_1__1__2_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__2_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__2_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__2_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__2_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__2_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__2_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__2_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__2_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__2_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__2_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__2_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__2_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__2_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__2_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__2_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_2_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_2_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_2_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_2_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_2_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_2_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_2_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_2_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_2_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_2_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_2_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_2_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_2_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_2_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_2_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_2_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__2_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__2_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__2_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__2_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__2_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__2_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__2_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__2_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__2_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[2] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_2_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_2_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_2_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_2_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_2_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_2_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_2_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_2_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_2_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_2_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_2_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_2_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__2_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_2_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_2_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_2_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_2_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__2_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__2_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__2_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__2_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__2_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__2_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_1__4_ (.SC_IN_TOP(\scff_Wires[9] ),
    .SC_OUT_BOT(\scff_Wires[10] ),
    .Test_en_E_in(\Test_enWires[58] ),
    .Test_en_W_in(\Test_enWires[58] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[2] ),
    .ccff_head(grid_io_left_3_ccff_tail),
    .ccff_tail(grid_clb_3_ccff_tail),
    .clk_0_N_in(\clk_1_wires[10] ),
    .clk_0_S_in(\clk_1_wires[10] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[17] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[10] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[10] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[16] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[19] ),
    .right_width_0_height_0__pin_16_(cby_1__1__3_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__3_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__3_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__3_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__3_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__3_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__3_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__3_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__3_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__3_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__3_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__3_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__3_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__3_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__3_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__3_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_3_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_3_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_3_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_3_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_3_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_3_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_3_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_3_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_3_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_3_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_3_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_3_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_3_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_3_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_3_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_3_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__3_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__3_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__3_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__3_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__3_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__3_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__3_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__3_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__3_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[3] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_3_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_3_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_3_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_3_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_3_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_3_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_3_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_3_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_3_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_3_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_3_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_3_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__3_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_3_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_3_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_3_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_3_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__3_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__3_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__3_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__3_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__3_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__3_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_1__5_ (.SC_IN_TOP(\scff_Wires[7] ),
    .SC_OUT_BOT(\scff_Wires[8] ),
    .Test_en_E_in(\Test_enWires[72] ),
    .Test_en_W_in(\Test_enWires[72] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[3] ),
    .ccff_head(grid_io_left_4_ccff_tail),
    .ccff_tail(grid_clb_4_ccff_tail),
    .clk_0_N_in(\clk_1_wires[18] ),
    .clk_0_S_in(\clk_1_wires[18] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[22] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[18] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[18] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[21] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[24] ),
    .right_width_0_height_0__pin_16_(cby_1__1__4_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__4_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__4_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__4_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__4_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__4_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__4_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__4_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__4_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__4_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__4_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__4_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__4_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__4_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__4_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__4_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_4_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_4_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_4_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_4_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_4_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_4_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_4_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_4_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_4_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_4_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_4_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_4_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_4_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_4_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_4_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_4_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__4_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__4_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__4_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__4_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__4_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__4_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__4_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__4_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__4_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[4] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_4_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_4_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_4_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_4_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_4_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_4_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_4_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_4_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_4_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_4_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_4_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_4_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__4_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_4_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_4_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_4_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_4_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__4_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__4_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__4_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__4_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__4_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__4_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_1__6_ (.SC_IN_TOP(\scff_Wires[5] ),
    .SC_OUT_BOT(\scff_Wires[6] ),
    .Test_en_E_in(\Test_enWires[86] ),
    .Test_en_W_in(\Test_enWires[86] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[4] ),
    .ccff_head(grid_io_left_5_ccff_tail),
    .ccff_tail(grid_clb_5_ccff_tail),
    .clk_0_N_in(\clk_1_wires[17] ),
    .clk_0_S_in(\clk_1_wires[17] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[27] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[17] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[17] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[26] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[29] ),
    .right_width_0_height_0__pin_16_(cby_1__1__5_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__5_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__5_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__5_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__5_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__5_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__5_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__5_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__5_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__5_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__5_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__5_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__5_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__5_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__5_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__5_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_5_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_5_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_5_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_5_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_5_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_5_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_5_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_5_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_5_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_5_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_5_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_5_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_5_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_5_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_5_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_5_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__5_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__5_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__5_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__5_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__5_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__5_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__5_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__5_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__5_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[5] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_5_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_5_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_5_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_5_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_5_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_5_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_5_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_5_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_5_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_5_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_5_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_5_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__5_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_5_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_5_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_5_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_5_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__5_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__5_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__5_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__5_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__5_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__5_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_1__7_ (.SC_IN_TOP(\scff_Wires[3] ),
    .SC_OUT_BOT(\scff_Wires[4] ),
    .Test_en_E_in(\Test_enWires[100] ),
    .Test_en_W_in(\Test_enWires[100] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[5] ),
    .ccff_head(grid_io_left_6_ccff_tail),
    .ccff_tail(grid_clb_6_ccff_tail),
    .clk_0_N_in(\clk_1_wires[25] ),
    .clk_0_S_in(\clk_1_wires[25] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[32] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[25] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[25] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[31] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[34] ),
    .right_width_0_height_0__pin_16_(cby_1__1__6_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__6_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__6_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__6_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__6_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__6_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__6_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__6_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__6_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__6_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__6_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__6_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__6_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__6_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__6_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__6_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_6_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_6_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_6_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_6_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_6_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_6_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_6_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_6_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_6_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_6_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_6_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_6_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_6_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_6_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_6_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_6_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__6_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__6_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__6_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__6_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__6_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__6_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__6_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__6_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__6_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[6] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_6_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_6_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_6_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_6_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_6_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_6_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_6_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_6_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_6_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_6_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_6_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_6_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__6_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_6_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_6_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_6_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_6_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__6_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__6_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__6_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__6_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__6_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__6_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_1__8_ (.SC_IN_TOP(\scff_Wires[1] ),
    .SC_OUT_BOT(\scff_Wires[2] ),
    .Test_en_E_in(\Test_enWires[114] ),
    .Test_en_W_in(\Test_enWires[114] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[6] ),
    .ccff_head(grid_io_left_7_ccff_tail),
    .ccff_tail(grid_clb_7_ccff_tail),
    .clk_0_N_in(\clk_1_wires[24] ),
    .clk_0_S_in(\clk_1_wires[24] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[37] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[24] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[39] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[24] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[36] ),
    .prog_clk_0_W_out(\prog_clk_0_wires[41] ),
    .right_width_0_height_0__pin_16_(cby_1__1__7_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__7_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__7_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__7_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__7_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__7_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__7_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__7_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__7_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__7_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__7_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__7_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__7_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__7_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__7_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__7_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_7_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_7_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_7_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_7_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_7_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_7_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_7_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_7_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_7_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_7_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_7_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_7_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_7_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_7_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_7_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_7_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__0_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__0_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__0_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__0_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__0_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__0_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__0_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__0_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__0_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[0] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_7_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_7_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_7_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_7_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_7_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_7_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_7_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_7_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_7_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_7_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_7_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_7_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__0_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_7_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_7_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_7_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_7_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__0_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__0_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__0_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__0_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__0_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__0_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__1_ (.SC_IN_TOP(\scff_Wires[20] ),
    .SC_OUT_TOP(\scff_Wires[21] ),
    .Test_en_E_in(\Test_enWires[17] ),
    .Test_en_W_in(\Test_enWires[17] ),
    .Test_en_W_out(\Test_enWires[18] ),
    .ccff_head(cby_1__1__0_ccff_tail),
    .ccff_tail(grid_clb_8_ccff_tail),
    .clk_0_N_in(\clk_1_wires[6] ),
    .clk_0_S_in(\clk_1_wires[6] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[44] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[6] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[6] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[43] ),
    .right_width_0_height_0__pin_16_(cby_1__1__8_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__8_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__8_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__8_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__8_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__8_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__8_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__8_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__8_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__8_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__8_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__8_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__8_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__8_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__8_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__8_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_8_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_8_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_8_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_8_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_8_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_8_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_8_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_8_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_8_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_8_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_8_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_8_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_8_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_8_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_8_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_8_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__7_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__7_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__7_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__7_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__7_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__7_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__7_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__7_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__7_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[7] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_8_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_8_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_8_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_8_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_8_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_8_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_8_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_8_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_8_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_8_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_8_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_8_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__7_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_8_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_8_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_8_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_8_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__7_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__7_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__7_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__7_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__7_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__7_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__2_ (.SC_IN_TOP(\scff_Wires[22] ),
    .SC_OUT_TOP(\scff_Wires[23] ),
    .Test_en_E_in(\Test_enWires[31] ),
    .Test_en_W_in(\Test_enWires[31] ),
    .Test_en_W_out(\Test_enWires[32] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[7] ),
    .ccff_head(cby_1__1__1_ccff_tail),
    .ccff_tail(grid_clb_9_ccff_tail),
    .clk_0_N_in(\clk_1_wires[5] ),
    .clk_0_S_in(\clk_1_wires[5] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[47] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[5] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[5] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[46] ),
    .right_width_0_height_0__pin_16_(cby_1__1__9_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__9_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__9_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__9_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__9_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__9_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__9_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__9_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__9_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__9_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__9_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__9_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__9_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__9_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__9_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__9_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_9_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_9_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_9_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_9_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_9_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_9_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_9_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_9_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_9_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_9_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_9_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_9_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_9_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_9_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_9_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_9_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__8_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__8_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__8_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__8_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__8_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__8_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__8_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__8_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__8_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[8] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_9_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_9_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_9_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_9_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_9_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_9_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_9_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_9_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_9_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_9_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_9_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_9_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__8_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_9_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_9_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_9_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_9_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__8_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__8_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__8_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__8_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__8_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__8_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__3_ (.SC_IN_TOP(\scff_Wires[24] ),
    .SC_OUT_TOP(\scff_Wires[25] ),
    .Test_en_E_in(\Test_enWires[45] ),
    .Test_en_W_in(\Test_enWires[45] ),
    .Test_en_W_out(\Test_enWires[46] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[8] ),
    .ccff_head(cby_1__1__2_ccff_tail),
    .ccff_tail(grid_clb_10_ccff_tail),
    .clk_0_N_in(\clk_1_wires[13] ),
    .clk_0_S_in(\clk_1_wires[13] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[50] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[13] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[13] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[49] ),
    .right_width_0_height_0__pin_16_(cby_1__1__10_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__10_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__10_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__10_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__10_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__10_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__10_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__10_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__10_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__10_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__10_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__10_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__10_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__10_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__10_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__10_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_10_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_10_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_10_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_10_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_10_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_10_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_10_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_10_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_10_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_10_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_10_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_10_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_10_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_10_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_10_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_10_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__9_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__9_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__9_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__9_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__9_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__9_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__9_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__9_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__9_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[9] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_10_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_10_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_10_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_10_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_10_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_10_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_10_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_10_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_10_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_10_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_10_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_10_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__9_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_10_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_10_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_10_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_10_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__9_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__9_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__9_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__9_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__9_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__9_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__4_ (.SC_IN_TOP(\scff_Wires[26] ),
    .SC_OUT_TOP(\scff_Wires[27] ),
    .Test_en_E_in(\Test_enWires[59] ),
    .Test_en_W_in(\Test_enWires[59] ),
    .Test_en_W_out(\Test_enWires[60] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[9] ),
    .ccff_head(cby_1__1__3_ccff_tail),
    .ccff_tail(grid_clb_11_ccff_tail),
    .clk_0_N_in(\clk_1_wires[12] ),
    .clk_0_S_in(\clk_1_wires[12] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[53] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[12] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[12] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[52] ),
    .right_width_0_height_0__pin_16_(cby_1__1__11_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__11_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__11_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__11_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__11_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__11_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__11_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__11_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__11_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__11_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__11_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__11_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__11_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__11_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__11_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__11_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_11_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_11_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_11_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_11_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_11_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_11_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_11_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_11_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_11_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_11_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_11_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_11_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_11_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_11_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_11_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_11_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__10_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__10_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__10_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__10_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__10_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__10_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__10_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__10_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__10_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[10] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_11_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_11_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_11_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_11_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_11_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_11_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_11_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_11_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_11_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_11_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_11_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_11_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__10_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_11_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_11_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_11_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_11_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__10_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__10_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__10_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__10_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__10_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__10_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__5_ (.SC_IN_TOP(\scff_Wires[28] ),
    .SC_OUT_TOP(\scff_Wires[29] ),
    .Test_en_E_in(\Test_enWires[73] ),
    .Test_en_W_in(\Test_enWires[73] ),
    .Test_en_W_out(\Test_enWires[74] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[10] ),
    .ccff_head(cby_1__1__4_ccff_tail),
    .ccff_tail(grid_clb_12_ccff_tail),
    .clk_0_N_in(\clk_1_wires[20] ),
    .clk_0_S_in(\clk_1_wires[20] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[56] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[20] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[20] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[55] ),
    .right_width_0_height_0__pin_16_(cby_1__1__12_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__12_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__12_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__12_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__12_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__12_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__12_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__12_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__12_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__12_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__12_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__12_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__12_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__12_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__12_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__12_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_12_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_12_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_12_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_12_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_12_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_12_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_12_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_12_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_12_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_12_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_12_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_12_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_12_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_12_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_12_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_12_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__11_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__11_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__11_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__11_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__11_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__11_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__11_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__11_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__11_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[11] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_12_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_12_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_12_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_12_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_12_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_12_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_12_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_12_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_12_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_12_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_12_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_12_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__11_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_12_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_12_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_12_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_12_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__11_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__11_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__11_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__11_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__11_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__11_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__6_ (.SC_IN_TOP(\scff_Wires[30] ),
    .SC_OUT_TOP(\scff_Wires[31] ),
    .Test_en_E_in(\Test_enWires[87] ),
    .Test_en_W_in(\Test_enWires[87] ),
    .Test_en_W_out(\Test_enWires[88] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[11] ),
    .ccff_head(cby_1__1__5_ccff_tail),
    .ccff_tail(grid_clb_13_ccff_tail),
    .clk_0_N_in(\clk_1_wires[19] ),
    .clk_0_S_in(\clk_1_wires[19] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[59] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[19] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[19] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[58] ),
    .right_width_0_height_0__pin_16_(cby_1__1__13_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__13_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__13_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__13_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__13_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__13_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__13_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__13_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__13_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__13_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__13_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__13_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__13_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__13_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__13_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__13_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_13_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_13_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_13_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_13_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_13_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_13_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_13_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_13_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_13_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_13_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_13_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_13_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_13_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_13_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_13_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_13_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__12_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__12_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__12_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__12_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__12_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__12_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__12_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__12_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__12_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[12] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_13_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_13_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_13_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_13_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_13_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_13_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_13_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_13_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_13_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_13_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_13_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_13_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__12_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_13_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_13_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_13_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_13_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__12_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__12_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__12_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__12_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__12_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__12_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__7_ (.SC_IN_TOP(\scff_Wires[32] ),
    .SC_OUT_TOP(\scff_Wires[33] ),
    .Test_en_E_in(\Test_enWires[101] ),
    .Test_en_W_in(\Test_enWires[101] ),
    .Test_en_W_out(\Test_enWires[102] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[12] ),
    .ccff_head(cby_1__1__6_ccff_tail),
    .ccff_tail(grid_clb_14_ccff_tail),
    .clk_0_N_in(\clk_1_wires[27] ),
    .clk_0_S_in(\clk_1_wires[27] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[62] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[27] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[27] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[61] ),
    .right_width_0_height_0__pin_16_(cby_1__1__14_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__14_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__14_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__14_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__14_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__14_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__14_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__14_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__14_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__14_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__14_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__14_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__14_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__14_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__14_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__14_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_14_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_14_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_14_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_14_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_14_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_14_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_14_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_14_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_14_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_14_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_14_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_14_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_14_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_14_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_14_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_14_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__13_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__13_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__13_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__13_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__13_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__13_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__13_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__13_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__13_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[13] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_14_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_14_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_14_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_14_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_14_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_14_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_14_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_14_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_14_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_14_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_14_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_14_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__13_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_14_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_14_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_14_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_14_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__13_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__13_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__13_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__13_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__13_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__13_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_2__8_ (.SC_IN_TOP(\scff_Wires[34] ),
    .SC_OUT_TOP(\scff_Wires[35] ),
    .Test_en_E_in(\Test_enWires[115] ),
    .Test_en_W_in(\Test_enWires[115] ),
    .Test_en_W_out(\Test_enWires[116] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[13] ),
    .ccff_head(cby_1__1__7_ccff_tail),
    .ccff_tail(grid_clb_15_ccff_tail),
    .clk_0_N_in(\clk_1_wires[26] ),
    .clk_0_S_in(\clk_1_wires[26] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[65] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[26] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[67] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[26] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[64] ),
    .right_width_0_height_0__pin_16_(cby_1__1__15_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__15_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__15_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__15_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__15_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__15_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__15_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__15_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__15_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__15_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__15_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__15_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__15_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__15_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__15_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__15_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_15_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_15_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_15_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_15_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_15_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_15_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_15_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_15_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_15_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_15_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_15_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_15_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_15_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_15_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_15_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_15_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__1_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__1_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__1_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__1_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__1_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__1_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__1_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__1_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__1_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[1] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_15_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_15_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_15_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_15_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_15_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_15_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_15_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_15_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_15_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_15_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_15_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_15_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__1_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_15_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_15_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_15_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_15_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__1_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__1_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__1_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__1_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__1_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__1_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__1_ (.SC_IN_TOP(\scff_Wires[52] ),
    .SC_OUT_BOT(\scff_Wires[54] ),
    .Test_en_E_in(\Test_enWires[19] ),
    .Test_en_W_in(\Test_enWires[19] ),
    .Test_en_W_out(\Test_enWires[20] ),
    .ccff_head(cby_1__1__8_ccff_tail),
    .ccff_tail(grid_clb_16_ccff_tail),
    .clk_0_N_in(\clk_1_wires[32] ),
    .clk_0_S_in(\clk_1_wires[32] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[70] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[32] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[32] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[69] ),
    .right_width_0_height_0__pin_16_(cby_1__1__16_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__16_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__16_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__16_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__16_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__16_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__16_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__16_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__16_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__16_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__16_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__16_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__16_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__16_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__16_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__16_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_16_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_16_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_16_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_16_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_16_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_16_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_16_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_16_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_16_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_16_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_16_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_16_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_16_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_16_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_16_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_16_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__14_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__14_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__14_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__14_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__14_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__14_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__14_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__14_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__14_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[14] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_16_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_16_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_16_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_16_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_16_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_16_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_16_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_16_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_16_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_16_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_16_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_16_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__14_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_16_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_16_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_16_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_16_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__14_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__14_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__14_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__14_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__14_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__14_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__2_ (.SC_IN_TOP(\scff_Wires[50] ),
    .SC_OUT_BOT(\scff_Wires[51] ),
    .Test_en_E_in(\Test_enWires[33] ),
    .Test_en_W_in(\Test_enWires[33] ),
    .Test_en_W_out(\Test_enWires[34] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[14] ),
    .ccff_head(cby_1__1__9_ccff_tail),
    .ccff_tail(grid_clb_17_ccff_tail),
    .clk_0_N_in(\clk_1_wires[31] ),
    .clk_0_S_in(\clk_1_wires[31] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[73] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[31] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[31] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[72] ),
    .right_width_0_height_0__pin_16_(cby_1__1__17_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__17_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__17_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__17_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__17_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__17_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__17_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__17_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__17_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__17_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__17_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__17_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__17_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__17_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__17_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__17_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_17_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_17_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_17_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_17_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_17_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_17_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_17_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_17_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_17_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_17_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_17_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_17_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_17_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_17_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_17_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_17_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__15_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__15_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__15_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__15_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__15_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__15_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__15_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__15_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__15_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[15] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_17_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_17_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_17_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_17_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_17_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_17_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_17_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_17_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_17_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_17_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_17_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_17_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__15_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_17_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_17_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_17_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_17_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__15_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__15_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__15_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__15_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__15_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__15_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__3_ (.SC_IN_TOP(\scff_Wires[48] ),
    .SC_OUT_BOT(\scff_Wires[49] ),
    .Test_en_E_in(\Test_enWires[47] ),
    .Test_en_W_in(\Test_enWires[47] ),
    .Test_en_W_out(\Test_enWires[48] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[15] ),
    .ccff_head(cby_1__1__10_ccff_tail),
    .ccff_tail(grid_clb_18_ccff_tail),
    .clk_0_N_in(\clk_1_wires[39] ),
    .clk_0_S_in(\clk_1_wires[39] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[76] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[39] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[39] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[75] ),
    .right_width_0_height_0__pin_16_(cby_1__1__18_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__18_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__18_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__18_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__18_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__18_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__18_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__18_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__18_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__18_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__18_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__18_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__18_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__18_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__18_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__18_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_18_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_18_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_18_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_18_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_18_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_18_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_18_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_18_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_18_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_18_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_18_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_18_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_18_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_18_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_18_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_18_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__16_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__16_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__16_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__16_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__16_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__16_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__16_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__16_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__16_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[16] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_18_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_18_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_18_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_18_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_18_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_18_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_18_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_18_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_18_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_18_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_18_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_18_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__16_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_18_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_18_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_18_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_18_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__16_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__16_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__16_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__16_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__16_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__16_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__4_ (.SC_IN_TOP(\scff_Wires[46] ),
    .SC_OUT_BOT(\scff_Wires[47] ),
    .Test_en_E_in(\Test_enWires[61] ),
    .Test_en_W_in(\Test_enWires[61] ),
    .Test_en_W_out(\Test_enWires[62] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[16] ),
    .ccff_head(cby_1__1__11_ccff_tail),
    .ccff_tail(grid_clb_19_ccff_tail),
    .clk_0_N_in(\clk_1_wires[38] ),
    .clk_0_S_in(\clk_1_wires[38] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[79] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[38] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[38] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[78] ),
    .right_width_0_height_0__pin_16_(cby_1__1__19_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__19_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__19_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__19_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__19_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__19_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__19_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__19_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__19_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__19_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__19_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__19_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__19_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__19_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__19_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__19_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_19_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_19_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_19_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_19_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_19_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_19_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_19_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_19_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_19_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_19_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_19_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_19_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_19_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_19_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_19_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_19_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__17_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__17_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__17_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__17_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__17_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__17_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__17_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__17_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__17_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[17] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_19_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_19_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_19_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_19_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_19_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_19_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_19_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_19_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_19_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_19_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_19_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_19_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__17_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_19_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_19_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_19_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_19_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__17_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__17_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__17_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__17_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__17_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__17_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__5_ (.SC_IN_TOP(\scff_Wires[44] ),
    .SC_OUT_BOT(\scff_Wires[45] ),
    .Test_en_E_in(\Test_enWires[75] ),
    .Test_en_W_in(\Test_enWires[75] ),
    .Test_en_W_out(\Test_enWires[76] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[17] ),
    .ccff_head(cby_1__1__12_ccff_tail),
    .ccff_tail(grid_clb_20_ccff_tail),
    .clk_0_N_in(\clk_1_wires[46] ),
    .clk_0_S_in(\clk_1_wires[46] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[82] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[46] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[46] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[81] ),
    .right_width_0_height_0__pin_16_(cby_1__1__20_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__20_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__20_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__20_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__20_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__20_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__20_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__20_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__20_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__20_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__20_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__20_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__20_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__20_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__20_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__20_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_20_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_20_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_20_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_20_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_20_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_20_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_20_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_20_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_20_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_20_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_20_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_20_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_20_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_20_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_20_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_20_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__18_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__18_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__18_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__18_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__18_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__18_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__18_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__18_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__18_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[18] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_20_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_20_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_20_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_20_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_20_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_20_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_20_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_20_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_20_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_20_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_20_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_20_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__18_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_20_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_20_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_20_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_20_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__18_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__18_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__18_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__18_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__18_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__18_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__6_ (.SC_IN_TOP(\scff_Wires[42] ),
    .SC_OUT_BOT(\scff_Wires[43] ),
    .Test_en_E_in(\Test_enWires[89] ),
    .Test_en_W_in(\Test_enWires[89] ),
    .Test_en_W_out(\Test_enWires[90] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[18] ),
    .ccff_head(cby_1__1__13_ccff_tail),
    .ccff_tail(grid_clb_21_ccff_tail),
    .clk_0_N_in(\clk_1_wires[45] ),
    .clk_0_S_in(\clk_1_wires[45] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[85] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[45] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[45] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[84] ),
    .right_width_0_height_0__pin_16_(cby_1__1__21_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__21_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__21_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__21_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__21_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__21_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__21_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__21_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__21_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__21_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__21_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__21_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__21_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__21_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__21_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__21_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_21_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_21_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_21_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_21_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_21_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_21_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_21_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_21_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_21_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_21_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_21_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_21_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_21_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_21_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_21_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_21_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__19_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__19_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__19_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__19_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__19_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__19_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__19_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__19_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__19_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[19] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_21_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_21_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_21_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_21_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_21_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_21_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_21_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_21_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_21_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_21_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_21_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_21_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__19_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_21_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_21_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_21_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_21_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__19_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__19_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__19_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__19_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__19_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__19_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__7_ (.SC_IN_TOP(\scff_Wires[40] ),
    .SC_OUT_BOT(\scff_Wires[41] ),
    .Test_en_E_in(\Test_enWires[103] ),
    .Test_en_W_in(\Test_enWires[103] ),
    .Test_en_W_out(\Test_enWires[104] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[19] ),
    .ccff_head(cby_1__1__14_ccff_tail),
    .ccff_tail(grid_clb_22_ccff_tail),
    .clk_0_N_in(\clk_1_wires[53] ),
    .clk_0_S_in(\clk_1_wires[53] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[88] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[53] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[53] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[87] ),
    .right_width_0_height_0__pin_16_(cby_1__1__22_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__22_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__22_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__22_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__22_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__22_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__22_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__22_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__22_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__22_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__22_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__22_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__22_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__22_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__22_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__22_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_22_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_22_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_22_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_22_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_22_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_22_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_22_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_22_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_22_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_22_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_22_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_22_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_22_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_22_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_22_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_22_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__20_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__20_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__20_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__20_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__20_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__20_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__20_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__20_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__20_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[20] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_22_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_22_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_22_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_22_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_22_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_22_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_22_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_22_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_22_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_22_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_22_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_22_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__20_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_22_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_22_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_22_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_22_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__20_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__20_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__20_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__20_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__20_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__20_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_3__8_ (.SC_IN_TOP(\scff_Wires[38] ),
    .SC_OUT_BOT(\scff_Wires[39] ),
    .Test_en_E_in(\Test_enWires[117] ),
    .Test_en_W_in(\Test_enWires[117] ),
    .Test_en_W_out(\Test_enWires[118] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[20] ),
    .ccff_head(cby_1__1__15_ccff_tail),
    .ccff_tail(grid_clb_23_ccff_tail),
    .clk_0_N_in(\clk_1_wires[52] ),
    .clk_0_S_in(\clk_1_wires[52] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[91] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[52] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[93] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[52] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[90] ),
    .right_width_0_height_0__pin_16_(cby_1__1__23_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__23_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__23_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__23_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__23_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__23_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__23_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__23_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__23_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__23_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__23_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__23_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__23_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__23_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__23_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__23_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_23_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_23_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_23_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_23_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_23_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_23_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_23_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_23_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_23_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_23_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_23_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_23_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_23_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_23_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_23_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_23_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__2_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__2_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__2_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__2_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__2_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__2_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__2_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__2_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__2_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[2] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_23_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_23_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_23_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_23_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_23_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_23_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_23_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_23_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_23_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_23_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_23_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_23_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__2_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_23_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_23_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_23_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_23_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__2_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__2_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__2_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__2_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__2_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__2_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__1_ (.SC_IN_TOP(\scff_Wires[57] ),
    .SC_OUT_TOP(\scff_Wires[58] ),
    .Test_en_E_in(\Test_enWires[21] ),
    .Test_en_W_in(\Test_enWires[21] ),
    .Test_en_W_out(\Test_enWires[22] ),
    .ccff_head(cby_1__1__16_ccff_tail),
    .ccff_tail(grid_clb_24_ccff_tail),
    .clk_0_N_in(\clk_1_wires[34] ),
    .clk_0_S_in(\clk_1_wires[34] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[96] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[34] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[34] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[95] ),
    .right_width_0_height_0__pin_16_(cby_1__1__24_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__24_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__24_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__24_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__24_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__24_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__24_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__24_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__24_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__24_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__24_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__24_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__24_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__24_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__24_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__24_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_24_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_24_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_24_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_24_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_24_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_24_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_24_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_24_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_24_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_24_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_24_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_24_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_24_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_24_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_24_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_24_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__21_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__21_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__21_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__21_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__21_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__21_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__21_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__21_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__21_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[21] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_24_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_24_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_24_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_24_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_24_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_24_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_24_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_24_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_24_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_24_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_24_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_24_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__21_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_24_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_24_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_24_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_24_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__21_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__21_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__21_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__21_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__21_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__21_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__2_ (.SC_IN_TOP(\scff_Wires[59] ),
    .SC_OUT_TOP(\scff_Wires[60] ),
    .Test_en_E_in(\Test_enWires[35] ),
    .Test_en_W_in(\Test_enWires[35] ),
    .Test_en_W_out(\Test_enWires[36] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[21] ),
    .ccff_head(cby_1__1__17_ccff_tail),
    .ccff_tail(grid_clb_25_ccff_tail),
    .clk_0_N_in(\clk_1_wires[33] ),
    .clk_0_S_in(\clk_1_wires[33] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[99] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[33] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[33] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[98] ),
    .right_width_0_height_0__pin_16_(cby_1__1__25_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__25_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__25_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__25_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__25_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__25_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__25_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__25_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__25_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__25_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__25_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__25_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__25_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__25_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__25_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__25_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_25_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_25_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_25_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_25_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_25_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_25_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_25_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_25_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_25_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_25_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_25_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_25_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_25_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_25_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_25_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_25_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__22_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__22_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__22_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__22_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__22_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__22_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__22_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__22_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__22_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[22] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_25_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_25_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_25_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_25_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_25_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_25_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_25_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_25_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_25_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_25_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_25_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_25_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__22_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_25_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_25_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_25_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_25_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__22_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__22_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__22_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__22_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__22_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__22_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__3_ (.SC_IN_TOP(\scff_Wires[61] ),
    .SC_OUT_TOP(\scff_Wires[62] ),
    .Test_en_E_in(\Test_enWires[49] ),
    .Test_en_W_in(\Test_enWires[49] ),
    .Test_en_W_out(\Test_enWires[50] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[22] ),
    .ccff_head(cby_1__1__18_ccff_tail),
    .ccff_tail(grid_clb_26_ccff_tail),
    .clk_0_N_in(\clk_1_wires[41] ),
    .clk_0_S_in(\clk_1_wires[41] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[102] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[41] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[41] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[101] ),
    .right_width_0_height_0__pin_16_(cby_1__1__26_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__26_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__26_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__26_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__26_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__26_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__26_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__26_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__26_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__26_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__26_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__26_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__26_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__26_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__26_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__26_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_26_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_26_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_26_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_26_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_26_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_26_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_26_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_26_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_26_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_26_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_26_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_26_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_26_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_26_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_26_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_26_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__23_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__23_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__23_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__23_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__23_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__23_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__23_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__23_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__23_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[23] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_26_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_26_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_26_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_26_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_26_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_26_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_26_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_26_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_26_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_26_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_26_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_26_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__23_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_26_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_26_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_26_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_26_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__23_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__23_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__23_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__23_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__23_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__23_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__4_ (.SC_IN_TOP(\scff_Wires[63] ),
    .SC_OUT_TOP(\scff_Wires[64] ),
    .Test_en_E_in(\Test_enWires[63] ),
    .Test_en_W_in(\Test_enWires[63] ),
    .Test_en_W_out(\Test_enWires[64] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[23] ),
    .ccff_head(cby_1__1__19_ccff_tail),
    .ccff_tail(grid_clb_27_ccff_tail),
    .clk_0_N_in(\clk_1_wires[40] ),
    .clk_0_S_in(\clk_1_wires[40] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[105] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[40] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[40] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[104] ),
    .right_width_0_height_0__pin_16_(cby_1__1__27_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__27_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__27_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__27_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__27_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__27_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__27_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__27_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__27_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__27_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__27_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__27_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__27_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__27_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__27_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__27_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_27_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_27_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_27_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_27_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_27_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_27_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_27_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_27_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_27_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_27_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_27_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_27_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_27_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_27_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_27_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_27_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__24_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__24_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__24_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__24_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__24_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__24_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__24_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__24_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__24_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[24] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_27_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_27_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_27_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_27_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_27_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_27_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_27_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_27_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_27_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_27_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_27_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_27_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__24_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_27_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_27_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_27_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_27_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__24_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__24_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__24_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__24_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__24_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__24_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__5_ (.SC_IN_TOP(\scff_Wires[65] ),
    .SC_OUT_TOP(\scff_Wires[66] ),
    .Test_en_E_in(\Test_enWires[77] ),
    .Test_en_W_in(\Test_enWires[77] ),
    .Test_en_W_out(\Test_enWires[78] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[24] ),
    .ccff_head(cby_1__1__20_ccff_tail),
    .ccff_tail(grid_clb_28_ccff_tail),
    .clk_0_N_in(\clk_1_wires[48] ),
    .clk_0_S_in(\clk_1_wires[48] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[108] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[48] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[48] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[107] ),
    .right_width_0_height_0__pin_16_(cby_1__1__28_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__28_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__28_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__28_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__28_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__28_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__28_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__28_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__28_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__28_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__28_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__28_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__28_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__28_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__28_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__28_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_28_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_28_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_28_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_28_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_28_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_28_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_28_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_28_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_28_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_28_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_28_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_28_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_28_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_28_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_28_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_28_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__25_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__25_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__25_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__25_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__25_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__25_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__25_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__25_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__25_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[25] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_28_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_28_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_28_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_28_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_28_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_28_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_28_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_28_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_28_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_28_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_28_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_28_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__25_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_28_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_28_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_28_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_28_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__25_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__25_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__25_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__25_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__25_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__25_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__6_ (.SC_IN_TOP(\scff_Wires[67] ),
    .SC_OUT_TOP(\scff_Wires[68] ),
    .Test_en_E_in(\Test_enWires[91] ),
    .Test_en_W_in(\Test_enWires[91] ),
    .Test_en_W_out(\Test_enWires[92] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[25] ),
    .ccff_head(cby_1__1__21_ccff_tail),
    .ccff_tail(grid_clb_29_ccff_tail),
    .clk_0_N_in(\clk_1_wires[47] ),
    .clk_0_S_in(\clk_1_wires[47] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[111] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[47] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[47] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[110] ),
    .right_width_0_height_0__pin_16_(cby_1__1__29_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__29_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__29_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__29_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__29_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__29_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__29_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__29_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__29_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__29_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__29_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__29_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__29_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__29_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__29_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__29_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_29_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_29_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_29_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_29_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_29_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_29_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_29_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_29_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_29_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_29_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_29_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_29_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_29_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_29_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_29_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_29_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__26_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__26_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__26_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__26_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__26_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__26_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__26_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__26_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__26_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[26] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_29_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_29_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_29_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_29_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_29_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_29_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_29_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_29_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_29_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_29_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_29_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_29_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__26_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_29_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_29_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_29_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_29_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__26_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__26_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__26_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__26_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__26_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__26_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__7_ (.SC_IN_TOP(\scff_Wires[69] ),
    .SC_OUT_TOP(\scff_Wires[70] ),
    .Test_en_E_in(\Test_enWires[105] ),
    .Test_en_W_in(\Test_enWires[105] ),
    .Test_en_W_out(\Test_enWires[106] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[26] ),
    .ccff_head(cby_1__1__22_ccff_tail),
    .ccff_tail(grid_clb_30_ccff_tail),
    .clk_0_N_in(\clk_1_wires[55] ),
    .clk_0_S_in(\clk_1_wires[55] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[114] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[55] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[55] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[113] ),
    .right_width_0_height_0__pin_16_(cby_1__1__30_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__30_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__30_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__30_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__30_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__30_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__30_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__30_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__30_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__30_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__30_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__30_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__30_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__30_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__30_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__30_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_30_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_30_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_30_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_30_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_30_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_30_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_30_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_30_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_30_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_30_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_30_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_30_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_30_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_30_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_30_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_30_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__27_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__27_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__27_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__27_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__27_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__27_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__27_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__27_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__27_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[27] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_30_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_30_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_30_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_30_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_30_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_30_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_30_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_30_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_30_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_30_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_30_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_30_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__27_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_30_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_30_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_30_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_30_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__27_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__27_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__27_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__27_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__27_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__27_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_4__8_ (.SC_IN_TOP(\scff_Wires[71] ),
    .SC_OUT_TOP(\scff_Wires[72] ),
    .Test_en_E_in(\Test_enWires[119] ),
    .Test_en_W_in(\Test_enWires[119] ),
    .Test_en_W_out(\Test_enWires[120] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[27] ),
    .ccff_head(cby_1__1__23_ccff_tail),
    .ccff_tail(grid_clb_31_ccff_tail),
    .clk_0_N_in(\clk_1_wires[54] ),
    .clk_0_S_in(\clk_1_wires[54] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[117] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[54] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[119] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[54] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[116] ),
    .right_width_0_height_0__pin_16_(cby_1__1__31_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__31_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__31_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__31_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__31_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__31_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__31_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__31_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__31_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__31_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__31_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__31_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__31_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__31_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__31_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__31_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_31_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_31_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_31_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_31_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_31_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_31_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_31_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_31_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_31_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_31_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_31_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_31_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_31_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_31_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_31_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_31_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__3_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__3_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__3_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__3_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__3_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__3_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__3_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__3_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__3_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[3] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_31_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_31_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_31_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_31_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_31_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_31_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_31_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_31_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_31_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_31_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_31_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_31_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__3_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_31_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_31_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_31_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_31_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__3_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__3_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__3_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__3_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__3_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__3_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__1_ (.SC_IN_TOP(\scff_Wires[89] ),
    .SC_OUT_BOT(\scff_Wires[91] ),
    .Test_en_E_in(\Test_enWires[23] ),
    .Test_en_E_out(\Test_enWires[24] ),
    .Test_en_W_in(\Test_enWires[23] ),
    .ccff_head(cby_1__1__24_ccff_tail),
    .ccff_tail(grid_clb_32_ccff_tail),
    .clk_0_N_in(\clk_1_wires[60] ),
    .clk_0_S_in(\clk_1_wires[60] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[122] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[60] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[60] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[121] ),
    .right_width_0_height_0__pin_16_(cby_1__1__32_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__32_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__32_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__32_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__32_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__32_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__32_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__32_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__32_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__32_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__32_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__32_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__32_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__32_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__32_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__32_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_32_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_32_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_32_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_32_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_32_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_32_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_32_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_32_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_32_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_32_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_32_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_32_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_32_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_32_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_32_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_32_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__28_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__28_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__28_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__28_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__28_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__28_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__28_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__28_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__28_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[28] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_32_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_32_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_32_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_32_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_32_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_32_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_32_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_32_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_32_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_32_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_32_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_32_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__28_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_32_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_32_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_32_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_32_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__28_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__28_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__28_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__28_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__28_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__28_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__2_ (.SC_IN_TOP(\scff_Wires[87] ),
    .SC_OUT_BOT(\scff_Wires[88] ),
    .Test_en_E_in(\Test_enWires[37] ),
    .Test_en_E_out(\Test_enWires[38] ),
    .Test_en_W_in(\Test_enWires[37] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[28] ),
    .ccff_head(cby_1__1__25_ccff_tail),
    .ccff_tail(grid_clb_33_ccff_tail),
    .clk_0_N_in(\clk_1_wires[59] ),
    .clk_0_S_in(\clk_1_wires[59] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[125] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[59] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[59] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[124] ),
    .right_width_0_height_0__pin_16_(cby_1__1__33_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__33_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__33_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__33_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__33_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__33_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__33_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__33_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__33_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__33_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__33_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__33_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__33_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__33_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__33_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__33_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_33_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_33_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_33_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_33_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_33_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_33_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_33_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_33_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_33_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_33_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_33_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_33_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_33_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_33_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_33_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_33_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__29_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__29_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__29_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__29_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__29_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__29_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__29_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__29_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__29_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[29] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_33_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_33_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_33_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_33_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_33_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_33_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_33_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_33_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_33_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_33_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_33_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_33_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__29_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_33_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_33_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_33_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_33_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__29_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__29_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__29_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__29_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__29_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__29_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__3_ (.SC_IN_TOP(\scff_Wires[85] ),
    .SC_OUT_BOT(\scff_Wires[86] ),
    .Test_en_E_in(\Test_enWires[51] ),
    .Test_en_E_out(\Test_enWires[52] ),
    .Test_en_W_in(\Test_enWires[51] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[29] ),
    .ccff_head(cby_1__1__26_ccff_tail),
    .ccff_tail(grid_clb_34_ccff_tail),
    .clk_0_N_in(\clk_1_wires[67] ),
    .clk_0_S_in(\clk_1_wires[67] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[128] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[67] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[67] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[127] ),
    .right_width_0_height_0__pin_16_(cby_1__1__34_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__34_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__34_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__34_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__34_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__34_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__34_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__34_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__34_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__34_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__34_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__34_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__34_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__34_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__34_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__34_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_34_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_34_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_34_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_34_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_34_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_34_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_34_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_34_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_34_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_34_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_34_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_34_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_34_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_34_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_34_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_34_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__30_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__30_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__30_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__30_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__30_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__30_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__30_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__30_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__30_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[30] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_34_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_34_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_34_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_34_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_34_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_34_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_34_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_34_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_34_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_34_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_34_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_34_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__30_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_34_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_34_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_34_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_34_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__30_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__30_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__30_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__30_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__30_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__30_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__4_ (.SC_IN_TOP(\scff_Wires[83] ),
    .SC_OUT_BOT(\scff_Wires[84] ),
    .Test_en_E_in(\Test_enWires[65] ),
    .Test_en_E_out(\Test_enWires[66] ),
    .Test_en_W_in(\Test_enWires[65] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[30] ),
    .ccff_head(cby_1__1__27_ccff_tail),
    .ccff_tail(grid_clb_35_ccff_tail),
    .clk_0_N_in(\clk_1_wires[66] ),
    .clk_0_S_in(\clk_1_wires[66] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[131] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[66] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[66] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[130] ),
    .right_width_0_height_0__pin_16_(cby_1__1__35_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__35_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__35_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__35_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__35_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__35_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__35_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__35_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__35_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__35_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__35_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__35_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__35_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__35_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__35_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__35_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_35_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_35_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_35_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_35_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_35_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_35_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_35_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_35_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_35_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_35_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_35_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_35_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_35_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_35_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_35_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_35_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__31_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__31_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__31_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__31_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__31_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__31_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__31_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__31_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__31_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[31] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_35_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_35_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_35_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_35_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_35_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_35_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_35_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_35_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_35_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_35_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_35_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_35_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__31_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_35_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_35_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_35_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_35_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__31_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__31_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__31_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__31_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__31_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__31_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__5_ (.SC_IN_TOP(\scff_Wires[81] ),
    .SC_OUT_BOT(\scff_Wires[82] ),
    .Test_en_E_in(\Test_enWires[79] ),
    .Test_en_E_out(\Test_enWires[80] ),
    .Test_en_W_in(\Test_enWires[79] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[31] ),
    .ccff_head(cby_1__1__28_ccff_tail),
    .ccff_tail(grid_clb_36_ccff_tail),
    .clk_0_N_in(\clk_1_wires[74] ),
    .clk_0_S_in(\clk_1_wires[74] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[134] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[74] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[74] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[133] ),
    .right_width_0_height_0__pin_16_(cby_1__1__36_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__36_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__36_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__36_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__36_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__36_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__36_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__36_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__36_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__36_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__36_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__36_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__36_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__36_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__36_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__36_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_36_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_36_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_36_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_36_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_36_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_36_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_36_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_36_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_36_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_36_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_36_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_36_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_36_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_36_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_36_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_36_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__32_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__32_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__32_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__32_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__32_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__32_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__32_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__32_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__32_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[32] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_36_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_36_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_36_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_36_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_36_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_36_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_36_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_36_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_36_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_36_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_36_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_36_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__32_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_36_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_36_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_36_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_36_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__32_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__32_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__32_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__32_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__32_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__32_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__6_ (.SC_IN_TOP(\scff_Wires[79] ),
    .SC_OUT_BOT(\scff_Wires[80] ),
    .Test_en_E_in(\Test_enWires[93] ),
    .Test_en_E_out(\Test_enWires[94] ),
    .Test_en_W_in(\Test_enWires[93] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[32] ),
    .ccff_head(cby_1__1__29_ccff_tail),
    .ccff_tail(grid_clb_37_ccff_tail),
    .clk_0_N_in(\clk_1_wires[73] ),
    .clk_0_S_in(\clk_1_wires[73] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[137] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[73] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[73] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[136] ),
    .right_width_0_height_0__pin_16_(cby_1__1__37_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__37_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__37_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__37_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__37_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__37_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__37_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__37_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__37_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__37_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__37_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__37_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__37_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__37_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__37_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__37_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_37_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_37_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_37_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_37_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_37_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_37_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_37_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_37_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_37_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_37_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_37_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_37_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_37_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_37_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_37_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_37_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__33_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__33_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__33_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__33_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__33_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__33_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__33_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__33_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__33_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[33] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_37_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_37_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_37_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_37_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_37_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_37_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_37_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_37_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_37_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_37_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_37_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_37_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__33_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_37_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_37_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_37_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_37_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__33_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__33_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__33_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__33_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__33_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__33_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__7_ (.SC_IN_TOP(\scff_Wires[77] ),
    .SC_OUT_BOT(\scff_Wires[78] ),
    .Test_en_E_in(\Test_enWires[107] ),
    .Test_en_E_out(\Test_enWires[108] ),
    .Test_en_W_in(\Test_enWires[107] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[33] ),
    .ccff_head(cby_1__1__30_ccff_tail),
    .ccff_tail(grid_clb_38_ccff_tail),
    .clk_0_N_in(\clk_1_wires[81] ),
    .clk_0_S_in(\clk_1_wires[81] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[140] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[81] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[81] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[139] ),
    .right_width_0_height_0__pin_16_(cby_1__1__38_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__38_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__38_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__38_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__38_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__38_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__38_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__38_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__38_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__38_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__38_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__38_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__38_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__38_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__38_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__38_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_38_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_38_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_38_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_38_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_38_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_38_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_38_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_38_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_38_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_38_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_38_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_38_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_38_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_38_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_38_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_38_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__34_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__34_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__34_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__34_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__34_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__34_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__34_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__34_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__34_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[34] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_38_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_38_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_38_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_38_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_38_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_38_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_38_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_38_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_38_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_38_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_38_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_38_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__34_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_38_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_38_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_38_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_38_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__34_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__34_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__34_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__34_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__34_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__34_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_5__8_ (.SC_IN_TOP(\scff_Wires[75] ),
    .SC_OUT_BOT(\scff_Wires[76] ),
    .Test_en_E_in(\Test_enWires[121] ),
    .Test_en_E_out(\Test_enWires[122] ),
    .Test_en_W_in(\Test_enWires[121] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[34] ),
    .ccff_head(cby_1__1__31_ccff_tail),
    .ccff_tail(grid_clb_39_ccff_tail),
    .clk_0_N_in(\clk_1_wires[80] ),
    .clk_0_S_in(\clk_1_wires[80] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[143] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[80] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[145] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[80] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[142] ),
    .right_width_0_height_0__pin_16_(cby_1__1__39_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__39_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__39_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__39_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__39_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__39_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__39_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__39_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__39_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__39_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__39_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__39_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__39_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__39_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__39_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__39_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_39_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_39_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_39_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_39_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_39_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_39_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_39_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_39_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_39_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_39_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_39_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_39_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_39_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_39_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_39_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_39_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__4_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__4_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__4_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__4_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__4_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__4_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__4_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__4_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__4_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[4] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_39_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_39_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_39_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_39_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_39_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_39_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_39_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_39_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_39_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_39_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_39_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_39_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__4_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_39_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_39_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_39_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_39_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__4_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__4_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__4_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__4_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__4_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__4_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__1_ (.SC_IN_TOP(\scff_Wires[94] ),
    .SC_OUT_TOP(\scff_Wires[95] ),
    .Test_en_E_in(\Test_enWires[25] ),
    .Test_en_E_out(\Test_enWires[26] ),
    .Test_en_W_in(\Test_enWires[25] ),
    .ccff_head(cby_1__1__32_ccff_tail),
    .ccff_tail(grid_clb_40_ccff_tail),
    .clk_0_N_in(\clk_1_wires[62] ),
    .clk_0_S_in(\clk_1_wires[62] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[148] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[62] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[62] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[147] ),
    .right_width_0_height_0__pin_16_(cby_1__1__40_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__40_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__40_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__40_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__40_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__40_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__40_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__40_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__40_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__40_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__40_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__40_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__40_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__40_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__40_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__40_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_40_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_40_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_40_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_40_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_40_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_40_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_40_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_40_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_40_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_40_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_40_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_40_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_40_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_40_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_40_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_40_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__35_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__35_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__35_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__35_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__35_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__35_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__35_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__35_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__35_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[35] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_40_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_40_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_40_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_40_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_40_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_40_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_40_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_40_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_40_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_40_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_40_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_40_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__35_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_40_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_40_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_40_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_40_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__35_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__35_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__35_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__35_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__35_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__35_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__2_ (.SC_IN_TOP(\scff_Wires[96] ),
    .SC_OUT_TOP(\scff_Wires[97] ),
    .Test_en_E_in(\Test_enWires[39] ),
    .Test_en_E_out(\Test_enWires[40] ),
    .Test_en_W_in(\Test_enWires[39] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[35] ),
    .ccff_head(cby_1__1__33_ccff_tail),
    .ccff_tail(grid_clb_41_ccff_tail),
    .clk_0_N_in(\clk_1_wires[61] ),
    .clk_0_S_in(\clk_1_wires[61] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[151] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[61] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[61] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[150] ),
    .right_width_0_height_0__pin_16_(cby_1__1__41_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__41_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__41_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__41_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__41_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__41_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__41_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__41_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__41_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__41_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__41_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__41_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__41_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__41_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__41_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__41_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_41_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_41_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_41_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_41_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_41_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_41_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_41_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_41_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_41_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_41_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_41_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_41_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_41_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_41_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_41_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_41_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__36_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__36_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__36_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__36_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__36_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__36_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__36_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__36_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__36_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[36] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_41_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_41_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_41_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_41_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_41_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_41_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_41_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_41_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_41_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_41_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_41_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_41_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__36_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_41_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_41_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_41_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_41_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__36_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__36_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__36_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__36_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__36_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__36_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__3_ (.SC_IN_TOP(\scff_Wires[98] ),
    .SC_OUT_TOP(\scff_Wires[99] ),
    .Test_en_E_in(\Test_enWires[53] ),
    .Test_en_E_out(\Test_enWires[54] ),
    .Test_en_W_in(\Test_enWires[53] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[36] ),
    .ccff_head(cby_1__1__34_ccff_tail),
    .ccff_tail(grid_clb_42_ccff_tail),
    .clk_0_N_in(\clk_1_wires[69] ),
    .clk_0_S_in(\clk_1_wires[69] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[154] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[69] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[69] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[153] ),
    .right_width_0_height_0__pin_16_(cby_1__1__42_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__42_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__42_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__42_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__42_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__42_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__42_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__42_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__42_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__42_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__42_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__42_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__42_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__42_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__42_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__42_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_42_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_42_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_42_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_42_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_42_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_42_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_42_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_42_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_42_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_42_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_42_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_42_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_42_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_42_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_42_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_42_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__37_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__37_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__37_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__37_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__37_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__37_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__37_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__37_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__37_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[37] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_42_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_42_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_42_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_42_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_42_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_42_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_42_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_42_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_42_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_42_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_42_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_42_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__37_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_42_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_42_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_42_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_42_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__37_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__37_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__37_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__37_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__37_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__37_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__4_ (.SC_IN_TOP(\scff_Wires[100] ),
    .SC_OUT_TOP(\scff_Wires[101] ),
    .Test_en_E_in(\Test_enWires[67] ),
    .Test_en_E_out(\Test_enWires[68] ),
    .Test_en_W_in(\Test_enWires[67] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[37] ),
    .ccff_head(cby_1__1__35_ccff_tail),
    .ccff_tail(grid_clb_43_ccff_tail),
    .clk_0_N_in(\clk_1_wires[68] ),
    .clk_0_S_in(\clk_1_wires[68] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[157] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[68] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[68] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[156] ),
    .right_width_0_height_0__pin_16_(cby_1__1__43_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__43_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__43_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__43_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__43_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__43_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__43_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__43_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__43_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__43_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__43_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__43_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__43_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__43_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__43_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__43_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_43_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_43_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_43_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_43_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_43_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_43_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_43_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_43_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_43_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_43_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_43_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_43_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_43_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_43_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_43_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_43_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__38_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__38_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__38_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__38_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__38_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__38_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__38_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__38_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__38_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[38] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_43_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_43_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_43_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_43_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_43_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_43_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_43_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_43_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_43_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_43_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_43_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_43_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__38_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_43_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_43_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_43_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_43_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__38_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__38_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__38_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__38_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__38_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__38_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__5_ (.SC_IN_TOP(\scff_Wires[102] ),
    .SC_OUT_TOP(\scff_Wires[103] ),
    .Test_en_E_in(\Test_enWires[81] ),
    .Test_en_E_out(\Test_enWires[82] ),
    .Test_en_W_in(\Test_enWires[81] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[38] ),
    .ccff_head(cby_1__1__36_ccff_tail),
    .ccff_tail(grid_clb_44_ccff_tail),
    .clk_0_N_in(\clk_1_wires[76] ),
    .clk_0_S_in(\clk_1_wires[76] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[160] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[76] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[76] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[159] ),
    .right_width_0_height_0__pin_16_(cby_1__1__44_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__44_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__44_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__44_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__44_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__44_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__44_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__44_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__44_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__44_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__44_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__44_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__44_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__44_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__44_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__44_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_44_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_44_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_44_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_44_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_44_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_44_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_44_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_44_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_44_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_44_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_44_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_44_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_44_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_44_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_44_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_44_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__39_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__39_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__39_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__39_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__39_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__39_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__39_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__39_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__39_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[39] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_44_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_44_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_44_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_44_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_44_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_44_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_44_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_44_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_44_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_44_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_44_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_44_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__39_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_44_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_44_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_44_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_44_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__39_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__39_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__39_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__39_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__39_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__39_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__6_ (.SC_IN_TOP(\scff_Wires[104] ),
    .SC_OUT_TOP(\scff_Wires[105] ),
    .Test_en_E_in(\Test_enWires[95] ),
    .Test_en_E_out(\Test_enWires[96] ),
    .Test_en_W_in(\Test_enWires[95] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[39] ),
    .ccff_head(cby_1__1__37_ccff_tail),
    .ccff_tail(grid_clb_45_ccff_tail),
    .clk_0_N_in(\clk_1_wires[75] ),
    .clk_0_S_in(\clk_1_wires[75] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[163] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[75] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[75] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[162] ),
    .right_width_0_height_0__pin_16_(cby_1__1__45_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__45_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__45_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__45_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__45_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__45_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__45_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__45_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__45_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__45_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__45_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__45_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__45_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__45_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__45_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__45_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_45_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_45_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_45_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_45_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_45_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_45_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_45_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_45_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_45_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_45_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_45_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_45_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_45_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_45_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_45_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_45_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__40_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__40_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__40_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__40_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__40_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__40_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__40_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__40_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__40_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[40] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_45_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_45_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_45_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_45_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_45_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_45_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_45_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_45_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_45_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_45_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_45_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_45_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__40_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_45_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_45_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_45_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_45_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__40_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__40_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__40_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__40_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__40_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__40_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__7_ (.SC_IN_TOP(\scff_Wires[106] ),
    .SC_OUT_TOP(\scff_Wires[107] ),
    .Test_en_E_in(\Test_enWires[109] ),
    .Test_en_E_out(\Test_enWires[110] ),
    .Test_en_W_in(\Test_enWires[109] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[40] ),
    .ccff_head(cby_1__1__38_ccff_tail),
    .ccff_tail(grid_clb_46_ccff_tail),
    .clk_0_N_in(\clk_1_wires[83] ),
    .clk_0_S_in(\clk_1_wires[83] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[166] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[83] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[83] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[165] ),
    .right_width_0_height_0__pin_16_(cby_1__1__46_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__46_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__46_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__46_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__46_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__46_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__46_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__46_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__46_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__46_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__46_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__46_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__46_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__46_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__46_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__46_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_46_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_46_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_46_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_46_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_46_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_46_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_46_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_46_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_46_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_46_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_46_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_46_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_46_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_46_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_46_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_46_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__41_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__41_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__41_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__41_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__41_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__41_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__41_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__41_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__41_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[41] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_46_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_46_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_46_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_46_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_46_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_46_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_46_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_46_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_46_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_46_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_46_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_46_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__41_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_46_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_46_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_46_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_46_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__41_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__41_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__41_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__41_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__41_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__41_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_6__8_ (.SC_IN_TOP(\scff_Wires[108] ),
    .SC_OUT_TOP(\scff_Wires[109] ),
    .Test_en_E_in(\Test_enWires[123] ),
    .Test_en_E_out(\Test_enWires[124] ),
    .Test_en_W_in(\Test_enWires[123] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[41] ),
    .ccff_head(cby_1__1__39_ccff_tail),
    .ccff_tail(grid_clb_47_ccff_tail),
    .clk_0_N_in(\clk_1_wires[82] ),
    .clk_0_S_in(\clk_1_wires[82] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[169] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[82] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[171] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[82] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[168] ),
    .right_width_0_height_0__pin_16_(cby_1__1__47_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__47_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__47_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__47_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__47_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__47_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__47_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__47_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__47_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__47_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__47_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__47_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__47_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__47_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__47_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__47_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_47_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_47_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_47_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_47_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_47_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_47_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_47_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_47_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_47_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_47_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_47_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_47_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_47_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_47_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_47_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_47_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__5_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__5_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__5_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__5_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__5_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__5_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__5_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__5_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__5_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[5] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_47_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_47_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_47_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_47_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_47_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_47_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_47_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_47_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_47_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_47_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_47_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_47_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__5_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_47_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_47_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_47_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_47_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__5_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__5_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__5_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__5_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__5_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__5_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__1_ (.SC_IN_TOP(\scff_Wires[126] ),
    .SC_OUT_BOT(\scff_Wires[128] ),
    .Test_en_E_in(\Test_enWires[27] ),
    .Test_en_E_out(\Test_enWires[28] ),
    .Test_en_W_in(\Test_enWires[27] ),
    .ccff_head(cby_1__1__40_ccff_tail),
    .ccff_tail(grid_clb_48_ccff_tail),
    .clk_0_N_in(\clk_1_wires[88] ),
    .clk_0_S_in(\clk_1_wires[88] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[174] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[88] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[88] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[173] ),
    .right_width_0_height_0__pin_16_(cby_1__1__48_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__48_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__48_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__48_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__48_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__48_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__48_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__48_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__48_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__48_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__48_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__48_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__48_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__48_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__48_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__48_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_48_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_48_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_48_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_48_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_48_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_48_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_48_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_48_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_48_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_48_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_48_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_48_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_48_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_48_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_48_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_48_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__42_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__42_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__42_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__42_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__42_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__42_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__42_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__42_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__42_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[42] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_48_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_48_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_48_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_48_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_48_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_48_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_48_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_48_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_48_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_48_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_48_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_48_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__42_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_48_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_48_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_48_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_48_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__42_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__42_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__42_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__42_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__42_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__42_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__2_ (.SC_IN_TOP(\scff_Wires[124] ),
    .SC_OUT_BOT(\scff_Wires[125] ),
    .Test_en_E_in(\Test_enWires[41] ),
    .Test_en_E_out(\Test_enWires[42] ),
    .Test_en_W_in(\Test_enWires[41] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[42] ),
    .ccff_head(cby_1__1__41_ccff_tail),
    .ccff_tail(grid_clb_49_ccff_tail),
    .clk_0_N_in(\clk_1_wires[87] ),
    .clk_0_S_in(\clk_1_wires[87] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[177] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[87] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[87] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[176] ),
    .right_width_0_height_0__pin_16_(cby_1__1__49_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__49_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__49_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__49_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__49_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__49_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__49_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__49_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__49_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__49_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__49_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__49_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__49_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__49_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__49_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__49_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_49_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_49_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_49_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_49_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_49_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_49_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_49_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_49_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_49_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_49_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_49_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_49_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_49_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_49_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_49_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_49_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__43_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__43_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__43_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__43_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__43_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__43_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__43_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__43_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__43_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[43] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_49_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_49_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_49_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_49_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_49_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_49_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_49_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_49_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_49_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_49_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_49_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_49_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__43_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_49_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_49_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_49_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_49_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__43_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__43_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__43_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__43_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__43_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__43_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__3_ (.SC_IN_TOP(\scff_Wires[122] ),
    .SC_OUT_BOT(\scff_Wires[123] ),
    .Test_en_E_in(\Test_enWires[55] ),
    .Test_en_E_out(\Test_enWires[56] ),
    .Test_en_W_in(\Test_enWires[55] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[43] ),
    .ccff_head(cby_1__1__42_ccff_tail),
    .ccff_tail(grid_clb_50_ccff_tail),
    .clk_0_N_in(\clk_1_wires[95] ),
    .clk_0_S_in(\clk_1_wires[95] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[180] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[95] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[95] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[179] ),
    .right_width_0_height_0__pin_16_(cby_1__1__50_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__50_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__50_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__50_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__50_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__50_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__50_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__50_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__50_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__50_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__50_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__50_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__50_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__50_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__50_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__50_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_50_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_50_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_50_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_50_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_50_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_50_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_50_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_50_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_50_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_50_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_50_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_50_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_50_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_50_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_50_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_50_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__44_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__44_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__44_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__44_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__44_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__44_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__44_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__44_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__44_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[44] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_50_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_50_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_50_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_50_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_50_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_50_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_50_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_50_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_50_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_50_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_50_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_50_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__44_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_50_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_50_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_50_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_50_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__44_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__44_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__44_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__44_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__44_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__44_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__4_ (.SC_IN_TOP(\scff_Wires[120] ),
    .SC_OUT_BOT(\scff_Wires[121] ),
    .Test_en_E_in(\Test_enWires[69] ),
    .Test_en_E_out(\Test_enWires[70] ),
    .Test_en_W_in(\Test_enWires[69] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[44] ),
    .ccff_head(cby_1__1__43_ccff_tail),
    .ccff_tail(grid_clb_51_ccff_tail),
    .clk_0_N_in(\clk_1_wires[94] ),
    .clk_0_S_in(\clk_1_wires[94] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[183] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[94] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[94] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[182] ),
    .right_width_0_height_0__pin_16_(cby_1__1__51_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__51_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__51_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__51_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__51_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__51_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__51_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__51_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__51_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__51_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__51_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__51_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__51_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__51_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__51_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__51_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_51_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_51_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_51_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_51_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_51_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_51_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_51_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_51_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_51_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_51_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_51_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_51_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_51_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_51_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_51_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_51_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__45_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__45_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__45_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__45_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__45_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__45_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__45_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__45_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__45_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[45] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_51_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_51_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_51_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_51_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_51_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_51_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_51_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_51_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_51_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_51_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_51_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_51_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__45_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_51_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_51_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_51_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_51_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__45_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__45_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__45_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__45_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__45_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__45_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__5_ (.SC_IN_TOP(\scff_Wires[118] ),
    .SC_OUT_BOT(\scff_Wires[119] ),
    .Test_en_E_in(\Test_enWires[83] ),
    .Test_en_E_out(\Test_enWires[84] ),
    .Test_en_W_in(\Test_enWires[83] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[45] ),
    .ccff_head(cby_1__1__44_ccff_tail),
    .ccff_tail(grid_clb_52_ccff_tail),
    .clk_0_N_in(\clk_1_wires[102] ),
    .clk_0_S_in(\clk_1_wires[102] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[186] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[102] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[102] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[185] ),
    .right_width_0_height_0__pin_16_(cby_1__1__52_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__52_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__52_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__52_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__52_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__52_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__52_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__52_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__52_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__52_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__52_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__52_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__52_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__52_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__52_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__52_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_52_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_52_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_52_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_52_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_52_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_52_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_52_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_52_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_52_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_52_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_52_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_52_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_52_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_52_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_52_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_52_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__46_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__46_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__46_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__46_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__46_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__46_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__46_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__46_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__46_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[46] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_52_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_52_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_52_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_52_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_52_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_52_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_52_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_52_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_52_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_52_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_52_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_52_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__46_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_52_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_52_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_52_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_52_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__46_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__46_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__46_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__46_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__46_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__46_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__6_ (.SC_IN_TOP(\scff_Wires[116] ),
    .SC_OUT_BOT(\scff_Wires[117] ),
    .Test_en_E_in(\Test_enWires[97] ),
    .Test_en_E_out(\Test_enWires[98] ),
    .Test_en_W_in(\Test_enWires[97] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[46] ),
    .ccff_head(cby_1__1__45_ccff_tail),
    .ccff_tail(grid_clb_53_ccff_tail),
    .clk_0_N_in(\clk_1_wires[101] ),
    .clk_0_S_in(\clk_1_wires[101] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[189] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[101] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[101] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[188] ),
    .right_width_0_height_0__pin_16_(cby_1__1__53_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__53_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__53_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__53_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__53_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__53_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__53_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__53_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__53_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__53_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__53_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__53_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__53_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__53_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__53_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__53_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_53_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_53_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_53_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_53_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_53_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_53_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_53_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_53_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_53_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_53_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_53_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_53_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_53_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_53_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_53_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_53_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__47_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__47_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__47_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__47_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__47_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__47_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__47_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__47_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__47_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[47] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_53_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_53_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_53_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_53_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_53_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_53_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_53_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_53_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_53_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_53_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_53_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_53_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__47_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_53_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_53_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_53_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_53_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__47_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__47_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__47_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__47_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__47_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__47_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__7_ (.SC_IN_TOP(\scff_Wires[114] ),
    .SC_OUT_BOT(\scff_Wires[115] ),
    .Test_en_E_in(\Test_enWires[111] ),
    .Test_en_E_out(\Test_enWires[112] ),
    .Test_en_W_in(\Test_enWires[111] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[47] ),
    .ccff_head(cby_1__1__46_ccff_tail),
    .ccff_tail(grid_clb_54_ccff_tail),
    .clk_0_N_in(\clk_1_wires[109] ),
    .clk_0_S_in(\clk_1_wires[109] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[192] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[109] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[109] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[191] ),
    .right_width_0_height_0__pin_16_(cby_1__1__54_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__54_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__54_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__54_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__54_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__54_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__54_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__54_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__54_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__54_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__54_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__54_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__54_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__54_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__54_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__54_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_54_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_54_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_54_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_54_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_54_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_54_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_54_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_54_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_54_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_54_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_54_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_54_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_54_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_54_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_54_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_54_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__48_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__48_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__48_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__48_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__48_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__48_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__48_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__48_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__48_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[48] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_54_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_54_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_54_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_54_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_54_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_54_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_54_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_54_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_54_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_54_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_54_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_54_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__48_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_54_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_54_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_54_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_54_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__48_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__48_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__48_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__48_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__48_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__48_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_7__8_ (.SC_IN_TOP(\scff_Wires[112] ),
    .SC_OUT_BOT(\scff_Wires[113] ),
    .Test_en_E_in(\Test_enWires[125] ),
    .Test_en_E_out(\Test_enWires[126] ),
    .Test_en_W_in(\Test_enWires[125] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[48] ),
    .ccff_head(cby_1__1__47_ccff_tail),
    .ccff_tail(grid_clb_55_ccff_tail),
    .clk_0_N_in(\clk_1_wires[108] ),
    .clk_0_S_in(\clk_1_wires[108] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[195] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[108] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[197] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[108] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[194] ),
    .right_width_0_height_0__pin_16_(cby_1__1__55_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_1__1__55_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_1__1__55_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_1__1__55_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_1__1__55_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_1__1__55_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_1__1__55_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_1__1__55_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_1__1__55_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_1__1__55_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_1__1__55_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_1__1__55_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_1__1__55_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_1__1__55_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_1__1__55_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_1__1__55_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_55_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_55_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_55_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_55_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_55_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_55_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_55_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_55_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_55_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_55_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_55_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_55_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_55_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_55_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_55_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_55_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__6_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__6_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__6_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__6_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__6_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__6_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__6_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__6_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__6_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[6] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_55_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_55_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_55_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_55_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_55_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_55_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_55_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_55_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_55_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_55_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_55_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_55_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__6_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_55_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_55_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_55_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_55_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__6_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__6_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__6_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__6_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__6_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__6_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__1_ (.SC_IN_TOP(\scff_Wires[131] ),
    .SC_OUT_TOP(\scff_Wires[132] ),
    .Test_en_E_in(\Test_enWires[29] ),
    .Test_en_W_in(\Test_enWires[29] ),
    .ccff_head(cby_1__1__48_ccff_tail),
    .ccff_tail(grid_clb_56_ccff_tail),
    .clk_0_N_in(\clk_1_wires[90] ),
    .clk_0_S_in(\clk_1_wires[90] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[200] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[90] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[90] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[199] ),
    .right_width_0_height_0__pin_16_(cby_8__1__0_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__0_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__0_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__0_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__0_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__0_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__0_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__0_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__0_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__0_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__0_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__0_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__0_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__0_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__0_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__0_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_56_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_56_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_56_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_56_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_56_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_56_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_56_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_56_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_56_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_56_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_56_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_56_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_56_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_56_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_56_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_56_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__49_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__49_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__49_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__49_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__49_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__49_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__49_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__49_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__49_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[49] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_56_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_56_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_56_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_56_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_56_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_56_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_56_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_56_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_56_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_56_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_56_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_56_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__49_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_56_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_56_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_56_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_56_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__49_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__49_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__49_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__49_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__49_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__49_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__2_ (.SC_IN_TOP(\scff_Wires[133] ),
    .SC_OUT_TOP(\scff_Wires[134] ),
    .Test_en_E_in(\Test_enWires[43] ),
    .Test_en_W_in(\Test_enWires[43] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[49] ),
    .ccff_head(cby_1__1__49_ccff_tail),
    .ccff_tail(grid_clb_57_ccff_tail),
    .clk_0_N_in(\clk_1_wires[89] ),
    .clk_0_S_in(\clk_1_wires[89] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[203] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[89] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[89] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[202] ),
    .right_width_0_height_0__pin_16_(cby_8__1__1_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__1_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__1_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__1_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__1_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__1_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__1_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__1_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__1_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__1_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__1_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__1_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__1_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__1_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__1_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__1_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_57_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_57_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_57_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_57_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_57_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_57_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_57_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_57_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_57_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_57_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_57_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_57_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_57_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_57_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_57_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_57_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__50_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__50_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__50_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__50_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__50_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__50_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__50_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__50_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__50_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[50] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_57_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_57_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_57_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_57_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_57_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_57_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_57_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_57_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_57_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_57_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_57_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_57_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__50_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_57_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_57_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_57_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_57_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__50_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__50_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__50_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__50_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__50_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__50_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__3_ (.SC_IN_TOP(\scff_Wires[135] ),
    .SC_OUT_TOP(\scff_Wires[136] ),
    .Test_en_E_in(\Test_enWires[57] ),
    .Test_en_W_in(\Test_enWires[57] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[50] ),
    .ccff_head(cby_1__1__50_ccff_tail),
    .ccff_tail(grid_clb_58_ccff_tail),
    .clk_0_N_in(\clk_1_wires[97] ),
    .clk_0_S_in(\clk_1_wires[97] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[206] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[97] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[97] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[205] ),
    .right_width_0_height_0__pin_16_(cby_8__1__2_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__2_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__2_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__2_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__2_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__2_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__2_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__2_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__2_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__2_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__2_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__2_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__2_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__2_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__2_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__2_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_58_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_58_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_58_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_58_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_58_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_58_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_58_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_58_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_58_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_58_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_58_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_58_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_58_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_58_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_58_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_58_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__51_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__51_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__51_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__51_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__51_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__51_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__51_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__51_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__51_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[51] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_58_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_58_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_58_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_58_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_58_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_58_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_58_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_58_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_58_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_58_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_58_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_58_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__51_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_58_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_58_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_58_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_58_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__51_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__51_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__51_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__51_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__51_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__51_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__4_ (.SC_IN_TOP(\scff_Wires[137] ),
    .SC_OUT_TOP(\scff_Wires[138] ),
    .Test_en_E_in(\Test_enWires[71] ),
    .Test_en_W_in(\Test_enWires[71] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[51] ),
    .ccff_head(cby_1__1__51_ccff_tail),
    .ccff_tail(grid_clb_59_ccff_tail),
    .clk_0_N_in(\clk_1_wires[96] ),
    .clk_0_S_in(\clk_1_wires[96] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[209] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[96] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[96] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[208] ),
    .right_width_0_height_0__pin_16_(cby_8__1__3_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__3_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__3_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__3_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__3_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__3_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__3_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__3_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__3_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__3_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__3_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__3_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__3_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__3_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__3_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__3_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_59_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_59_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_59_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_59_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_59_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_59_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_59_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_59_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_59_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_59_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_59_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_59_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_59_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_59_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_59_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_59_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__52_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__52_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__52_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__52_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__52_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__52_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__52_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__52_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__52_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[52] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_59_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_59_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_59_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_59_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_59_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_59_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_59_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_59_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_59_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_59_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_59_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_59_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__52_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_59_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_59_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_59_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_59_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__52_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__52_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__52_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__52_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__52_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__52_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__5_ (.SC_IN_TOP(\scff_Wires[139] ),
    .SC_OUT_TOP(\scff_Wires[140] ),
    .Test_en_E_in(\Test_enWires[85] ),
    .Test_en_W_in(\Test_enWires[85] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[52] ),
    .ccff_head(cby_1__1__52_ccff_tail),
    .ccff_tail(grid_clb_60_ccff_tail),
    .clk_0_N_in(\clk_1_wires[104] ),
    .clk_0_S_in(\clk_1_wires[104] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[212] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[104] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[104] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[211] ),
    .right_width_0_height_0__pin_16_(cby_8__1__4_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__4_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__4_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__4_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__4_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__4_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__4_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__4_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__4_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__4_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__4_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__4_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__4_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__4_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__4_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__4_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_60_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_60_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_60_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_60_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_60_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_60_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_60_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_60_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_60_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_60_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_60_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_60_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_60_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_60_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_60_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_60_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__53_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__53_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__53_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__53_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__53_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__53_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__53_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__53_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__53_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[53] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_60_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_60_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_60_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_60_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_60_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_60_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_60_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_60_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_60_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_60_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_60_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_60_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__53_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_60_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_60_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_60_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_60_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__53_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__53_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__53_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__53_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__53_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__53_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__6_ (.SC_IN_TOP(\scff_Wires[141] ),
    .SC_OUT_TOP(\scff_Wires[142] ),
    .Test_en_E_in(\Test_enWires[99] ),
    .Test_en_W_in(\Test_enWires[99] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[53] ),
    .ccff_head(cby_1__1__53_ccff_tail),
    .ccff_tail(grid_clb_61_ccff_tail),
    .clk_0_N_in(\clk_1_wires[103] ),
    .clk_0_S_in(\clk_1_wires[103] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[215] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[103] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[103] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[214] ),
    .right_width_0_height_0__pin_16_(cby_8__1__5_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__5_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__5_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__5_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__5_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__5_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__5_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__5_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__5_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__5_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__5_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__5_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__5_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__5_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__5_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__5_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_61_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_61_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_61_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_61_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_61_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_61_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_61_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_61_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_61_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_61_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_61_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_61_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_61_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_61_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_61_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_61_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__54_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__54_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__54_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__54_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__54_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__54_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__54_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__54_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__54_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[54] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_61_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_61_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_61_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_61_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_61_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_61_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_61_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_61_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_61_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_61_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_61_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_61_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__54_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_61_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_61_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_61_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_61_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__54_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__54_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__54_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__54_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__54_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__54_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__7_ (.SC_IN_TOP(\scff_Wires[143] ),
    .SC_OUT_TOP(\scff_Wires[144] ),
    .Test_en_E_in(\Test_enWires[113] ),
    .Test_en_W_in(\Test_enWires[113] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[54] ),
    .ccff_head(cby_1__1__54_ccff_tail),
    .ccff_tail(grid_clb_62_ccff_tail),
    .clk_0_N_in(\clk_1_wires[111] ),
    .clk_0_S_in(\clk_1_wires[111] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[218] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[111] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[111] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[217] ),
    .right_width_0_height_0__pin_16_(cby_8__1__6_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__6_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__6_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__6_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__6_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__6_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__6_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__6_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__6_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__6_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__6_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__6_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__6_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__6_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__6_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__6_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_62_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_62_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_62_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_62_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_62_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_62_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_62_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_62_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_62_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_62_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_62_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_62_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_62_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_62_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_62_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_62_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__1__55_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__1__55_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__1__55_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__1__55_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__1__55_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__1__55_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__1__55_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__1__55_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__1__55_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\regout_feedthrough_wires[55] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_62_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_62_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_62_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_62_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_62_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_62_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_62_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_62_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_62_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_62_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_62_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_62_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__1__55_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_62_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_62_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_62_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_62_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__1__55_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__1__55_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__1__55_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__1__55_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__1__55_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__1__55_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 grid_clb grid_clb_8__8_ (.SC_IN_TOP(\scff_Wires[145] ),
    .SC_OUT_TOP(\scff_Wires[146] ),
    .Test_en_E_in(\Test_enWires[127] ),
    .Test_en_W_in(\Test_enWires[127] ),
    .bottom_width_0_height_0__pin_50_(\regin_feedthrough_wires[55] ),
    .ccff_head(cby_1__1__55_ccff_tail),
    .ccff_tail(grid_clb_63_ccff_tail),
    .clk_0_N_in(\clk_1_wires[110] ),
    .clk_0_S_in(\clk_1_wires[110] ),
    .prog_clk_0_E_out(\prog_clk_0_wires[221] ),
    .prog_clk_0_N_in(\prog_clk_1_wires[110] ),
    .prog_clk_0_N_out(\prog_clk_0_wires[223] ),
    .prog_clk_0_S_in(\prog_clk_1_wires[110] ),
    .prog_clk_0_S_out(\prog_clk_0_wires[220] ),
    .right_width_0_height_0__pin_16_(cby_8__1__7_left_grid_pin_16_),
    .right_width_0_height_0__pin_17_(cby_8__1__7_left_grid_pin_17_),
    .right_width_0_height_0__pin_18_(cby_8__1__7_left_grid_pin_18_),
    .right_width_0_height_0__pin_19_(cby_8__1__7_left_grid_pin_19_),
    .right_width_0_height_0__pin_20_(cby_8__1__7_left_grid_pin_20_),
    .right_width_0_height_0__pin_21_(cby_8__1__7_left_grid_pin_21_),
    .right_width_0_height_0__pin_22_(cby_8__1__7_left_grid_pin_22_),
    .right_width_0_height_0__pin_23_(cby_8__1__7_left_grid_pin_23_),
    .right_width_0_height_0__pin_24_(cby_8__1__7_left_grid_pin_24_),
    .right_width_0_height_0__pin_25_(cby_8__1__7_left_grid_pin_25_),
    .right_width_0_height_0__pin_26_(cby_8__1__7_left_grid_pin_26_),
    .right_width_0_height_0__pin_27_(cby_8__1__7_left_grid_pin_27_),
    .right_width_0_height_0__pin_28_(cby_8__1__7_left_grid_pin_28_),
    .right_width_0_height_0__pin_29_(cby_8__1__7_left_grid_pin_29_),
    .right_width_0_height_0__pin_30_(cby_8__1__7_left_grid_pin_30_),
    .right_width_0_height_0__pin_31_(cby_8__1__7_left_grid_pin_31_),
    .right_width_0_height_0__pin_42_lower(grid_clb_63_right_width_0_height_0__pin_42_lower),
    .right_width_0_height_0__pin_42_upper(grid_clb_63_right_width_0_height_0__pin_42_upper),
    .right_width_0_height_0__pin_43_lower(grid_clb_63_right_width_0_height_0__pin_43_lower),
    .right_width_0_height_0__pin_43_upper(grid_clb_63_right_width_0_height_0__pin_43_upper),
    .right_width_0_height_0__pin_44_lower(grid_clb_63_right_width_0_height_0__pin_44_lower),
    .right_width_0_height_0__pin_44_upper(grid_clb_63_right_width_0_height_0__pin_44_upper),
    .right_width_0_height_0__pin_45_lower(grid_clb_63_right_width_0_height_0__pin_45_lower),
    .right_width_0_height_0__pin_45_upper(grid_clb_63_right_width_0_height_0__pin_45_upper),
    .right_width_0_height_0__pin_46_lower(grid_clb_63_right_width_0_height_0__pin_46_lower),
    .right_width_0_height_0__pin_46_upper(grid_clb_63_right_width_0_height_0__pin_46_upper),
    .right_width_0_height_0__pin_47_lower(grid_clb_63_right_width_0_height_0__pin_47_lower),
    .right_width_0_height_0__pin_47_upper(grid_clb_63_right_width_0_height_0__pin_47_upper),
    .right_width_0_height_0__pin_48_lower(grid_clb_63_right_width_0_height_0__pin_48_lower),
    .right_width_0_height_0__pin_48_upper(grid_clb_63_right_width_0_height_0__pin_48_upper),
    .right_width_0_height_0__pin_49_lower(grid_clb_63_right_width_0_height_0__pin_49_lower),
    .right_width_0_height_0__pin_49_upper(grid_clb_63_right_width_0_height_0__pin_49_upper),
    .top_width_0_height_0__pin_0_(cbx_1__8__7_bottom_grid_pin_0_),
    .top_width_0_height_0__pin_10_(cbx_1__8__7_bottom_grid_pin_10_),
    .top_width_0_height_0__pin_11_(cbx_1__8__7_bottom_grid_pin_11_),
    .top_width_0_height_0__pin_12_(cbx_1__8__7_bottom_grid_pin_12_),
    .top_width_0_height_0__pin_13_(cbx_1__8__7_bottom_grid_pin_13_),
    .top_width_0_height_0__pin_14_(cbx_1__8__7_bottom_grid_pin_14_),
    .top_width_0_height_0__pin_15_(cbx_1__8__7_bottom_grid_pin_15_),
    .top_width_0_height_0__pin_1_(cbx_1__8__7_bottom_grid_pin_1_),
    .top_width_0_height_0__pin_2_(cbx_1__8__7_bottom_grid_pin_2_),
    .top_width_0_height_0__pin_32_(\logic_zero_tie[7] ),
    .top_width_0_height_0__pin_34_lower(grid_clb_63_top_width_0_height_0__pin_34_lower),
    .top_width_0_height_0__pin_34_upper(grid_clb_63_top_width_0_height_0__pin_34_upper),
    .top_width_0_height_0__pin_35_lower(grid_clb_63_top_width_0_height_0__pin_35_lower),
    .top_width_0_height_0__pin_35_upper(grid_clb_63_top_width_0_height_0__pin_35_upper),
    .top_width_0_height_0__pin_36_lower(grid_clb_63_top_width_0_height_0__pin_36_lower),
    .top_width_0_height_0__pin_36_upper(grid_clb_63_top_width_0_height_0__pin_36_upper),
    .top_width_0_height_0__pin_37_lower(grid_clb_63_top_width_0_height_0__pin_37_lower),
    .top_width_0_height_0__pin_37_upper(grid_clb_63_top_width_0_height_0__pin_37_upper),
    .top_width_0_height_0__pin_38_lower(grid_clb_63_top_width_0_height_0__pin_38_lower),
    .top_width_0_height_0__pin_38_upper(grid_clb_63_top_width_0_height_0__pin_38_upper),
    .top_width_0_height_0__pin_39_lower(grid_clb_63_top_width_0_height_0__pin_39_lower),
    .top_width_0_height_0__pin_39_upper(grid_clb_63_top_width_0_height_0__pin_39_upper),
    .top_width_0_height_0__pin_3_(cbx_1__8__7_bottom_grid_pin_3_),
    .top_width_0_height_0__pin_40_lower(grid_clb_63_top_width_0_height_0__pin_40_lower),
    .top_width_0_height_0__pin_40_upper(grid_clb_63_top_width_0_height_0__pin_40_upper),
    .top_width_0_height_0__pin_41_lower(grid_clb_63_top_width_0_height_0__pin_41_lower),
    .top_width_0_height_0__pin_41_upper(grid_clb_63_top_width_0_height_0__pin_41_upper),
    .top_width_0_height_0__pin_4_(cbx_1__8__7_bottom_grid_pin_4_),
    .top_width_0_height_0__pin_5_(cbx_1__8__7_bottom_grid_pin_5_),
    .top_width_0_height_0__pin_6_(cbx_1__8__7_bottom_grid_pin_6_),
    .top_width_0_height_0__pin_7_(cbx_1__8__7_bottom_grid_pin_7_),
    .top_width_0_height_0__pin_8_(cbx_1__8__7_bottom_grid_pin_8_),
    .top_width_0_height_0__pin_9_(cbx_1__8__7_bottom_grid_pin_9_),
    .VPWR(VPWR),
    .VGND(VGND));
 sb_0__0_ sb_0__0_ (.ccff_head(grid_io_bottom_7_ccff_tail),
    .ccff_tail(ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[5] ),
    .right_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__0__0_chanx_left_out[0] ,
    \cbx_1__0__0_chanx_left_out[1] ,
    \cbx_1__0__0_chanx_left_out[2] ,
    \cbx_1__0__0_chanx_left_out[3] ,
    \cbx_1__0__0_chanx_left_out[4] ,
    \cbx_1__0__0_chanx_left_out[5] ,
    \cbx_1__0__0_chanx_left_out[6] ,
    \cbx_1__0__0_chanx_left_out[7] ,
    \cbx_1__0__0_chanx_left_out[8] ,
    \cbx_1__0__0_chanx_left_out[9] ,
    \cbx_1__0__0_chanx_left_out[10] ,
    \cbx_1__0__0_chanx_left_out[11] ,
    \cbx_1__0__0_chanx_left_out[12] ,
    \cbx_1__0__0_chanx_left_out[13] ,
    \cbx_1__0__0_chanx_left_out[14] ,
    \cbx_1__0__0_chanx_left_out[15] ,
    \cbx_1__0__0_chanx_left_out[16] ,
    \cbx_1__0__0_chanx_left_out[17] ,
    \cbx_1__0__0_chanx_left_out[18] ,
    \cbx_1__0__0_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__0__0_chanx_right_out[0] ,
    \sb_0__0__0_chanx_right_out[1] ,
    \sb_0__0__0_chanx_right_out[2] ,
    \sb_0__0__0_chanx_right_out[3] ,
    \sb_0__0__0_chanx_right_out[4] ,
    \sb_0__0__0_chanx_right_out[5] ,
    \sb_0__0__0_chanx_right_out[6] ,
    \sb_0__0__0_chanx_right_out[7] ,
    \sb_0__0__0_chanx_right_out[8] ,
    \sb_0__0__0_chanx_right_out[9] ,
    \sb_0__0__0_chanx_right_out[10] ,
    \sb_0__0__0_chanx_right_out[11] ,
    \sb_0__0__0_chanx_right_out[12] ,
    \sb_0__0__0_chanx_right_out[13] ,
    \sb_0__0__0_chanx_right_out[14] ,
    \sb_0__0__0_chanx_right_out[15] ,
    \sb_0__0__0_chanx_right_out[16] ,
    \sb_0__0__0_chanx_right_out[17] ,
    \sb_0__0__0_chanx_right_out[18] ,
    \sb_0__0__0_chanx_right_out[19] }),
    .chany_top_in({\cby_0__1__0_chany_bottom_out[0] ,
    \cby_0__1__0_chany_bottom_out[1] ,
    \cby_0__1__0_chany_bottom_out[2] ,
    \cby_0__1__0_chany_bottom_out[3] ,
    \cby_0__1__0_chany_bottom_out[4] ,
    \cby_0__1__0_chany_bottom_out[5] ,
    \cby_0__1__0_chany_bottom_out[6] ,
    \cby_0__1__0_chany_bottom_out[7] ,
    \cby_0__1__0_chany_bottom_out[8] ,
    \cby_0__1__0_chany_bottom_out[9] ,
    \cby_0__1__0_chany_bottom_out[10] ,
    \cby_0__1__0_chany_bottom_out[11] ,
    \cby_0__1__0_chany_bottom_out[12] ,
    \cby_0__1__0_chany_bottom_out[13] ,
    \cby_0__1__0_chany_bottom_out[14] ,
    \cby_0__1__0_chany_bottom_out[15] ,
    \cby_0__1__0_chany_bottom_out[16] ,
    \cby_0__1__0_chany_bottom_out[17] ,
    \cby_0__1__0_chany_bottom_out[18] ,
    \cby_0__1__0_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__0__0_chany_top_out[0] ,
    \sb_0__0__0_chany_top_out[1] ,
    \sb_0__0__0_chany_top_out[2] ,
    \sb_0__0__0_chany_top_out[3] ,
    \sb_0__0__0_chany_top_out[4] ,
    \sb_0__0__0_chany_top_out[5] ,
    \sb_0__0__0_chany_top_out[6] ,
    \sb_0__0__0_chany_top_out[7] ,
    \sb_0__0__0_chany_top_out[8] ,
    \sb_0__0__0_chany_top_out[9] ,
    \sb_0__0__0_chany_top_out[10] ,
    \sb_0__0__0_chany_top_out[11] ,
    \sb_0__0__0_chany_top_out[12] ,
    \sb_0__0__0_chany_top_out[13] ,
    \sb_0__0__0_chany_top_out[14] ,
    \sb_0__0__0_chany_top_out[15] ,
    \sb_0__0__0_chany_top_out[16] ,
    \sb_0__0__0_chany_top_out[17] ,
    \sb_0__0__0_chany_top_out[18] ,
    \sb_0__0__0_chany_top_out[19] }));
 sb_0__1_ sb_0__1_ (.bottom_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_upper),
    .ccff_head(cbx_1__1__0_ccff_tail),
    .ccff_tail(sb_0__1__0_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[4] ),
    .right_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__1__0_chanx_left_out[0] ,
    \cbx_1__1__0_chanx_left_out[1] ,
    \cbx_1__1__0_chanx_left_out[2] ,
    \cbx_1__1__0_chanx_left_out[3] ,
    \cbx_1__1__0_chanx_left_out[4] ,
    \cbx_1__1__0_chanx_left_out[5] ,
    \cbx_1__1__0_chanx_left_out[6] ,
    \cbx_1__1__0_chanx_left_out[7] ,
    \cbx_1__1__0_chanx_left_out[8] ,
    \cbx_1__1__0_chanx_left_out[9] ,
    \cbx_1__1__0_chanx_left_out[10] ,
    \cbx_1__1__0_chanx_left_out[11] ,
    \cbx_1__1__0_chanx_left_out[12] ,
    \cbx_1__1__0_chanx_left_out[13] ,
    \cbx_1__1__0_chanx_left_out[14] ,
    \cbx_1__1__0_chanx_left_out[15] ,
    \cbx_1__1__0_chanx_left_out[16] ,
    \cbx_1__1__0_chanx_left_out[17] ,
    \cbx_1__1__0_chanx_left_out[18] ,
    \cbx_1__1__0_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__1__0_chanx_right_out[0] ,
    \sb_0__1__0_chanx_right_out[1] ,
    \sb_0__1__0_chanx_right_out[2] ,
    \sb_0__1__0_chanx_right_out[3] ,
    \sb_0__1__0_chanx_right_out[4] ,
    \sb_0__1__0_chanx_right_out[5] ,
    \sb_0__1__0_chanx_right_out[6] ,
    \sb_0__1__0_chanx_right_out[7] ,
    \sb_0__1__0_chanx_right_out[8] ,
    \sb_0__1__0_chanx_right_out[9] ,
    \sb_0__1__0_chanx_right_out[10] ,
    \sb_0__1__0_chanx_right_out[11] ,
    \sb_0__1__0_chanx_right_out[12] ,
    \sb_0__1__0_chanx_right_out[13] ,
    \sb_0__1__0_chanx_right_out[14] ,
    \sb_0__1__0_chanx_right_out[15] ,
    \sb_0__1__0_chanx_right_out[16] ,
    \sb_0__1__0_chanx_right_out[17] ,
    \sb_0__1__0_chanx_right_out[18] ,
    \sb_0__1__0_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__0_chany_top_out[0] ,
    \cby_0__1__0_chany_top_out[1] ,
    \cby_0__1__0_chany_top_out[2] ,
    \cby_0__1__0_chany_top_out[3] ,
    \cby_0__1__0_chany_top_out[4] ,
    \cby_0__1__0_chany_top_out[5] ,
    \cby_0__1__0_chany_top_out[6] ,
    \cby_0__1__0_chany_top_out[7] ,
    \cby_0__1__0_chany_top_out[8] ,
    \cby_0__1__0_chany_top_out[9] ,
    \cby_0__1__0_chany_top_out[10] ,
    \cby_0__1__0_chany_top_out[11] ,
    \cby_0__1__0_chany_top_out[12] ,
    \cby_0__1__0_chany_top_out[13] ,
    \cby_0__1__0_chany_top_out[14] ,
    \cby_0__1__0_chany_top_out[15] ,
    \cby_0__1__0_chany_top_out[16] ,
    \cby_0__1__0_chany_top_out[17] ,
    \cby_0__1__0_chany_top_out[18] ,
    \cby_0__1__0_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__1__0_chany_bottom_out[0] ,
    \sb_0__1__0_chany_bottom_out[1] ,
    \sb_0__1__0_chany_bottom_out[2] ,
    \sb_0__1__0_chany_bottom_out[3] ,
    \sb_0__1__0_chany_bottom_out[4] ,
    \sb_0__1__0_chany_bottom_out[5] ,
    \sb_0__1__0_chany_bottom_out[6] ,
    \sb_0__1__0_chany_bottom_out[7] ,
    \sb_0__1__0_chany_bottom_out[8] ,
    \sb_0__1__0_chany_bottom_out[9] ,
    \sb_0__1__0_chany_bottom_out[10] ,
    \sb_0__1__0_chany_bottom_out[11] ,
    \sb_0__1__0_chany_bottom_out[12] ,
    \sb_0__1__0_chany_bottom_out[13] ,
    \sb_0__1__0_chany_bottom_out[14] ,
    \sb_0__1__0_chany_bottom_out[15] ,
    \sb_0__1__0_chany_bottom_out[16] ,
    \sb_0__1__0_chany_bottom_out[17] ,
    \sb_0__1__0_chany_bottom_out[18] ,
    \sb_0__1__0_chany_bottom_out[19] }),
    .chany_top_in({\cby_0__1__1_chany_bottom_out[0] ,
    \cby_0__1__1_chany_bottom_out[1] ,
    \cby_0__1__1_chany_bottom_out[2] ,
    \cby_0__1__1_chany_bottom_out[3] ,
    \cby_0__1__1_chany_bottom_out[4] ,
    \cby_0__1__1_chany_bottom_out[5] ,
    \cby_0__1__1_chany_bottom_out[6] ,
    \cby_0__1__1_chany_bottom_out[7] ,
    \cby_0__1__1_chany_bottom_out[8] ,
    \cby_0__1__1_chany_bottom_out[9] ,
    \cby_0__1__1_chany_bottom_out[10] ,
    \cby_0__1__1_chany_bottom_out[11] ,
    \cby_0__1__1_chany_bottom_out[12] ,
    \cby_0__1__1_chany_bottom_out[13] ,
    \cby_0__1__1_chany_bottom_out[14] ,
    \cby_0__1__1_chany_bottom_out[15] ,
    \cby_0__1__1_chany_bottom_out[16] ,
    \cby_0__1__1_chany_bottom_out[17] ,
    \cby_0__1__1_chany_bottom_out[18] ,
    \cby_0__1__1_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__1__0_chany_top_out[0] ,
    \sb_0__1__0_chany_top_out[1] ,
    \sb_0__1__0_chany_top_out[2] ,
    \sb_0__1__0_chany_top_out[3] ,
    \sb_0__1__0_chany_top_out[4] ,
    \sb_0__1__0_chany_top_out[5] ,
    \sb_0__1__0_chany_top_out[6] ,
    \sb_0__1__0_chany_top_out[7] ,
    \sb_0__1__0_chany_top_out[8] ,
    \sb_0__1__0_chany_top_out[9] ,
    \sb_0__1__0_chany_top_out[10] ,
    \sb_0__1__0_chany_top_out[11] ,
    \sb_0__1__0_chany_top_out[12] ,
    \sb_0__1__0_chany_top_out[13] ,
    \sb_0__1__0_chany_top_out[14] ,
    \sb_0__1__0_chany_top_out[15] ,
    \sb_0__1__0_chany_top_out[16] ,
    \sb_0__1__0_chany_top_out[17] ,
    \sb_0__1__0_chany_top_out[18] ,
    \sb_0__1__0_chany_top_out[19] }));
 sb_0__1_ sb_0__2_ (.bottom_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_upper),
    .ccff_head(cbx_1__1__1_ccff_tail),
    .ccff_tail(sb_0__1__1_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[10] ),
    .right_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__1__1_chanx_left_out[0] ,
    \cbx_1__1__1_chanx_left_out[1] ,
    \cbx_1__1__1_chanx_left_out[2] ,
    \cbx_1__1__1_chanx_left_out[3] ,
    \cbx_1__1__1_chanx_left_out[4] ,
    \cbx_1__1__1_chanx_left_out[5] ,
    \cbx_1__1__1_chanx_left_out[6] ,
    \cbx_1__1__1_chanx_left_out[7] ,
    \cbx_1__1__1_chanx_left_out[8] ,
    \cbx_1__1__1_chanx_left_out[9] ,
    \cbx_1__1__1_chanx_left_out[10] ,
    \cbx_1__1__1_chanx_left_out[11] ,
    \cbx_1__1__1_chanx_left_out[12] ,
    \cbx_1__1__1_chanx_left_out[13] ,
    \cbx_1__1__1_chanx_left_out[14] ,
    \cbx_1__1__1_chanx_left_out[15] ,
    \cbx_1__1__1_chanx_left_out[16] ,
    \cbx_1__1__1_chanx_left_out[17] ,
    \cbx_1__1__1_chanx_left_out[18] ,
    \cbx_1__1__1_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__1__1_chanx_right_out[0] ,
    \sb_0__1__1_chanx_right_out[1] ,
    \sb_0__1__1_chanx_right_out[2] ,
    \sb_0__1__1_chanx_right_out[3] ,
    \sb_0__1__1_chanx_right_out[4] ,
    \sb_0__1__1_chanx_right_out[5] ,
    \sb_0__1__1_chanx_right_out[6] ,
    \sb_0__1__1_chanx_right_out[7] ,
    \sb_0__1__1_chanx_right_out[8] ,
    \sb_0__1__1_chanx_right_out[9] ,
    \sb_0__1__1_chanx_right_out[10] ,
    \sb_0__1__1_chanx_right_out[11] ,
    \sb_0__1__1_chanx_right_out[12] ,
    \sb_0__1__1_chanx_right_out[13] ,
    \sb_0__1__1_chanx_right_out[14] ,
    \sb_0__1__1_chanx_right_out[15] ,
    \sb_0__1__1_chanx_right_out[16] ,
    \sb_0__1__1_chanx_right_out[17] ,
    \sb_0__1__1_chanx_right_out[18] ,
    \sb_0__1__1_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__1_chany_top_out[0] ,
    \cby_0__1__1_chany_top_out[1] ,
    \cby_0__1__1_chany_top_out[2] ,
    \cby_0__1__1_chany_top_out[3] ,
    \cby_0__1__1_chany_top_out[4] ,
    \cby_0__1__1_chany_top_out[5] ,
    \cby_0__1__1_chany_top_out[6] ,
    \cby_0__1__1_chany_top_out[7] ,
    \cby_0__1__1_chany_top_out[8] ,
    \cby_0__1__1_chany_top_out[9] ,
    \cby_0__1__1_chany_top_out[10] ,
    \cby_0__1__1_chany_top_out[11] ,
    \cby_0__1__1_chany_top_out[12] ,
    \cby_0__1__1_chany_top_out[13] ,
    \cby_0__1__1_chany_top_out[14] ,
    \cby_0__1__1_chany_top_out[15] ,
    \cby_0__1__1_chany_top_out[16] ,
    \cby_0__1__1_chany_top_out[17] ,
    \cby_0__1__1_chany_top_out[18] ,
    \cby_0__1__1_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__1__1_chany_bottom_out[0] ,
    \sb_0__1__1_chany_bottom_out[1] ,
    \sb_0__1__1_chany_bottom_out[2] ,
    \sb_0__1__1_chany_bottom_out[3] ,
    \sb_0__1__1_chany_bottom_out[4] ,
    \sb_0__1__1_chany_bottom_out[5] ,
    \sb_0__1__1_chany_bottom_out[6] ,
    \sb_0__1__1_chany_bottom_out[7] ,
    \sb_0__1__1_chany_bottom_out[8] ,
    \sb_0__1__1_chany_bottom_out[9] ,
    \sb_0__1__1_chany_bottom_out[10] ,
    \sb_0__1__1_chany_bottom_out[11] ,
    \sb_0__1__1_chany_bottom_out[12] ,
    \sb_0__1__1_chany_bottom_out[13] ,
    \sb_0__1__1_chany_bottom_out[14] ,
    \sb_0__1__1_chany_bottom_out[15] ,
    \sb_0__1__1_chany_bottom_out[16] ,
    \sb_0__1__1_chany_bottom_out[17] ,
    \sb_0__1__1_chany_bottom_out[18] ,
    \sb_0__1__1_chany_bottom_out[19] }),
    .chany_top_in({\cby_0__1__2_chany_bottom_out[0] ,
    \cby_0__1__2_chany_bottom_out[1] ,
    \cby_0__1__2_chany_bottom_out[2] ,
    \cby_0__1__2_chany_bottom_out[3] ,
    \cby_0__1__2_chany_bottom_out[4] ,
    \cby_0__1__2_chany_bottom_out[5] ,
    \cby_0__1__2_chany_bottom_out[6] ,
    \cby_0__1__2_chany_bottom_out[7] ,
    \cby_0__1__2_chany_bottom_out[8] ,
    \cby_0__1__2_chany_bottom_out[9] ,
    \cby_0__1__2_chany_bottom_out[10] ,
    \cby_0__1__2_chany_bottom_out[11] ,
    \cby_0__1__2_chany_bottom_out[12] ,
    \cby_0__1__2_chany_bottom_out[13] ,
    \cby_0__1__2_chany_bottom_out[14] ,
    \cby_0__1__2_chany_bottom_out[15] ,
    \cby_0__1__2_chany_bottom_out[16] ,
    \cby_0__1__2_chany_bottom_out[17] ,
    \cby_0__1__2_chany_bottom_out[18] ,
    \cby_0__1__2_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__1__1_chany_top_out[0] ,
    \sb_0__1__1_chany_top_out[1] ,
    \sb_0__1__1_chany_top_out[2] ,
    \sb_0__1__1_chany_top_out[3] ,
    \sb_0__1__1_chany_top_out[4] ,
    \sb_0__1__1_chany_top_out[5] ,
    \sb_0__1__1_chany_top_out[6] ,
    \sb_0__1__1_chany_top_out[7] ,
    \sb_0__1__1_chany_top_out[8] ,
    \sb_0__1__1_chany_top_out[9] ,
    \sb_0__1__1_chany_top_out[10] ,
    \sb_0__1__1_chany_top_out[11] ,
    \sb_0__1__1_chany_top_out[12] ,
    \sb_0__1__1_chany_top_out[13] ,
    \sb_0__1__1_chany_top_out[14] ,
    \sb_0__1__1_chany_top_out[15] ,
    \sb_0__1__1_chany_top_out[16] ,
    \sb_0__1__1_chany_top_out[17] ,
    \sb_0__1__1_chany_top_out[18] ,
    \sb_0__1__1_chany_top_out[19] }));
 sb_0__1_ sb_0__3_ (.bottom_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_upper),
    .ccff_head(cbx_1__1__2_ccff_tail),
    .ccff_tail(sb_0__1__2_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[15] ),
    .right_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__1__2_chanx_left_out[0] ,
    \cbx_1__1__2_chanx_left_out[1] ,
    \cbx_1__1__2_chanx_left_out[2] ,
    \cbx_1__1__2_chanx_left_out[3] ,
    \cbx_1__1__2_chanx_left_out[4] ,
    \cbx_1__1__2_chanx_left_out[5] ,
    \cbx_1__1__2_chanx_left_out[6] ,
    \cbx_1__1__2_chanx_left_out[7] ,
    \cbx_1__1__2_chanx_left_out[8] ,
    \cbx_1__1__2_chanx_left_out[9] ,
    \cbx_1__1__2_chanx_left_out[10] ,
    \cbx_1__1__2_chanx_left_out[11] ,
    \cbx_1__1__2_chanx_left_out[12] ,
    \cbx_1__1__2_chanx_left_out[13] ,
    \cbx_1__1__2_chanx_left_out[14] ,
    \cbx_1__1__2_chanx_left_out[15] ,
    \cbx_1__1__2_chanx_left_out[16] ,
    \cbx_1__1__2_chanx_left_out[17] ,
    \cbx_1__1__2_chanx_left_out[18] ,
    \cbx_1__1__2_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__1__2_chanx_right_out[0] ,
    \sb_0__1__2_chanx_right_out[1] ,
    \sb_0__1__2_chanx_right_out[2] ,
    \sb_0__1__2_chanx_right_out[3] ,
    \sb_0__1__2_chanx_right_out[4] ,
    \sb_0__1__2_chanx_right_out[5] ,
    \sb_0__1__2_chanx_right_out[6] ,
    \sb_0__1__2_chanx_right_out[7] ,
    \sb_0__1__2_chanx_right_out[8] ,
    \sb_0__1__2_chanx_right_out[9] ,
    \sb_0__1__2_chanx_right_out[10] ,
    \sb_0__1__2_chanx_right_out[11] ,
    \sb_0__1__2_chanx_right_out[12] ,
    \sb_0__1__2_chanx_right_out[13] ,
    \sb_0__1__2_chanx_right_out[14] ,
    \sb_0__1__2_chanx_right_out[15] ,
    \sb_0__1__2_chanx_right_out[16] ,
    \sb_0__1__2_chanx_right_out[17] ,
    \sb_0__1__2_chanx_right_out[18] ,
    \sb_0__1__2_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__2_chany_top_out[0] ,
    \cby_0__1__2_chany_top_out[1] ,
    \cby_0__1__2_chany_top_out[2] ,
    \cby_0__1__2_chany_top_out[3] ,
    \cby_0__1__2_chany_top_out[4] ,
    \cby_0__1__2_chany_top_out[5] ,
    \cby_0__1__2_chany_top_out[6] ,
    \cby_0__1__2_chany_top_out[7] ,
    \cby_0__1__2_chany_top_out[8] ,
    \cby_0__1__2_chany_top_out[9] ,
    \cby_0__1__2_chany_top_out[10] ,
    \cby_0__1__2_chany_top_out[11] ,
    \cby_0__1__2_chany_top_out[12] ,
    \cby_0__1__2_chany_top_out[13] ,
    \cby_0__1__2_chany_top_out[14] ,
    \cby_0__1__2_chany_top_out[15] ,
    \cby_0__1__2_chany_top_out[16] ,
    \cby_0__1__2_chany_top_out[17] ,
    \cby_0__1__2_chany_top_out[18] ,
    \cby_0__1__2_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__1__2_chany_bottom_out[0] ,
    \sb_0__1__2_chany_bottom_out[1] ,
    \sb_0__1__2_chany_bottom_out[2] ,
    \sb_0__1__2_chany_bottom_out[3] ,
    \sb_0__1__2_chany_bottom_out[4] ,
    \sb_0__1__2_chany_bottom_out[5] ,
    \sb_0__1__2_chany_bottom_out[6] ,
    \sb_0__1__2_chany_bottom_out[7] ,
    \sb_0__1__2_chany_bottom_out[8] ,
    \sb_0__1__2_chany_bottom_out[9] ,
    \sb_0__1__2_chany_bottom_out[10] ,
    \sb_0__1__2_chany_bottom_out[11] ,
    \sb_0__1__2_chany_bottom_out[12] ,
    \sb_0__1__2_chany_bottom_out[13] ,
    \sb_0__1__2_chany_bottom_out[14] ,
    \sb_0__1__2_chany_bottom_out[15] ,
    \sb_0__1__2_chany_bottom_out[16] ,
    \sb_0__1__2_chany_bottom_out[17] ,
    \sb_0__1__2_chany_bottom_out[18] ,
    \sb_0__1__2_chany_bottom_out[19] }),
    .chany_top_in({\cby_0__1__3_chany_bottom_out[0] ,
    \cby_0__1__3_chany_bottom_out[1] ,
    \cby_0__1__3_chany_bottom_out[2] ,
    \cby_0__1__3_chany_bottom_out[3] ,
    \cby_0__1__3_chany_bottom_out[4] ,
    \cby_0__1__3_chany_bottom_out[5] ,
    \cby_0__1__3_chany_bottom_out[6] ,
    \cby_0__1__3_chany_bottom_out[7] ,
    \cby_0__1__3_chany_bottom_out[8] ,
    \cby_0__1__3_chany_bottom_out[9] ,
    \cby_0__1__3_chany_bottom_out[10] ,
    \cby_0__1__3_chany_bottom_out[11] ,
    \cby_0__1__3_chany_bottom_out[12] ,
    \cby_0__1__3_chany_bottom_out[13] ,
    \cby_0__1__3_chany_bottom_out[14] ,
    \cby_0__1__3_chany_bottom_out[15] ,
    \cby_0__1__3_chany_bottom_out[16] ,
    \cby_0__1__3_chany_bottom_out[17] ,
    \cby_0__1__3_chany_bottom_out[18] ,
    \cby_0__1__3_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__1__2_chany_top_out[0] ,
    \sb_0__1__2_chany_top_out[1] ,
    \sb_0__1__2_chany_top_out[2] ,
    \sb_0__1__2_chany_top_out[3] ,
    \sb_0__1__2_chany_top_out[4] ,
    \sb_0__1__2_chany_top_out[5] ,
    \sb_0__1__2_chany_top_out[6] ,
    \sb_0__1__2_chany_top_out[7] ,
    \sb_0__1__2_chany_top_out[8] ,
    \sb_0__1__2_chany_top_out[9] ,
    \sb_0__1__2_chany_top_out[10] ,
    \sb_0__1__2_chany_top_out[11] ,
    \sb_0__1__2_chany_top_out[12] ,
    \sb_0__1__2_chany_top_out[13] ,
    \sb_0__1__2_chany_top_out[14] ,
    \sb_0__1__2_chany_top_out[15] ,
    \sb_0__1__2_chany_top_out[16] ,
    \sb_0__1__2_chany_top_out[17] ,
    \sb_0__1__2_chany_top_out[18] ,
    \sb_0__1__2_chany_top_out[19] }));
 sb_0__1_ sb_0__4_ (.bottom_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_upper),
    .ccff_head(cbx_1__1__3_ccff_tail),
    .ccff_tail(sb_0__1__3_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[20] ),
    .right_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__1__3_chanx_left_out[0] ,
    \cbx_1__1__3_chanx_left_out[1] ,
    \cbx_1__1__3_chanx_left_out[2] ,
    \cbx_1__1__3_chanx_left_out[3] ,
    \cbx_1__1__3_chanx_left_out[4] ,
    \cbx_1__1__3_chanx_left_out[5] ,
    \cbx_1__1__3_chanx_left_out[6] ,
    \cbx_1__1__3_chanx_left_out[7] ,
    \cbx_1__1__3_chanx_left_out[8] ,
    \cbx_1__1__3_chanx_left_out[9] ,
    \cbx_1__1__3_chanx_left_out[10] ,
    \cbx_1__1__3_chanx_left_out[11] ,
    \cbx_1__1__3_chanx_left_out[12] ,
    \cbx_1__1__3_chanx_left_out[13] ,
    \cbx_1__1__3_chanx_left_out[14] ,
    \cbx_1__1__3_chanx_left_out[15] ,
    \cbx_1__1__3_chanx_left_out[16] ,
    \cbx_1__1__3_chanx_left_out[17] ,
    \cbx_1__1__3_chanx_left_out[18] ,
    \cbx_1__1__3_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__1__3_chanx_right_out[0] ,
    \sb_0__1__3_chanx_right_out[1] ,
    \sb_0__1__3_chanx_right_out[2] ,
    \sb_0__1__3_chanx_right_out[3] ,
    \sb_0__1__3_chanx_right_out[4] ,
    \sb_0__1__3_chanx_right_out[5] ,
    \sb_0__1__3_chanx_right_out[6] ,
    \sb_0__1__3_chanx_right_out[7] ,
    \sb_0__1__3_chanx_right_out[8] ,
    \sb_0__1__3_chanx_right_out[9] ,
    \sb_0__1__3_chanx_right_out[10] ,
    \sb_0__1__3_chanx_right_out[11] ,
    \sb_0__1__3_chanx_right_out[12] ,
    \sb_0__1__3_chanx_right_out[13] ,
    \sb_0__1__3_chanx_right_out[14] ,
    \sb_0__1__3_chanx_right_out[15] ,
    \sb_0__1__3_chanx_right_out[16] ,
    \sb_0__1__3_chanx_right_out[17] ,
    \sb_0__1__3_chanx_right_out[18] ,
    \sb_0__1__3_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__3_chany_top_out[0] ,
    \cby_0__1__3_chany_top_out[1] ,
    \cby_0__1__3_chany_top_out[2] ,
    \cby_0__1__3_chany_top_out[3] ,
    \cby_0__1__3_chany_top_out[4] ,
    \cby_0__1__3_chany_top_out[5] ,
    \cby_0__1__3_chany_top_out[6] ,
    \cby_0__1__3_chany_top_out[7] ,
    \cby_0__1__3_chany_top_out[8] ,
    \cby_0__1__3_chany_top_out[9] ,
    \cby_0__1__3_chany_top_out[10] ,
    \cby_0__1__3_chany_top_out[11] ,
    \cby_0__1__3_chany_top_out[12] ,
    \cby_0__1__3_chany_top_out[13] ,
    \cby_0__1__3_chany_top_out[14] ,
    \cby_0__1__3_chany_top_out[15] ,
    \cby_0__1__3_chany_top_out[16] ,
    \cby_0__1__3_chany_top_out[17] ,
    \cby_0__1__3_chany_top_out[18] ,
    \cby_0__1__3_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__1__3_chany_bottom_out[0] ,
    \sb_0__1__3_chany_bottom_out[1] ,
    \sb_0__1__3_chany_bottom_out[2] ,
    \sb_0__1__3_chany_bottom_out[3] ,
    \sb_0__1__3_chany_bottom_out[4] ,
    \sb_0__1__3_chany_bottom_out[5] ,
    \sb_0__1__3_chany_bottom_out[6] ,
    \sb_0__1__3_chany_bottom_out[7] ,
    \sb_0__1__3_chany_bottom_out[8] ,
    \sb_0__1__3_chany_bottom_out[9] ,
    \sb_0__1__3_chany_bottom_out[10] ,
    \sb_0__1__3_chany_bottom_out[11] ,
    \sb_0__1__3_chany_bottom_out[12] ,
    \sb_0__1__3_chany_bottom_out[13] ,
    \sb_0__1__3_chany_bottom_out[14] ,
    \sb_0__1__3_chany_bottom_out[15] ,
    \sb_0__1__3_chany_bottom_out[16] ,
    \sb_0__1__3_chany_bottom_out[17] ,
    \sb_0__1__3_chany_bottom_out[18] ,
    \sb_0__1__3_chany_bottom_out[19] }),
    .chany_top_in({\cby_0__1__4_chany_bottom_out[0] ,
    \cby_0__1__4_chany_bottom_out[1] ,
    \cby_0__1__4_chany_bottom_out[2] ,
    \cby_0__1__4_chany_bottom_out[3] ,
    \cby_0__1__4_chany_bottom_out[4] ,
    \cby_0__1__4_chany_bottom_out[5] ,
    \cby_0__1__4_chany_bottom_out[6] ,
    \cby_0__1__4_chany_bottom_out[7] ,
    \cby_0__1__4_chany_bottom_out[8] ,
    \cby_0__1__4_chany_bottom_out[9] ,
    \cby_0__1__4_chany_bottom_out[10] ,
    \cby_0__1__4_chany_bottom_out[11] ,
    \cby_0__1__4_chany_bottom_out[12] ,
    \cby_0__1__4_chany_bottom_out[13] ,
    \cby_0__1__4_chany_bottom_out[14] ,
    \cby_0__1__4_chany_bottom_out[15] ,
    \cby_0__1__4_chany_bottom_out[16] ,
    \cby_0__1__4_chany_bottom_out[17] ,
    \cby_0__1__4_chany_bottom_out[18] ,
    \cby_0__1__4_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__1__3_chany_top_out[0] ,
    \sb_0__1__3_chany_top_out[1] ,
    \sb_0__1__3_chany_top_out[2] ,
    \sb_0__1__3_chany_top_out[3] ,
    \sb_0__1__3_chany_top_out[4] ,
    \sb_0__1__3_chany_top_out[5] ,
    \sb_0__1__3_chany_top_out[6] ,
    \sb_0__1__3_chany_top_out[7] ,
    \sb_0__1__3_chany_top_out[8] ,
    \sb_0__1__3_chany_top_out[9] ,
    \sb_0__1__3_chany_top_out[10] ,
    \sb_0__1__3_chany_top_out[11] ,
    \sb_0__1__3_chany_top_out[12] ,
    \sb_0__1__3_chany_top_out[13] ,
    \sb_0__1__3_chany_top_out[14] ,
    \sb_0__1__3_chany_top_out[15] ,
    \sb_0__1__3_chany_top_out[16] ,
    \sb_0__1__3_chany_top_out[17] ,
    \sb_0__1__3_chany_top_out[18] ,
    \sb_0__1__3_chany_top_out[19] }));
 sb_0__1_ sb_0__5_ (.bottom_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_upper),
    .ccff_head(cbx_1__1__4_ccff_tail),
    .ccff_tail(sb_0__1__4_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[25] ),
    .right_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__1__4_chanx_left_out[0] ,
    \cbx_1__1__4_chanx_left_out[1] ,
    \cbx_1__1__4_chanx_left_out[2] ,
    \cbx_1__1__4_chanx_left_out[3] ,
    \cbx_1__1__4_chanx_left_out[4] ,
    \cbx_1__1__4_chanx_left_out[5] ,
    \cbx_1__1__4_chanx_left_out[6] ,
    \cbx_1__1__4_chanx_left_out[7] ,
    \cbx_1__1__4_chanx_left_out[8] ,
    \cbx_1__1__4_chanx_left_out[9] ,
    \cbx_1__1__4_chanx_left_out[10] ,
    \cbx_1__1__4_chanx_left_out[11] ,
    \cbx_1__1__4_chanx_left_out[12] ,
    \cbx_1__1__4_chanx_left_out[13] ,
    \cbx_1__1__4_chanx_left_out[14] ,
    \cbx_1__1__4_chanx_left_out[15] ,
    \cbx_1__1__4_chanx_left_out[16] ,
    \cbx_1__1__4_chanx_left_out[17] ,
    \cbx_1__1__4_chanx_left_out[18] ,
    \cbx_1__1__4_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__1__4_chanx_right_out[0] ,
    \sb_0__1__4_chanx_right_out[1] ,
    \sb_0__1__4_chanx_right_out[2] ,
    \sb_0__1__4_chanx_right_out[3] ,
    \sb_0__1__4_chanx_right_out[4] ,
    \sb_0__1__4_chanx_right_out[5] ,
    \sb_0__1__4_chanx_right_out[6] ,
    \sb_0__1__4_chanx_right_out[7] ,
    \sb_0__1__4_chanx_right_out[8] ,
    \sb_0__1__4_chanx_right_out[9] ,
    \sb_0__1__4_chanx_right_out[10] ,
    \sb_0__1__4_chanx_right_out[11] ,
    \sb_0__1__4_chanx_right_out[12] ,
    \sb_0__1__4_chanx_right_out[13] ,
    \sb_0__1__4_chanx_right_out[14] ,
    \sb_0__1__4_chanx_right_out[15] ,
    \sb_0__1__4_chanx_right_out[16] ,
    \sb_0__1__4_chanx_right_out[17] ,
    \sb_0__1__4_chanx_right_out[18] ,
    \sb_0__1__4_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__4_chany_top_out[0] ,
    \cby_0__1__4_chany_top_out[1] ,
    \cby_0__1__4_chany_top_out[2] ,
    \cby_0__1__4_chany_top_out[3] ,
    \cby_0__1__4_chany_top_out[4] ,
    \cby_0__1__4_chany_top_out[5] ,
    \cby_0__1__4_chany_top_out[6] ,
    \cby_0__1__4_chany_top_out[7] ,
    \cby_0__1__4_chany_top_out[8] ,
    \cby_0__1__4_chany_top_out[9] ,
    \cby_0__1__4_chany_top_out[10] ,
    \cby_0__1__4_chany_top_out[11] ,
    \cby_0__1__4_chany_top_out[12] ,
    \cby_0__1__4_chany_top_out[13] ,
    \cby_0__1__4_chany_top_out[14] ,
    \cby_0__1__4_chany_top_out[15] ,
    \cby_0__1__4_chany_top_out[16] ,
    \cby_0__1__4_chany_top_out[17] ,
    \cby_0__1__4_chany_top_out[18] ,
    \cby_0__1__4_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__1__4_chany_bottom_out[0] ,
    \sb_0__1__4_chany_bottom_out[1] ,
    \sb_0__1__4_chany_bottom_out[2] ,
    \sb_0__1__4_chany_bottom_out[3] ,
    \sb_0__1__4_chany_bottom_out[4] ,
    \sb_0__1__4_chany_bottom_out[5] ,
    \sb_0__1__4_chany_bottom_out[6] ,
    \sb_0__1__4_chany_bottom_out[7] ,
    \sb_0__1__4_chany_bottom_out[8] ,
    \sb_0__1__4_chany_bottom_out[9] ,
    \sb_0__1__4_chany_bottom_out[10] ,
    \sb_0__1__4_chany_bottom_out[11] ,
    \sb_0__1__4_chany_bottom_out[12] ,
    \sb_0__1__4_chany_bottom_out[13] ,
    \sb_0__1__4_chany_bottom_out[14] ,
    \sb_0__1__4_chany_bottom_out[15] ,
    \sb_0__1__4_chany_bottom_out[16] ,
    \sb_0__1__4_chany_bottom_out[17] ,
    \sb_0__1__4_chany_bottom_out[18] ,
    \sb_0__1__4_chany_bottom_out[19] }),
    .chany_top_in({\cby_0__1__5_chany_bottom_out[0] ,
    \cby_0__1__5_chany_bottom_out[1] ,
    \cby_0__1__5_chany_bottom_out[2] ,
    \cby_0__1__5_chany_bottom_out[3] ,
    \cby_0__1__5_chany_bottom_out[4] ,
    \cby_0__1__5_chany_bottom_out[5] ,
    \cby_0__1__5_chany_bottom_out[6] ,
    \cby_0__1__5_chany_bottom_out[7] ,
    \cby_0__1__5_chany_bottom_out[8] ,
    \cby_0__1__5_chany_bottom_out[9] ,
    \cby_0__1__5_chany_bottom_out[10] ,
    \cby_0__1__5_chany_bottom_out[11] ,
    \cby_0__1__5_chany_bottom_out[12] ,
    \cby_0__1__5_chany_bottom_out[13] ,
    \cby_0__1__5_chany_bottom_out[14] ,
    \cby_0__1__5_chany_bottom_out[15] ,
    \cby_0__1__5_chany_bottom_out[16] ,
    \cby_0__1__5_chany_bottom_out[17] ,
    \cby_0__1__5_chany_bottom_out[18] ,
    \cby_0__1__5_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__1__4_chany_top_out[0] ,
    \sb_0__1__4_chany_top_out[1] ,
    \sb_0__1__4_chany_top_out[2] ,
    \sb_0__1__4_chany_top_out[3] ,
    \sb_0__1__4_chany_top_out[4] ,
    \sb_0__1__4_chany_top_out[5] ,
    \sb_0__1__4_chany_top_out[6] ,
    \sb_0__1__4_chany_top_out[7] ,
    \sb_0__1__4_chany_top_out[8] ,
    \sb_0__1__4_chany_top_out[9] ,
    \sb_0__1__4_chany_top_out[10] ,
    \sb_0__1__4_chany_top_out[11] ,
    \sb_0__1__4_chany_top_out[12] ,
    \sb_0__1__4_chany_top_out[13] ,
    \sb_0__1__4_chany_top_out[14] ,
    \sb_0__1__4_chany_top_out[15] ,
    \sb_0__1__4_chany_top_out[16] ,
    \sb_0__1__4_chany_top_out[17] ,
    \sb_0__1__4_chany_top_out[18] ,
    \sb_0__1__4_chany_top_out[19] }));
 sb_0__1_ sb_0__6_ (.bottom_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_upper),
    .ccff_head(cbx_1__1__5_ccff_tail),
    .ccff_tail(sb_0__1__5_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[30] ),
    .right_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__1__5_chanx_left_out[0] ,
    \cbx_1__1__5_chanx_left_out[1] ,
    \cbx_1__1__5_chanx_left_out[2] ,
    \cbx_1__1__5_chanx_left_out[3] ,
    \cbx_1__1__5_chanx_left_out[4] ,
    \cbx_1__1__5_chanx_left_out[5] ,
    \cbx_1__1__5_chanx_left_out[6] ,
    \cbx_1__1__5_chanx_left_out[7] ,
    \cbx_1__1__5_chanx_left_out[8] ,
    \cbx_1__1__5_chanx_left_out[9] ,
    \cbx_1__1__5_chanx_left_out[10] ,
    \cbx_1__1__5_chanx_left_out[11] ,
    \cbx_1__1__5_chanx_left_out[12] ,
    \cbx_1__1__5_chanx_left_out[13] ,
    \cbx_1__1__5_chanx_left_out[14] ,
    \cbx_1__1__5_chanx_left_out[15] ,
    \cbx_1__1__5_chanx_left_out[16] ,
    \cbx_1__1__5_chanx_left_out[17] ,
    \cbx_1__1__5_chanx_left_out[18] ,
    \cbx_1__1__5_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__1__5_chanx_right_out[0] ,
    \sb_0__1__5_chanx_right_out[1] ,
    \sb_0__1__5_chanx_right_out[2] ,
    \sb_0__1__5_chanx_right_out[3] ,
    \sb_0__1__5_chanx_right_out[4] ,
    \sb_0__1__5_chanx_right_out[5] ,
    \sb_0__1__5_chanx_right_out[6] ,
    \sb_0__1__5_chanx_right_out[7] ,
    \sb_0__1__5_chanx_right_out[8] ,
    \sb_0__1__5_chanx_right_out[9] ,
    \sb_0__1__5_chanx_right_out[10] ,
    \sb_0__1__5_chanx_right_out[11] ,
    \sb_0__1__5_chanx_right_out[12] ,
    \sb_0__1__5_chanx_right_out[13] ,
    \sb_0__1__5_chanx_right_out[14] ,
    \sb_0__1__5_chanx_right_out[15] ,
    \sb_0__1__5_chanx_right_out[16] ,
    \sb_0__1__5_chanx_right_out[17] ,
    \sb_0__1__5_chanx_right_out[18] ,
    \sb_0__1__5_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__5_chany_top_out[0] ,
    \cby_0__1__5_chany_top_out[1] ,
    \cby_0__1__5_chany_top_out[2] ,
    \cby_0__1__5_chany_top_out[3] ,
    \cby_0__1__5_chany_top_out[4] ,
    \cby_0__1__5_chany_top_out[5] ,
    \cby_0__1__5_chany_top_out[6] ,
    \cby_0__1__5_chany_top_out[7] ,
    \cby_0__1__5_chany_top_out[8] ,
    \cby_0__1__5_chany_top_out[9] ,
    \cby_0__1__5_chany_top_out[10] ,
    \cby_0__1__5_chany_top_out[11] ,
    \cby_0__1__5_chany_top_out[12] ,
    \cby_0__1__5_chany_top_out[13] ,
    \cby_0__1__5_chany_top_out[14] ,
    \cby_0__1__5_chany_top_out[15] ,
    \cby_0__1__5_chany_top_out[16] ,
    \cby_0__1__5_chany_top_out[17] ,
    \cby_0__1__5_chany_top_out[18] ,
    \cby_0__1__5_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__1__5_chany_bottom_out[0] ,
    \sb_0__1__5_chany_bottom_out[1] ,
    \sb_0__1__5_chany_bottom_out[2] ,
    \sb_0__1__5_chany_bottom_out[3] ,
    \sb_0__1__5_chany_bottom_out[4] ,
    \sb_0__1__5_chany_bottom_out[5] ,
    \sb_0__1__5_chany_bottom_out[6] ,
    \sb_0__1__5_chany_bottom_out[7] ,
    \sb_0__1__5_chany_bottom_out[8] ,
    \sb_0__1__5_chany_bottom_out[9] ,
    \sb_0__1__5_chany_bottom_out[10] ,
    \sb_0__1__5_chany_bottom_out[11] ,
    \sb_0__1__5_chany_bottom_out[12] ,
    \sb_0__1__5_chany_bottom_out[13] ,
    \sb_0__1__5_chany_bottom_out[14] ,
    \sb_0__1__5_chany_bottom_out[15] ,
    \sb_0__1__5_chany_bottom_out[16] ,
    \sb_0__1__5_chany_bottom_out[17] ,
    \sb_0__1__5_chany_bottom_out[18] ,
    \sb_0__1__5_chany_bottom_out[19] }),
    .chany_top_in({\cby_0__1__6_chany_bottom_out[0] ,
    \cby_0__1__6_chany_bottom_out[1] ,
    \cby_0__1__6_chany_bottom_out[2] ,
    \cby_0__1__6_chany_bottom_out[3] ,
    \cby_0__1__6_chany_bottom_out[4] ,
    \cby_0__1__6_chany_bottom_out[5] ,
    \cby_0__1__6_chany_bottom_out[6] ,
    \cby_0__1__6_chany_bottom_out[7] ,
    \cby_0__1__6_chany_bottom_out[8] ,
    \cby_0__1__6_chany_bottom_out[9] ,
    \cby_0__1__6_chany_bottom_out[10] ,
    \cby_0__1__6_chany_bottom_out[11] ,
    \cby_0__1__6_chany_bottom_out[12] ,
    \cby_0__1__6_chany_bottom_out[13] ,
    \cby_0__1__6_chany_bottom_out[14] ,
    \cby_0__1__6_chany_bottom_out[15] ,
    \cby_0__1__6_chany_bottom_out[16] ,
    \cby_0__1__6_chany_bottom_out[17] ,
    \cby_0__1__6_chany_bottom_out[18] ,
    \cby_0__1__6_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__1__5_chany_top_out[0] ,
    \sb_0__1__5_chany_top_out[1] ,
    \sb_0__1__5_chany_top_out[2] ,
    \sb_0__1__5_chany_top_out[3] ,
    \sb_0__1__5_chany_top_out[4] ,
    \sb_0__1__5_chany_top_out[5] ,
    \sb_0__1__5_chany_top_out[6] ,
    \sb_0__1__5_chany_top_out[7] ,
    \sb_0__1__5_chany_top_out[8] ,
    \sb_0__1__5_chany_top_out[9] ,
    \sb_0__1__5_chany_top_out[10] ,
    \sb_0__1__5_chany_top_out[11] ,
    \sb_0__1__5_chany_top_out[12] ,
    \sb_0__1__5_chany_top_out[13] ,
    \sb_0__1__5_chany_top_out[14] ,
    \sb_0__1__5_chany_top_out[15] ,
    \sb_0__1__5_chany_top_out[16] ,
    \sb_0__1__5_chany_top_out[17] ,
    \sb_0__1__5_chany_top_out[18] ,
    \sb_0__1__5_chany_top_out[19] }));
 sb_0__1_ sb_0__7_ (.bottom_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_upper),
    .ccff_head(cbx_1__1__6_ccff_tail),
    .ccff_tail(sb_0__1__6_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[35] ),
    .right_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__1__6_chanx_left_out[0] ,
    \cbx_1__1__6_chanx_left_out[1] ,
    \cbx_1__1__6_chanx_left_out[2] ,
    \cbx_1__1__6_chanx_left_out[3] ,
    \cbx_1__1__6_chanx_left_out[4] ,
    \cbx_1__1__6_chanx_left_out[5] ,
    \cbx_1__1__6_chanx_left_out[6] ,
    \cbx_1__1__6_chanx_left_out[7] ,
    \cbx_1__1__6_chanx_left_out[8] ,
    \cbx_1__1__6_chanx_left_out[9] ,
    \cbx_1__1__6_chanx_left_out[10] ,
    \cbx_1__1__6_chanx_left_out[11] ,
    \cbx_1__1__6_chanx_left_out[12] ,
    \cbx_1__1__6_chanx_left_out[13] ,
    \cbx_1__1__6_chanx_left_out[14] ,
    \cbx_1__1__6_chanx_left_out[15] ,
    \cbx_1__1__6_chanx_left_out[16] ,
    \cbx_1__1__6_chanx_left_out[17] ,
    \cbx_1__1__6_chanx_left_out[18] ,
    \cbx_1__1__6_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__1__6_chanx_right_out[0] ,
    \sb_0__1__6_chanx_right_out[1] ,
    \sb_0__1__6_chanx_right_out[2] ,
    \sb_0__1__6_chanx_right_out[3] ,
    \sb_0__1__6_chanx_right_out[4] ,
    \sb_0__1__6_chanx_right_out[5] ,
    \sb_0__1__6_chanx_right_out[6] ,
    \sb_0__1__6_chanx_right_out[7] ,
    \sb_0__1__6_chanx_right_out[8] ,
    \sb_0__1__6_chanx_right_out[9] ,
    \sb_0__1__6_chanx_right_out[10] ,
    \sb_0__1__6_chanx_right_out[11] ,
    \sb_0__1__6_chanx_right_out[12] ,
    \sb_0__1__6_chanx_right_out[13] ,
    \sb_0__1__6_chanx_right_out[14] ,
    \sb_0__1__6_chanx_right_out[15] ,
    \sb_0__1__6_chanx_right_out[16] ,
    \sb_0__1__6_chanx_right_out[17] ,
    \sb_0__1__6_chanx_right_out[18] ,
    \sb_0__1__6_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__6_chany_top_out[0] ,
    \cby_0__1__6_chany_top_out[1] ,
    \cby_0__1__6_chany_top_out[2] ,
    \cby_0__1__6_chany_top_out[3] ,
    \cby_0__1__6_chany_top_out[4] ,
    \cby_0__1__6_chany_top_out[5] ,
    \cby_0__1__6_chany_top_out[6] ,
    \cby_0__1__6_chany_top_out[7] ,
    \cby_0__1__6_chany_top_out[8] ,
    \cby_0__1__6_chany_top_out[9] ,
    \cby_0__1__6_chany_top_out[10] ,
    \cby_0__1__6_chany_top_out[11] ,
    \cby_0__1__6_chany_top_out[12] ,
    \cby_0__1__6_chany_top_out[13] ,
    \cby_0__1__6_chany_top_out[14] ,
    \cby_0__1__6_chany_top_out[15] ,
    \cby_0__1__6_chany_top_out[16] ,
    \cby_0__1__6_chany_top_out[17] ,
    \cby_0__1__6_chany_top_out[18] ,
    \cby_0__1__6_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__1__6_chany_bottom_out[0] ,
    \sb_0__1__6_chany_bottom_out[1] ,
    \sb_0__1__6_chany_bottom_out[2] ,
    \sb_0__1__6_chany_bottom_out[3] ,
    \sb_0__1__6_chany_bottom_out[4] ,
    \sb_0__1__6_chany_bottom_out[5] ,
    \sb_0__1__6_chany_bottom_out[6] ,
    \sb_0__1__6_chany_bottom_out[7] ,
    \sb_0__1__6_chany_bottom_out[8] ,
    \sb_0__1__6_chany_bottom_out[9] ,
    \sb_0__1__6_chany_bottom_out[10] ,
    \sb_0__1__6_chany_bottom_out[11] ,
    \sb_0__1__6_chany_bottom_out[12] ,
    \sb_0__1__6_chany_bottom_out[13] ,
    \sb_0__1__6_chany_bottom_out[14] ,
    \sb_0__1__6_chany_bottom_out[15] ,
    \sb_0__1__6_chany_bottom_out[16] ,
    \sb_0__1__6_chany_bottom_out[17] ,
    \sb_0__1__6_chany_bottom_out[18] ,
    \sb_0__1__6_chany_bottom_out[19] }),
    .chany_top_in({\cby_0__1__7_chany_bottom_out[0] ,
    \cby_0__1__7_chany_bottom_out[1] ,
    \cby_0__1__7_chany_bottom_out[2] ,
    \cby_0__1__7_chany_bottom_out[3] ,
    \cby_0__1__7_chany_bottom_out[4] ,
    \cby_0__1__7_chany_bottom_out[5] ,
    \cby_0__1__7_chany_bottom_out[6] ,
    \cby_0__1__7_chany_bottom_out[7] ,
    \cby_0__1__7_chany_bottom_out[8] ,
    \cby_0__1__7_chany_bottom_out[9] ,
    \cby_0__1__7_chany_bottom_out[10] ,
    \cby_0__1__7_chany_bottom_out[11] ,
    \cby_0__1__7_chany_bottom_out[12] ,
    \cby_0__1__7_chany_bottom_out[13] ,
    \cby_0__1__7_chany_bottom_out[14] ,
    \cby_0__1__7_chany_bottom_out[15] ,
    \cby_0__1__7_chany_bottom_out[16] ,
    \cby_0__1__7_chany_bottom_out[17] ,
    \cby_0__1__7_chany_bottom_out[18] ,
    \cby_0__1__7_chany_bottom_out[19] }),
    .chany_top_out({\sb_0__1__6_chany_top_out[0] ,
    \sb_0__1__6_chany_top_out[1] ,
    \sb_0__1__6_chany_top_out[2] ,
    \sb_0__1__6_chany_top_out[3] ,
    \sb_0__1__6_chany_top_out[4] ,
    \sb_0__1__6_chany_top_out[5] ,
    \sb_0__1__6_chany_top_out[6] ,
    \sb_0__1__6_chany_top_out[7] ,
    \sb_0__1__6_chany_top_out[8] ,
    \sb_0__1__6_chany_top_out[9] ,
    \sb_0__1__6_chany_top_out[10] ,
    \sb_0__1__6_chany_top_out[11] ,
    \sb_0__1__6_chany_top_out[12] ,
    \sb_0__1__6_chany_top_out[13] ,
    \sb_0__1__6_chany_top_out[14] ,
    \sb_0__1__6_chany_top_out[15] ,
    \sb_0__1__6_chany_top_out[16] ,
    \sb_0__1__6_chany_top_out[17] ,
    \sb_0__1__6_chany_top_out[18] ,
    \sb_0__1__6_chany_top_out[19] }));
 sb_0__2_ sb_0__8_ (.SC_IN_TOP(sc_head),
    .SC_OUT_BOT(\scff_Wires[0] ),
    .bottom_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_top_0_ccff_tail),
    .ccff_tail(sb_0__8__0_ccff_tail),
    .prog_clk_0_E_in(\prog_clk_0_wires[42] ),
    .right_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_right_in({\cbx_1__8__0_chanx_left_out[0] ,
    \cbx_1__8__0_chanx_left_out[1] ,
    \cbx_1__8__0_chanx_left_out[2] ,
    \cbx_1__8__0_chanx_left_out[3] ,
    \cbx_1__8__0_chanx_left_out[4] ,
    \cbx_1__8__0_chanx_left_out[5] ,
    \cbx_1__8__0_chanx_left_out[6] ,
    \cbx_1__8__0_chanx_left_out[7] ,
    \cbx_1__8__0_chanx_left_out[8] ,
    \cbx_1__8__0_chanx_left_out[9] ,
    \cbx_1__8__0_chanx_left_out[10] ,
    \cbx_1__8__0_chanx_left_out[11] ,
    \cbx_1__8__0_chanx_left_out[12] ,
    \cbx_1__8__0_chanx_left_out[13] ,
    \cbx_1__8__0_chanx_left_out[14] ,
    \cbx_1__8__0_chanx_left_out[15] ,
    \cbx_1__8__0_chanx_left_out[16] ,
    \cbx_1__8__0_chanx_left_out[17] ,
    \cbx_1__8__0_chanx_left_out[18] ,
    \cbx_1__8__0_chanx_left_out[19] }),
    .chanx_right_out({\sb_0__8__0_chanx_right_out[0] ,
    \sb_0__8__0_chanx_right_out[1] ,
    \sb_0__8__0_chanx_right_out[2] ,
    \sb_0__8__0_chanx_right_out[3] ,
    \sb_0__8__0_chanx_right_out[4] ,
    \sb_0__8__0_chanx_right_out[5] ,
    \sb_0__8__0_chanx_right_out[6] ,
    \sb_0__8__0_chanx_right_out[7] ,
    \sb_0__8__0_chanx_right_out[8] ,
    \sb_0__8__0_chanx_right_out[9] ,
    \sb_0__8__0_chanx_right_out[10] ,
    \sb_0__8__0_chanx_right_out[11] ,
    \sb_0__8__0_chanx_right_out[12] ,
    \sb_0__8__0_chanx_right_out[13] ,
    \sb_0__8__0_chanx_right_out[14] ,
    \sb_0__8__0_chanx_right_out[15] ,
    \sb_0__8__0_chanx_right_out[16] ,
    \sb_0__8__0_chanx_right_out[17] ,
    \sb_0__8__0_chanx_right_out[18] ,
    \sb_0__8__0_chanx_right_out[19] }),
    .chany_bottom_in({\cby_0__1__7_chany_top_out[0] ,
    \cby_0__1__7_chany_top_out[1] ,
    \cby_0__1__7_chany_top_out[2] ,
    \cby_0__1__7_chany_top_out[3] ,
    \cby_0__1__7_chany_top_out[4] ,
    \cby_0__1__7_chany_top_out[5] ,
    \cby_0__1__7_chany_top_out[6] ,
    \cby_0__1__7_chany_top_out[7] ,
    \cby_0__1__7_chany_top_out[8] ,
    \cby_0__1__7_chany_top_out[9] ,
    \cby_0__1__7_chany_top_out[10] ,
    \cby_0__1__7_chany_top_out[11] ,
    \cby_0__1__7_chany_top_out[12] ,
    \cby_0__1__7_chany_top_out[13] ,
    \cby_0__1__7_chany_top_out[14] ,
    \cby_0__1__7_chany_top_out[15] ,
    \cby_0__1__7_chany_top_out[16] ,
    \cby_0__1__7_chany_top_out[17] ,
    \cby_0__1__7_chany_top_out[18] ,
    \cby_0__1__7_chany_top_out[19] }),
    .chany_bottom_out({\sb_0__8__0_chany_bottom_out[0] ,
    \sb_0__8__0_chany_bottom_out[1] ,
    \sb_0__8__0_chany_bottom_out[2] ,
    \sb_0__8__0_chany_bottom_out[3] ,
    \sb_0__8__0_chany_bottom_out[4] ,
    \sb_0__8__0_chany_bottom_out[5] ,
    \sb_0__8__0_chany_bottom_out[6] ,
    \sb_0__8__0_chany_bottom_out[7] ,
    \sb_0__8__0_chany_bottom_out[8] ,
    \sb_0__8__0_chany_bottom_out[9] ,
    \sb_0__8__0_chany_bottom_out[10] ,
    \sb_0__8__0_chany_bottom_out[11] ,
    \sb_0__8__0_chany_bottom_out[12] ,
    \sb_0__8__0_chany_bottom_out[13] ,
    \sb_0__8__0_chany_bottom_out[14] ,
    \sb_0__8__0_chany_bottom_out[15] ,
    \sb_0__8__0_chany_bottom_out[16] ,
    \sb_0__8__0_chany_bottom_out[17] ,
    \sb_0__8__0_chany_bottom_out[18] ,
    \sb_0__8__0_chany_bottom_out[19] }));
 sb_1__0_ sb_1__0_ (.SC_IN_TOP(\scff_Wires[18] ),
    .SC_OUT_TOP(\scff_Wires[19] ),
    .ccff_head(grid_io_bottom_6_ccff_tail),
    .ccff_tail(sb_1__0__0_ccff_tail),
    .left_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[2] ),
    .right_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__0_chanx_right_out[0] ,
    \cbx_1__0__0_chanx_right_out[1] ,
    \cbx_1__0__0_chanx_right_out[2] ,
    \cbx_1__0__0_chanx_right_out[3] ,
    \cbx_1__0__0_chanx_right_out[4] ,
    \cbx_1__0__0_chanx_right_out[5] ,
    \cbx_1__0__0_chanx_right_out[6] ,
    \cbx_1__0__0_chanx_right_out[7] ,
    \cbx_1__0__0_chanx_right_out[8] ,
    \cbx_1__0__0_chanx_right_out[9] ,
    \cbx_1__0__0_chanx_right_out[10] ,
    \cbx_1__0__0_chanx_right_out[11] ,
    \cbx_1__0__0_chanx_right_out[12] ,
    \cbx_1__0__0_chanx_right_out[13] ,
    \cbx_1__0__0_chanx_right_out[14] ,
    \cbx_1__0__0_chanx_right_out[15] ,
    \cbx_1__0__0_chanx_right_out[16] ,
    \cbx_1__0__0_chanx_right_out[17] ,
    \cbx_1__0__0_chanx_right_out[18] ,
    \cbx_1__0__0_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__0__0_chanx_left_out[0] ,
    \sb_1__0__0_chanx_left_out[1] ,
    \sb_1__0__0_chanx_left_out[2] ,
    \sb_1__0__0_chanx_left_out[3] ,
    \sb_1__0__0_chanx_left_out[4] ,
    \sb_1__0__0_chanx_left_out[5] ,
    \sb_1__0__0_chanx_left_out[6] ,
    \sb_1__0__0_chanx_left_out[7] ,
    \sb_1__0__0_chanx_left_out[8] ,
    \sb_1__0__0_chanx_left_out[9] ,
    \sb_1__0__0_chanx_left_out[10] ,
    \sb_1__0__0_chanx_left_out[11] ,
    \sb_1__0__0_chanx_left_out[12] ,
    \sb_1__0__0_chanx_left_out[13] ,
    \sb_1__0__0_chanx_left_out[14] ,
    \sb_1__0__0_chanx_left_out[15] ,
    \sb_1__0__0_chanx_left_out[16] ,
    \sb_1__0__0_chanx_left_out[17] ,
    \sb_1__0__0_chanx_left_out[18] ,
    \sb_1__0__0_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__0__1_chanx_left_out[0] ,
    \cbx_1__0__1_chanx_left_out[1] ,
    \cbx_1__0__1_chanx_left_out[2] ,
    \cbx_1__0__1_chanx_left_out[3] ,
    \cbx_1__0__1_chanx_left_out[4] ,
    \cbx_1__0__1_chanx_left_out[5] ,
    \cbx_1__0__1_chanx_left_out[6] ,
    \cbx_1__0__1_chanx_left_out[7] ,
    \cbx_1__0__1_chanx_left_out[8] ,
    \cbx_1__0__1_chanx_left_out[9] ,
    \cbx_1__0__1_chanx_left_out[10] ,
    \cbx_1__0__1_chanx_left_out[11] ,
    \cbx_1__0__1_chanx_left_out[12] ,
    \cbx_1__0__1_chanx_left_out[13] ,
    \cbx_1__0__1_chanx_left_out[14] ,
    \cbx_1__0__1_chanx_left_out[15] ,
    \cbx_1__0__1_chanx_left_out[16] ,
    \cbx_1__0__1_chanx_left_out[17] ,
    \cbx_1__0__1_chanx_left_out[18] ,
    \cbx_1__0__1_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__0__0_chanx_right_out[0] ,
    \sb_1__0__0_chanx_right_out[1] ,
    \sb_1__0__0_chanx_right_out[2] ,
    \sb_1__0__0_chanx_right_out[3] ,
    \sb_1__0__0_chanx_right_out[4] ,
    \sb_1__0__0_chanx_right_out[5] ,
    \sb_1__0__0_chanx_right_out[6] ,
    \sb_1__0__0_chanx_right_out[7] ,
    \sb_1__0__0_chanx_right_out[8] ,
    \sb_1__0__0_chanx_right_out[9] ,
    \sb_1__0__0_chanx_right_out[10] ,
    \sb_1__0__0_chanx_right_out[11] ,
    \sb_1__0__0_chanx_right_out[12] ,
    \sb_1__0__0_chanx_right_out[13] ,
    \sb_1__0__0_chanx_right_out[14] ,
    \sb_1__0__0_chanx_right_out[15] ,
    \sb_1__0__0_chanx_right_out[16] ,
    \sb_1__0__0_chanx_right_out[17] ,
    \sb_1__0__0_chanx_right_out[18] ,
    \sb_1__0__0_chanx_right_out[19] }),
    .chany_top_in({\cby_1__1__0_chany_bottom_out[0] ,
    \cby_1__1__0_chany_bottom_out[1] ,
    \cby_1__1__0_chany_bottom_out[2] ,
    \cby_1__1__0_chany_bottom_out[3] ,
    \cby_1__1__0_chany_bottom_out[4] ,
    \cby_1__1__0_chany_bottom_out[5] ,
    \cby_1__1__0_chany_bottom_out[6] ,
    \cby_1__1__0_chany_bottom_out[7] ,
    \cby_1__1__0_chany_bottom_out[8] ,
    \cby_1__1__0_chany_bottom_out[9] ,
    \cby_1__1__0_chany_bottom_out[10] ,
    \cby_1__1__0_chany_bottom_out[11] ,
    \cby_1__1__0_chany_bottom_out[12] ,
    \cby_1__1__0_chany_bottom_out[13] ,
    \cby_1__1__0_chany_bottom_out[14] ,
    \cby_1__1__0_chany_bottom_out[15] ,
    \cby_1__1__0_chany_bottom_out[16] ,
    \cby_1__1__0_chany_bottom_out[17] ,
    \cby_1__1__0_chany_bottom_out[18] ,
    \cby_1__1__0_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__0__0_chany_top_out[0] ,
    \sb_1__0__0_chany_top_out[1] ,
    \sb_1__0__0_chany_top_out[2] ,
    \sb_1__0__0_chany_top_out[3] ,
    \sb_1__0__0_chany_top_out[4] ,
    \sb_1__0__0_chany_top_out[5] ,
    \sb_1__0__0_chany_top_out[6] ,
    \sb_1__0__0_chany_top_out[7] ,
    \sb_1__0__0_chany_top_out[8] ,
    \sb_1__0__0_chany_top_out[9] ,
    \sb_1__0__0_chany_top_out[10] ,
    \sb_1__0__0_chany_top_out[11] ,
    \sb_1__0__0_chany_top_out[12] ,
    \sb_1__0__0_chany_top_out[13] ,
    \sb_1__0__0_chany_top_out[14] ,
    \sb_1__0__0_chany_top_out[15] ,
    \sb_1__0__0_chany_top_out[16] ,
    \sb_1__0__0_chany_top_out[17] ,
    \sb_1__0__0_chany_top_out[18] ,
    \sb_1__0__0_chany_top_out[19] }));
 sb_1__1_ sb_1__1_ (.bottom_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__7_ccff_tail),
    .ccff_tail(sb_1__1__0_ccff_tail),
    .clk_1_E_out(\clk_1_wires[1] ),
    .clk_1_N_in(\clk_2_wires[8] ),
    .clk_1_W_out(\clk_1_wires[2] ),
    .left_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[8] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[1] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[8] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[2] ),
    .right_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__0_chanx_right_out[0] ,
    \cbx_1__1__0_chanx_right_out[1] ,
    \cbx_1__1__0_chanx_right_out[2] ,
    \cbx_1__1__0_chanx_right_out[3] ,
    \cbx_1__1__0_chanx_right_out[4] ,
    \cbx_1__1__0_chanx_right_out[5] ,
    \cbx_1__1__0_chanx_right_out[6] ,
    \cbx_1__1__0_chanx_right_out[7] ,
    \cbx_1__1__0_chanx_right_out[8] ,
    \cbx_1__1__0_chanx_right_out[9] ,
    \cbx_1__1__0_chanx_right_out[10] ,
    \cbx_1__1__0_chanx_right_out[11] ,
    \cbx_1__1__0_chanx_right_out[12] ,
    \cbx_1__1__0_chanx_right_out[13] ,
    \cbx_1__1__0_chanx_right_out[14] ,
    \cbx_1__1__0_chanx_right_out[15] ,
    \cbx_1__1__0_chanx_right_out[16] ,
    \cbx_1__1__0_chanx_right_out[17] ,
    \cbx_1__1__0_chanx_right_out[18] ,
    \cbx_1__1__0_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__0_chanx_left_out[0] ,
    \sb_1__1__0_chanx_left_out[1] ,
    \sb_1__1__0_chanx_left_out[2] ,
    \sb_1__1__0_chanx_left_out[3] ,
    \sb_1__1__0_chanx_left_out[4] ,
    \sb_1__1__0_chanx_left_out[5] ,
    \sb_1__1__0_chanx_left_out[6] ,
    \sb_1__1__0_chanx_left_out[7] ,
    \sb_1__1__0_chanx_left_out[8] ,
    \sb_1__1__0_chanx_left_out[9] ,
    \sb_1__1__0_chanx_left_out[10] ,
    \sb_1__1__0_chanx_left_out[11] ,
    \sb_1__1__0_chanx_left_out[12] ,
    \sb_1__1__0_chanx_left_out[13] ,
    \sb_1__1__0_chanx_left_out[14] ,
    \sb_1__1__0_chanx_left_out[15] ,
    \sb_1__1__0_chanx_left_out[16] ,
    \sb_1__1__0_chanx_left_out[17] ,
    \sb_1__1__0_chanx_left_out[18] ,
    \sb_1__1__0_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__7_chanx_left_out[0] ,
    \cbx_1__1__7_chanx_left_out[1] ,
    \cbx_1__1__7_chanx_left_out[2] ,
    \cbx_1__1__7_chanx_left_out[3] ,
    \cbx_1__1__7_chanx_left_out[4] ,
    \cbx_1__1__7_chanx_left_out[5] ,
    \cbx_1__1__7_chanx_left_out[6] ,
    \cbx_1__1__7_chanx_left_out[7] ,
    \cbx_1__1__7_chanx_left_out[8] ,
    \cbx_1__1__7_chanx_left_out[9] ,
    \cbx_1__1__7_chanx_left_out[10] ,
    \cbx_1__1__7_chanx_left_out[11] ,
    \cbx_1__1__7_chanx_left_out[12] ,
    \cbx_1__1__7_chanx_left_out[13] ,
    \cbx_1__1__7_chanx_left_out[14] ,
    \cbx_1__1__7_chanx_left_out[15] ,
    \cbx_1__1__7_chanx_left_out[16] ,
    \cbx_1__1__7_chanx_left_out[17] ,
    \cbx_1__1__7_chanx_left_out[18] ,
    \cbx_1__1__7_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__0_chanx_right_out[0] ,
    \sb_1__1__0_chanx_right_out[1] ,
    \sb_1__1__0_chanx_right_out[2] ,
    \sb_1__1__0_chanx_right_out[3] ,
    \sb_1__1__0_chanx_right_out[4] ,
    \sb_1__1__0_chanx_right_out[5] ,
    \sb_1__1__0_chanx_right_out[6] ,
    \sb_1__1__0_chanx_right_out[7] ,
    \sb_1__1__0_chanx_right_out[8] ,
    \sb_1__1__0_chanx_right_out[9] ,
    \sb_1__1__0_chanx_right_out[10] ,
    \sb_1__1__0_chanx_right_out[11] ,
    \sb_1__1__0_chanx_right_out[12] ,
    \sb_1__1__0_chanx_right_out[13] ,
    \sb_1__1__0_chanx_right_out[14] ,
    \sb_1__1__0_chanx_right_out[15] ,
    \sb_1__1__0_chanx_right_out[16] ,
    \sb_1__1__0_chanx_right_out[17] ,
    \sb_1__1__0_chanx_right_out[18] ,
    \sb_1__1__0_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__0_chany_top_out[0] ,
    \cby_1__1__0_chany_top_out[1] ,
    \cby_1__1__0_chany_top_out[2] ,
    \cby_1__1__0_chany_top_out[3] ,
    \cby_1__1__0_chany_top_out[4] ,
    \cby_1__1__0_chany_top_out[5] ,
    \cby_1__1__0_chany_top_out[6] ,
    \cby_1__1__0_chany_top_out[7] ,
    \cby_1__1__0_chany_top_out[8] ,
    \cby_1__1__0_chany_top_out[9] ,
    \cby_1__1__0_chany_top_out[10] ,
    \cby_1__1__0_chany_top_out[11] ,
    \cby_1__1__0_chany_top_out[12] ,
    \cby_1__1__0_chany_top_out[13] ,
    \cby_1__1__0_chany_top_out[14] ,
    \cby_1__1__0_chany_top_out[15] ,
    \cby_1__1__0_chany_top_out[16] ,
    \cby_1__1__0_chany_top_out[17] ,
    \cby_1__1__0_chany_top_out[18] ,
    \cby_1__1__0_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__0_chany_bottom_out[0] ,
    \sb_1__1__0_chany_bottom_out[1] ,
    \sb_1__1__0_chany_bottom_out[2] ,
    \sb_1__1__0_chany_bottom_out[3] ,
    \sb_1__1__0_chany_bottom_out[4] ,
    \sb_1__1__0_chany_bottom_out[5] ,
    \sb_1__1__0_chany_bottom_out[6] ,
    \sb_1__1__0_chany_bottom_out[7] ,
    \sb_1__1__0_chany_bottom_out[8] ,
    \sb_1__1__0_chany_bottom_out[9] ,
    \sb_1__1__0_chany_bottom_out[10] ,
    \sb_1__1__0_chany_bottom_out[11] ,
    \sb_1__1__0_chany_bottom_out[12] ,
    \sb_1__1__0_chany_bottom_out[13] ,
    \sb_1__1__0_chany_bottom_out[14] ,
    \sb_1__1__0_chany_bottom_out[15] ,
    \sb_1__1__0_chany_bottom_out[16] ,
    \sb_1__1__0_chany_bottom_out[17] ,
    \sb_1__1__0_chany_bottom_out[18] ,
    \sb_1__1__0_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__1_chany_bottom_out[0] ,
    \cby_1__1__1_chany_bottom_out[1] ,
    \cby_1__1__1_chany_bottom_out[2] ,
    \cby_1__1__1_chany_bottom_out[3] ,
    \cby_1__1__1_chany_bottom_out[4] ,
    \cby_1__1__1_chany_bottom_out[5] ,
    \cby_1__1__1_chany_bottom_out[6] ,
    \cby_1__1__1_chany_bottom_out[7] ,
    \cby_1__1__1_chany_bottom_out[8] ,
    \cby_1__1__1_chany_bottom_out[9] ,
    \cby_1__1__1_chany_bottom_out[10] ,
    \cby_1__1__1_chany_bottom_out[11] ,
    \cby_1__1__1_chany_bottom_out[12] ,
    \cby_1__1__1_chany_bottom_out[13] ,
    \cby_1__1__1_chany_bottom_out[14] ,
    \cby_1__1__1_chany_bottom_out[15] ,
    \cby_1__1__1_chany_bottom_out[16] ,
    \cby_1__1__1_chany_bottom_out[17] ,
    \cby_1__1__1_chany_bottom_out[18] ,
    \cby_1__1__1_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__0_chany_top_out[0] ,
    \sb_1__1__0_chany_top_out[1] ,
    \sb_1__1__0_chany_top_out[2] ,
    \sb_1__1__0_chany_top_out[3] ,
    \sb_1__1__0_chany_top_out[4] ,
    \sb_1__1__0_chany_top_out[5] ,
    \sb_1__1__0_chany_top_out[6] ,
    \sb_1__1__0_chany_top_out[7] ,
    \sb_1__1__0_chany_top_out[8] ,
    \sb_1__1__0_chany_top_out[9] ,
    \sb_1__1__0_chany_top_out[10] ,
    \sb_1__1__0_chany_top_out[11] ,
    \sb_1__1__0_chany_top_out[12] ,
    \sb_1__1__0_chany_top_out[13] ,
    \sb_1__1__0_chany_top_out[14] ,
    \sb_1__1__0_chany_top_out[15] ,
    \sb_1__1__0_chany_top_out[16] ,
    \sb_1__1__0_chany_top_out[17] ,
    \sb_1__1__0_chany_top_out[18] ,
    \sb_1__1__0_chany_top_out[19] }));
 sb_1__1_ sb_1__2_ (.bottom_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__8_ccff_tail),
    .ccff_tail(sb_1__1__1_ccff_tail),
    .clk_2_N_in(\clk_2_wires[4] ),
    .clk_2_N_out(\clk_2_wires[5] ),
    .clk_2_S_out(\clk_2_wires[7] ),
    .left_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[13] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[4] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[5] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[7] ),
    .right_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__1_chanx_right_out[0] ,
    \cbx_1__1__1_chanx_right_out[1] ,
    \cbx_1__1__1_chanx_right_out[2] ,
    \cbx_1__1__1_chanx_right_out[3] ,
    \cbx_1__1__1_chanx_right_out[4] ,
    \cbx_1__1__1_chanx_right_out[5] ,
    \cbx_1__1__1_chanx_right_out[6] ,
    \cbx_1__1__1_chanx_right_out[7] ,
    \cbx_1__1__1_chanx_right_out[8] ,
    \cbx_1__1__1_chanx_right_out[9] ,
    \cbx_1__1__1_chanx_right_out[10] ,
    \cbx_1__1__1_chanx_right_out[11] ,
    \cbx_1__1__1_chanx_right_out[12] ,
    \cbx_1__1__1_chanx_right_out[13] ,
    \cbx_1__1__1_chanx_right_out[14] ,
    \cbx_1__1__1_chanx_right_out[15] ,
    \cbx_1__1__1_chanx_right_out[16] ,
    \cbx_1__1__1_chanx_right_out[17] ,
    \cbx_1__1__1_chanx_right_out[18] ,
    \cbx_1__1__1_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__1_chanx_left_out[0] ,
    \sb_1__1__1_chanx_left_out[1] ,
    \sb_1__1__1_chanx_left_out[2] ,
    \sb_1__1__1_chanx_left_out[3] ,
    \sb_1__1__1_chanx_left_out[4] ,
    \sb_1__1__1_chanx_left_out[5] ,
    \sb_1__1__1_chanx_left_out[6] ,
    \sb_1__1__1_chanx_left_out[7] ,
    \sb_1__1__1_chanx_left_out[8] ,
    \sb_1__1__1_chanx_left_out[9] ,
    \sb_1__1__1_chanx_left_out[10] ,
    \sb_1__1__1_chanx_left_out[11] ,
    \sb_1__1__1_chanx_left_out[12] ,
    \sb_1__1__1_chanx_left_out[13] ,
    \sb_1__1__1_chanx_left_out[14] ,
    \sb_1__1__1_chanx_left_out[15] ,
    \sb_1__1__1_chanx_left_out[16] ,
    \sb_1__1__1_chanx_left_out[17] ,
    \sb_1__1__1_chanx_left_out[18] ,
    \sb_1__1__1_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__8_chanx_left_out[0] ,
    \cbx_1__1__8_chanx_left_out[1] ,
    \cbx_1__1__8_chanx_left_out[2] ,
    \cbx_1__1__8_chanx_left_out[3] ,
    \cbx_1__1__8_chanx_left_out[4] ,
    \cbx_1__1__8_chanx_left_out[5] ,
    \cbx_1__1__8_chanx_left_out[6] ,
    \cbx_1__1__8_chanx_left_out[7] ,
    \cbx_1__1__8_chanx_left_out[8] ,
    \cbx_1__1__8_chanx_left_out[9] ,
    \cbx_1__1__8_chanx_left_out[10] ,
    \cbx_1__1__8_chanx_left_out[11] ,
    \cbx_1__1__8_chanx_left_out[12] ,
    \cbx_1__1__8_chanx_left_out[13] ,
    \cbx_1__1__8_chanx_left_out[14] ,
    \cbx_1__1__8_chanx_left_out[15] ,
    \cbx_1__1__8_chanx_left_out[16] ,
    \cbx_1__1__8_chanx_left_out[17] ,
    \cbx_1__1__8_chanx_left_out[18] ,
    \cbx_1__1__8_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__1_chanx_right_out[0] ,
    \sb_1__1__1_chanx_right_out[1] ,
    \sb_1__1__1_chanx_right_out[2] ,
    \sb_1__1__1_chanx_right_out[3] ,
    \sb_1__1__1_chanx_right_out[4] ,
    \sb_1__1__1_chanx_right_out[5] ,
    \sb_1__1__1_chanx_right_out[6] ,
    \sb_1__1__1_chanx_right_out[7] ,
    \sb_1__1__1_chanx_right_out[8] ,
    \sb_1__1__1_chanx_right_out[9] ,
    \sb_1__1__1_chanx_right_out[10] ,
    \sb_1__1__1_chanx_right_out[11] ,
    \sb_1__1__1_chanx_right_out[12] ,
    \sb_1__1__1_chanx_right_out[13] ,
    \sb_1__1__1_chanx_right_out[14] ,
    \sb_1__1__1_chanx_right_out[15] ,
    \sb_1__1__1_chanx_right_out[16] ,
    \sb_1__1__1_chanx_right_out[17] ,
    \sb_1__1__1_chanx_right_out[18] ,
    \sb_1__1__1_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__1_chany_top_out[0] ,
    \cby_1__1__1_chany_top_out[1] ,
    \cby_1__1__1_chany_top_out[2] ,
    \cby_1__1__1_chany_top_out[3] ,
    \cby_1__1__1_chany_top_out[4] ,
    \cby_1__1__1_chany_top_out[5] ,
    \cby_1__1__1_chany_top_out[6] ,
    \cby_1__1__1_chany_top_out[7] ,
    \cby_1__1__1_chany_top_out[8] ,
    \cby_1__1__1_chany_top_out[9] ,
    \cby_1__1__1_chany_top_out[10] ,
    \cby_1__1__1_chany_top_out[11] ,
    \cby_1__1__1_chany_top_out[12] ,
    \cby_1__1__1_chany_top_out[13] ,
    \cby_1__1__1_chany_top_out[14] ,
    \cby_1__1__1_chany_top_out[15] ,
    \cby_1__1__1_chany_top_out[16] ,
    \cby_1__1__1_chany_top_out[17] ,
    \cby_1__1__1_chany_top_out[18] ,
    \cby_1__1__1_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__1_chany_bottom_out[0] ,
    \sb_1__1__1_chany_bottom_out[1] ,
    \sb_1__1__1_chany_bottom_out[2] ,
    \sb_1__1__1_chany_bottom_out[3] ,
    \sb_1__1__1_chany_bottom_out[4] ,
    \sb_1__1__1_chany_bottom_out[5] ,
    \sb_1__1__1_chany_bottom_out[6] ,
    \sb_1__1__1_chany_bottom_out[7] ,
    \sb_1__1__1_chany_bottom_out[8] ,
    \sb_1__1__1_chany_bottom_out[9] ,
    \sb_1__1__1_chany_bottom_out[10] ,
    \sb_1__1__1_chany_bottom_out[11] ,
    \sb_1__1__1_chany_bottom_out[12] ,
    \sb_1__1__1_chany_bottom_out[13] ,
    \sb_1__1__1_chany_bottom_out[14] ,
    \sb_1__1__1_chany_bottom_out[15] ,
    \sb_1__1__1_chany_bottom_out[16] ,
    \sb_1__1__1_chany_bottom_out[17] ,
    \sb_1__1__1_chany_bottom_out[18] ,
    \sb_1__1__1_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__2_chany_bottom_out[0] ,
    \cby_1__1__2_chany_bottom_out[1] ,
    \cby_1__1__2_chany_bottom_out[2] ,
    \cby_1__1__2_chany_bottom_out[3] ,
    \cby_1__1__2_chany_bottom_out[4] ,
    \cby_1__1__2_chany_bottom_out[5] ,
    \cby_1__1__2_chany_bottom_out[6] ,
    \cby_1__1__2_chany_bottom_out[7] ,
    \cby_1__1__2_chany_bottom_out[8] ,
    \cby_1__1__2_chany_bottom_out[9] ,
    \cby_1__1__2_chany_bottom_out[10] ,
    \cby_1__1__2_chany_bottom_out[11] ,
    \cby_1__1__2_chany_bottom_out[12] ,
    \cby_1__1__2_chany_bottom_out[13] ,
    \cby_1__1__2_chany_bottom_out[14] ,
    \cby_1__1__2_chany_bottom_out[15] ,
    \cby_1__1__2_chany_bottom_out[16] ,
    \cby_1__1__2_chany_bottom_out[17] ,
    \cby_1__1__2_chany_bottom_out[18] ,
    \cby_1__1__2_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__1_chany_top_out[0] ,
    \sb_1__1__1_chany_top_out[1] ,
    \sb_1__1__1_chany_top_out[2] ,
    \sb_1__1__1_chany_top_out[3] ,
    \sb_1__1__1_chany_top_out[4] ,
    \sb_1__1__1_chany_top_out[5] ,
    \sb_1__1__1_chany_top_out[6] ,
    \sb_1__1__1_chany_top_out[7] ,
    \sb_1__1__1_chany_top_out[8] ,
    \sb_1__1__1_chany_top_out[9] ,
    \sb_1__1__1_chany_top_out[10] ,
    \sb_1__1__1_chany_top_out[11] ,
    \sb_1__1__1_chany_top_out[12] ,
    \sb_1__1__1_chany_top_out[13] ,
    \sb_1__1__1_chany_top_out[14] ,
    \sb_1__1__1_chany_top_out[15] ,
    \sb_1__1__1_chany_top_out[16] ,
    \sb_1__1__1_chany_top_out[17] ,
    \sb_1__1__1_chany_top_out[18] ,
    \sb_1__1__1_chany_top_out[19] }));
 sb_1__1_ sb_1__3_ (.bottom_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__9_ccff_tail),
    .ccff_tail(sb_1__1__2_ccff_tail),
    .clk_1_E_out(\clk_1_wires[8] ),
    .clk_1_N_in(\clk_2_wires[6] ),
    .clk_1_W_out(\clk_1_wires[9] ),
    .left_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[18] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[8] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[6] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[9] ),
    .right_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__2_chanx_right_out[0] ,
    \cbx_1__1__2_chanx_right_out[1] ,
    \cbx_1__1__2_chanx_right_out[2] ,
    \cbx_1__1__2_chanx_right_out[3] ,
    \cbx_1__1__2_chanx_right_out[4] ,
    \cbx_1__1__2_chanx_right_out[5] ,
    \cbx_1__1__2_chanx_right_out[6] ,
    \cbx_1__1__2_chanx_right_out[7] ,
    \cbx_1__1__2_chanx_right_out[8] ,
    \cbx_1__1__2_chanx_right_out[9] ,
    \cbx_1__1__2_chanx_right_out[10] ,
    \cbx_1__1__2_chanx_right_out[11] ,
    \cbx_1__1__2_chanx_right_out[12] ,
    \cbx_1__1__2_chanx_right_out[13] ,
    \cbx_1__1__2_chanx_right_out[14] ,
    \cbx_1__1__2_chanx_right_out[15] ,
    \cbx_1__1__2_chanx_right_out[16] ,
    \cbx_1__1__2_chanx_right_out[17] ,
    \cbx_1__1__2_chanx_right_out[18] ,
    \cbx_1__1__2_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__2_chanx_left_out[0] ,
    \sb_1__1__2_chanx_left_out[1] ,
    \sb_1__1__2_chanx_left_out[2] ,
    \sb_1__1__2_chanx_left_out[3] ,
    \sb_1__1__2_chanx_left_out[4] ,
    \sb_1__1__2_chanx_left_out[5] ,
    \sb_1__1__2_chanx_left_out[6] ,
    \sb_1__1__2_chanx_left_out[7] ,
    \sb_1__1__2_chanx_left_out[8] ,
    \sb_1__1__2_chanx_left_out[9] ,
    \sb_1__1__2_chanx_left_out[10] ,
    \sb_1__1__2_chanx_left_out[11] ,
    \sb_1__1__2_chanx_left_out[12] ,
    \sb_1__1__2_chanx_left_out[13] ,
    \sb_1__1__2_chanx_left_out[14] ,
    \sb_1__1__2_chanx_left_out[15] ,
    \sb_1__1__2_chanx_left_out[16] ,
    \sb_1__1__2_chanx_left_out[17] ,
    \sb_1__1__2_chanx_left_out[18] ,
    \sb_1__1__2_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__9_chanx_left_out[0] ,
    \cbx_1__1__9_chanx_left_out[1] ,
    \cbx_1__1__9_chanx_left_out[2] ,
    \cbx_1__1__9_chanx_left_out[3] ,
    \cbx_1__1__9_chanx_left_out[4] ,
    \cbx_1__1__9_chanx_left_out[5] ,
    \cbx_1__1__9_chanx_left_out[6] ,
    \cbx_1__1__9_chanx_left_out[7] ,
    \cbx_1__1__9_chanx_left_out[8] ,
    \cbx_1__1__9_chanx_left_out[9] ,
    \cbx_1__1__9_chanx_left_out[10] ,
    \cbx_1__1__9_chanx_left_out[11] ,
    \cbx_1__1__9_chanx_left_out[12] ,
    \cbx_1__1__9_chanx_left_out[13] ,
    \cbx_1__1__9_chanx_left_out[14] ,
    \cbx_1__1__9_chanx_left_out[15] ,
    \cbx_1__1__9_chanx_left_out[16] ,
    \cbx_1__1__9_chanx_left_out[17] ,
    \cbx_1__1__9_chanx_left_out[18] ,
    \cbx_1__1__9_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__2_chanx_right_out[0] ,
    \sb_1__1__2_chanx_right_out[1] ,
    \sb_1__1__2_chanx_right_out[2] ,
    \sb_1__1__2_chanx_right_out[3] ,
    \sb_1__1__2_chanx_right_out[4] ,
    \sb_1__1__2_chanx_right_out[5] ,
    \sb_1__1__2_chanx_right_out[6] ,
    \sb_1__1__2_chanx_right_out[7] ,
    \sb_1__1__2_chanx_right_out[8] ,
    \sb_1__1__2_chanx_right_out[9] ,
    \sb_1__1__2_chanx_right_out[10] ,
    \sb_1__1__2_chanx_right_out[11] ,
    \sb_1__1__2_chanx_right_out[12] ,
    \sb_1__1__2_chanx_right_out[13] ,
    \sb_1__1__2_chanx_right_out[14] ,
    \sb_1__1__2_chanx_right_out[15] ,
    \sb_1__1__2_chanx_right_out[16] ,
    \sb_1__1__2_chanx_right_out[17] ,
    \sb_1__1__2_chanx_right_out[18] ,
    \sb_1__1__2_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__2_chany_top_out[0] ,
    \cby_1__1__2_chany_top_out[1] ,
    \cby_1__1__2_chany_top_out[2] ,
    \cby_1__1__2_chany_top_out[3] ,
    \cby_1__1__2_chany_top_out[4] ,
    \cby_1__1__2_chany_top_out[5] ,
    \cby_1__1__2_chany_top_out[6] ,
    \cby_1__1__2_chany_top_out[7] ,
    \cby_1__1__2_chany_top_out[8] ,
    \cby_1__1__2_chany_top_out[9] ,
    \cby_1__1__2_chany_top_out[10] ,
    \cby_1__1__2_chany_top_out[11] ,
    \cby_1__1__2_chany_top_out[12] ,
    \cby_1__1__2_chany_top_out[13] ,
    \cby_1__1__2_chany_top_out[14] ,
    \cby_1__1__2_chany_top_out[15] ,
    \cby_1__1__2_chany_top_out[16] ,
    \cby_1__1__2_chany_top_out[17] ,
    \cby_1__1__2_chany_top_out[18] ,
    \cby_1__1__2_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__2_chany_bottom_out[0] ,
    \sb_1__1__2_chany_bottom_out[1] ,
    \sb_1__1__2_chany_bottom_out[2] ,
    \sb_1__1__2_chany_bottom_out[3] ,
    \sb_1__1__2_chany_bottom_out[4] ,
    \sb_1__1__2_chany_bottom_out[5] ,
    \sb_1__1__2_chany_bottom_out[6] ,
    \sb_1__1__2_chany_bottom_out[7] ,
    \sb_1__1__2_chany_bottom_out[8] ,
    \sb_1__1__2_chany_bottom_out[9] ,
    \sb_1__1__2_chany_bottom_out[10] ,
    \sb_1__1__2_chany_bottom_out[11] ,
    \sb_1__1__2_chany_bottom_out[12] ,
    \sb_1__1__2_chany_bottom_out[13] ,
    \sb_1__1__2_chany_bottom_out[14] ,
    \sb_1__1__2_chany_bottom_out[15] ,
    \sb_1__1__2_chany_bottom_out[16] ,
    \sb_1__1__2_chany_bottom_out[17] ,
    \sb_1__1__2_chany_bottom_out[18] ,
    \sb_1__1__2_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__3_chany_bottom_out[0] ,
    \cby_1__1__3_chany_bottom_out[1] ,
    \cby_1__1__3_chany_bottom_out[2] ,
    \cby_1__1__3_chany_bottom_out[3] ,
    \cby_1__1__3_chany_bottom_out[4] ,
    \cby_1__1__3_chany_bottom_out[5] ,
    \cby_1__1__3_chany_bottom_out[6] ,
    \cby_1__1__3_chany_bottom_out[7] ,
    \cby_1__1__3_chany_bottom_out[8] ,
    \cby_1__1__3_chany_bottom_out[9] ,
    \cby_1__1__3_chany_bottom_out[10] ,
    \cby_1__1__3_chany_bottom_out[11] ,
    \cby_1__1__3_chany_bottom_out[12] ,
    \cby_1__1__3_chany_bottom_out[13] ,
    \cby_1__1__3_chany_bottom_out[14] ,
    \cby_1__1__3_chany_bottom_out[15] ,
    \cby_1__1__3_chany_bottom_out[16] ,
    \cby_1__1__3_chany_bottom_out[17] ,
    \cby_1__1__3_chany_bottom_out[18] ,
    \cby_1__1__3_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__2_chany_top_out[0] ,
    \sb_1__1__2_chany_top_out[1] ,
    \sb_1__1__2_chany_top_out[2] ,
    \sb_1__1__2_chany_top_out[3] ,
    \sb_1__1__2_chany_top_out[4] ,
    \sb_1__1__2_chany_top_out[5] ,
    \sb_1__1__2_chany_top_out[6] ,
    \sb_1__1__2_chany_top_out[7] ,
    \sb_1__1__2_chany_top_out[8] ,
    \sb_1__1__2_chany_top_out[9] ,
    \sb_1__1__2_chany_top_out[10] ,
    \sb_1__1__2_chany_top_out[11] ,
    \sb_1__1__2_chany_top_out[12] ,
    \sb_1__1__2_chany_top_out[13] ,
    \sb_1__1__2_chany_top_out[14] ,
    \sb_1__1__2_chany_top_out[15] ,
    \sb_1__1__2_chany_top_out[16] ,
    \sb_1__1__2_chany_top_out[17] ,
    \sb_1__1__2_chany_top_out[18] ,
    \sb_1__1__2_chany_top_out[19] }));
 sb_1__1_ sb_1__4_ (.bottom_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__10_ccff_tail),
    .ccff_tail(sb_1__1__3_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[23] ),
    .right_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__3_chanx_right_out[0] ,
    \cbx_1__1__3_chanx_right_out[1] ,
    \cbx_1__1__3_chanx_right_out[2] ,
    \cbx_1__1__3_chanx_right_out[3] ,
    \cbx_1__1__3_chanx_right_out[4] ,
    \cbx_1__1__3_chanx_right_out[5] ,
    \cbx_1__1__3_chanx_right_out[6] ,
    \cbx_1__1__3_chanx_right_out[7] ,
    \cbx_1__1__3_chanx_right_out[8] ,
    \cbx_1__1__3_chanx_right_out[9] ,
    \cbx_1__1__3_chanx_right_out[10] ,
    \cbx_1__1__3_chanx_right_out[11] ,
    \cbx_1__1__3_chanx_right_out[12] ,
    \cbx_1__1__3_chanx_right_out[13] ,
    \cbx_1__1__3_chanx_right_out[14] ,
    \cbx_1__1__3_chanx_right_out[15] ,
    \cbx_1__1__3_chanx_right_out[16] ,
    \cbx_1__1__3_chanx_right_out[17] ,
    \cbx_1__1__3_chanx_right_out[18] ,
    \cbx_1__1__3_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__3_chanx_left_out[0] ,
    \sb_1__1__3_chanx_left_out[1] ,
    \sb_1__1__3_chanx_left_out[2] ,
    \sb_1__1__3_chanx_left_out[3] ,
    \sb_1__1__3_chanx_left_out[4] ,
    \sb_1__1__3_chanx_left_out[5] ,
    \sb_1__1__3_chanx_left_out[6] ,
    \sb_1__1__3_chanx_left_out[7] ,
    \sb_1__1__3_chanx_left_out[8] ,
    \sb_1__1__3_chanx_left_out[9] ,
    \sb_1__1__3_chanx_left_out[10] ,
    \sb_1__1__3_chanx_left_out[11] ,
    \sb_1__1__3_chanx_left_out[12] ,
    \sb_1__1__3_chanx_left_out[13] ,
    \sb_1__1__3_chanx_left_out[14] ,
    \sb_1__1__3_chanx_left_out[15] ,
    \sb_1__1__3_chanx_left_out[16] ,
    \sb_1__1__3_chanx_left_out[17] ,
    \sb_1__1__3_chanx_left_out[18] ,
    \sb_1__1__3_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__10_chanx_left_out[0] ,
    \cbx_1__1__10_chanx_left_out[1] ,
    \cbx_1__1__10_chanx_left_out[2] ,
    \cbx_1__1__10_chanx_left_out[3] ,
    \cbx_1__1__10_chanx_left_out[4] ,
    \cbx_1__1__10_chanx_left_out[5] ,
    \cbx_1__1__10_chanx_left_out[6] ,
    \cbx_1__1__10_chanx_left_out[7] ,
    \cbx_1__1__10_chanx_left_out[8] ,
    \cbx_1__1__10_chanx_left_out[9] ,
    \cbx_1__1__10_chanx_left_out[10] ,
    \cbx_1__1__10_chanx_left_out[11] ,
    \cbx_1__1__10_chanx_left_out[12] ,
    \cbx_1__1__10_chanx_left_out[13] ,
    \cbx_1__1__10_chanx_left_out[14] ,
    \cbx_1__1__10_chanx_left_out[15] ,
    \cbx_1__1__10_chanx_left_out[16] ,
    \cbx_1__1__10_chanx_left_out[17] ,
    \cbx_1__1__10_chanx_left_out[18] ,
    \cbx_1__1__10_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__3_chanx_right_out[0] ,
    \sb_1__1__3_chanx_right_out[1] ,
    \sb_1__1__3_chanx_right_out[2] ,
    \sb_1__1__3_chanx_right_out[3] ,
    \sb_1__1__3_chanx_right_out[4] ,
    \sb_1__1__3_chanx_right_out[5] ,
    \sb_1__1__3_chanx_right_out[6] ,
    \sb_1__1__3_chanx_right_out[7] ,
    \sb_1__1__3_chanx_right_out[8] ,
    \sb_1__1__3_chanx_right_out[9] ,
    \sb_1__1__3_chanx_right_out[10] ,
    \sb_1__1__3_chanx_right_out[11] ,
    \sb_1__1__3_chanx_right_out[12] ,
    \sb_1__1__3_chanx_right_out[13] ,
    \sb_1__1__3_chanx_right_out[14] ,
    \sb_1__1__3_chanx_right_out[15] ,
    \sb_1__1__3_chanx_right_out[16] ,
    \sb_1__1__3_chanx_right_out[17] ,
    \sb_1__1__3_chanx_right_out[18] ,
    \sb_1__1__3_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__3_chany_top_out[0] ,
    \cby_1__1__3_chany_top_out[1] ,
    \cby_1__1__3_chany_top_out[2] ,
    \cby_1__1__3_chany_top_out[3] ,
    \cby_1__1__3_chany_top_out[4] ,
    \cby_1__1__3_chany_top_out[5] ,
    \cby_1__1__3_chany_top_out[6] ,
    \cby_1__1__3_chany_top_out[7] ,
    \cby_1__1__3_chany_top_out[8] ,
    \cby_1__1__3_chany_top_out[9] ,
    \cby_1__1__3_chany_top_out[10] ,
    \cby_1__1__3_chany_top_out[11] ,
    \cby_1__1__3_chany_top_out[12] ,
    \cby_1__1__3_chany_top_out[13] ,
    \cby_1__1__3_chany_top_out[14] ,
    \cby_1__1__3_chany_top_out[15] ,
    \cby_1__1__3_chany_top_out[16] ,
    \cby_1__1__3_chany_top_out[17] ,
    \cby_1__1__3_chany_top_out[18] ,
    \cby_1__1__3_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__3_chany_bottom_out[0] ,
    \sb_1__1__3_chany_bottom_out[1] ,
    \sb_1__1__3_chany_bottom_out[2] ,
    \sb_1__1__3_chany_bottom_out[3] ,
    \sb_1__1__3_chany_bottom_out[4] ,
    \sb_1__1__3_chany_bottom_out[5] ,
    \sb_1__1__3_chany_bottom_out[6] ,
    \sb_1__1__3_chany_bottom_out[7] ,
    \sb_1__1__3_chany_bottom_out[8] ,
    \sb_1__1__3_chany_bottom_out[9] ,
    \sb_1__1__3_chany_bottom_out[10] ,
    \sb_1__1__3_chany_bottom_out[11] ,
    \sb_1__1__3_chany_bottom_out[12] ,
    \sb_1__1__3_chany_bottom_out[13] ,
    \sb_1__1__3_chany_bottom_out[14] ,
    \sb_1__1__3_chany_bottom_out[15] ,
    \sb_1__1__3_chany_bottom_out[16] ,
    \sb_1__1__3_chany_bottom_out[17] ,
    \sb_1__1__3_chany_bottom_out[18] ,
    \sb_1__1__3_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__4_chany_bottom_out[0] ,
    \cby_1__1__4_chany_bottom_out[1] ,
    \cby_1__1__4_chany_bottom_out[2] ,
    \cby_1__1__4_chany_bottom_out[3] ,
    \cby_1__1__4_chany_bottom_out[4] ,
    \cby_1__1__4_chany_bottom_out[5] ,
    \cby_1__1__4_chany_bottom_out[6] ,
    \cby_1__1__4_chany_bottom_out[7] ,
    \cby_1__1__4_chany_bottom_out[8] ,
    \cby_1__1__4_chany_bottom_out[9] ,
    \cby_1__1__4_chany_bottom_out[10] ,
    \cby_1__1__4_chany_bottom_out[11] ,
    \cby_1__1__4_chany_bottom_out[12] ,
    \cby_1__1__4_chany_bottom_out[13] ,
    \cby_1__1__4_chany_bottom_out[14] ,
    \cby_1__1__4_chany_bottom_out[15] ,
    \cby_1__1__4_chany_bottom_out[16] ,
    \cby_1__1__4_chany_bottom_out[17] ,
    \cby_1__1__4_chany_bottom_out[18] ,
    \cby_1__1__4_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__3_chany_top_out[0] ,
    \sb_1__1__3_chany_top_out[1] ,
    \sb_1__1__3_chany_top_out[2] ,
    \sb_1__1__3_chany_top_out[3] ,
    \sb_1__1__3_chany_top_out[4] ,
    \sb_1__1__3_chany_top_out[5] ,
    \sb_1__1__3_chany_top_out[6] ,
    \sb_1__1__3_chany_top_out[7] ,
    \sb_1__1__3_chany_top_out[8] ,
    \sb_1__1__3_chany_top_out[9] ,
    \sb_1__1__3_chany_top_out[10] ,
    \sb_1__1__3_chany_top_out[11] ,
    \sb_1__1__3_chany_top_out[12] ,
    \sb_1__1__3_chany_top_out[13] ,
    \sb_1__1__3_chany_top_out[14] ,
    \sb_1__1__3_chany_top_out[15] ,
    \sb_1__1__3_chany_top_out[16] ,
    \sb_1__1__3_chany_top_out[17] ,
    \sb_1__1__3_chany_top_out[18] ,
    \sb_1__1__3_chany_top_out[19] }));
 sb_1__1_ sb_1__5_ (.bottom_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__11_ccff_tail),
    .ccff_tail(sb_1__1__4_ccff_tail),
    .clk_1_E_out(\clk_1_wires[15] ),
    .clk_1_N_in(\clk_2_wires[21] ),
    .clk_1_W_out(\clk_1_wires[16] ),
    .left_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[28] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[15] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[21] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[16] ),
    .right_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__4_chanx_right_out[0] ,
    \cbx_1__1__4_chanx_right_out[1] ,
    \cbx_1__1__4_chanx_right_out[2] ,
    \cbx_1__1__4_chanx_right_out[3] ,
    \cbx_1__1__4_chanx_right_out[4] ,
    \cbx_1__1__4_chanx_right_out[5] ,
    \cbx_1__1__4_chanx_right_out[6] ,
    \cbx_1__1__4_chanx_right_out[7] ,
    \cbx_1__1__4_chanx_right_out[8] ,
    \cbx_1__1__4_chanx_right_out[9] ,
    \cbx_1__1__4_chanx_right_out[10] ,
    \cbx_1__1__4_chanx_right_out[11] ,
    \cbx_1__1__4_chanx_right_out[12] ,
    \cbx_1__1__4_chanx_right_out[13] ,
    \cbx_1__1__4_chanx_right_out[14] ,
    \cbx_1__1__4_chanx_right_out[15] ,
    \cbx_1__1__4_chanx_right_out[16] ,
    \cbx_1__1__4_chanx_right_out[17] ,
    \cbx_1__1__4_chanx_right_out[18] ,
    \cbx_1__1__4_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__4_chanx_left_out[0] ,
    \sb_1__1__4_chanx_left_out[1] ,
    \sb_1__1__4_chanx_left_out[2] ,
    \sb_1__1__4_chanx_left_out[3] ,
    \sb_1__1__4_chanx_left_out[4] ,
    \sb_1__1__4_chanx_left_out[5] ,
    \sb_1__1__4_chanx_left_out[6] ,
    \sb_1__1__4_chanx_left_out[7] ,
    \sb_1__1__4_chanx_left_out[8] ,
    \sb_1__1__4_chanx_left_out[9] ,
    \sb_1__1__4_chanx_left_out[10] ,
    \sb_1__1__4_chanx_left_out[11] ,
    \sb_1__1__4_chanx_left_out[12] ,
    \sb_1__1__4_chanx_left_out[13] ,
    \sb_1__1__4_chanx_left_out[14] ,
    \sb_1__1__4_chanx_left_out[15] ,
    \sb_1__1__4_chanx_left_out[16] ,
    \sb_1__1__4_chanx_left_out[17] ,
    \sb_1__1__4_chanx_left_out[18] ,
    \sb_1__1__4_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__11_chanx_left_out[0] ,
    \cbx_1__1__11_chanx_left_out[1] ,
    \cbx_1__1__11_chanx_left_out[2] ,
    \cbx_1__1__11_chanx_left_out[3] ,
    \cbx_1__1__11_chanx_left_out[4] ,
    \cbx_1__1__11_chanx_left_out[5] ,
    \cbx_1__1__11_chanx_left_out[6] ,
    \cbx_1__1__11_chanx_left_out[7] ,
    \cbx_1__1__11_chanx_left_out[8] ,
    \cbx_1__1__11_chanx_left_out[9] ,
    \cbx_1__1__11_chanx_left_out[10] ,
    \cbx_1__1__11_chanx_left_out[11] ,
    \cbx_1__1__11_chanx_left_out[12] ,
    \cbx_1__1__11_chanx_left_out[13] ,
    \cbx_1__1__11_chanx_left_out[14] ,
    \cbx_1__1__11_chanx_left_out[15] ,
    \cbx_1__1__11_chanx_left_out[16] ,
    \cbx_1__1__11_chanx_left_out[17] ,
    \cbx_1__1__11_chanx_left_out[18] ,
    \cbx_1__1__11_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__4_chanx_right_out[0] ,
    \sb_1__1__4_chanx_right_out[1] ,
    \sb_1__1__4_chanx_right_out[2] ,
    \sb_1__1__4_chanx_right_out[3] ,
    \sb_1__1__4_chanx_right_out[4] ,
    \sb_1__1__4_chanx_right_out[5] ,
    \sb_1__1__4_chanx_right_out[6] ,
    \sb_1__1__4_chanx_right_out[7] ,
    \sb_1__1__4_chanx_right_out[8] ,
    \sb_1__1__4_chanx_right_out[9] ,
    \sb_1__1__4_chanx_right_out[10] ,
    \sb_1__1__4_chanx_right_out[11] ,
    \sb_1__1__4_chanx_right_out[12] ,
    \sb_1__1__4_chanx_right_out[13] ,
    \sb_1__1__4_chanx_right_out[14] ,
    \sb_1__1__4_chanx_right_out[15] ,
    \sb_1__1__4_chanx_right_out[16] ,
    \sb_1__1__4_chanx_right_out[17] ,
    \sb_1__1__4_chanx_right_out[18] ,
    \sb_1__1__4_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__4_chany_top_out[0] ,
    \cby_1__1__4_chany_top_out[1] ,
    \cby_1__1__4_chany_top_out[2] ,
    \cby_1__1__4_chany_top_out[3] ,
    \cby_1__1__4_chany_top_out[4] ,
    \cby_1__1__4_chany_top_out[5] ,
    \cby_1__1__4_chany_top_out[6] ,
    \cby_1__1__4_chany_top_out[7] ,
    \cby_1__1__4_chany_top_out[8] ,
    \cby_1__1__4_chany_top_out[9] ,
    \cby_1__1__4_chany_top_out[10] ,
    \cby_1__1__4_chany_top_out[11] ,
    \cby_1__1__4_chany_top_out[12] ,
    \cby_1__1__4_chany_top_out[13] ,
    \cby_1__1__4_chany_top_out[14] ,
    \cby_1__1__4_chany_top_out[15] ,
    \cby_1__1__4_chany_top_out[16] ,
    \cby_1__1__4_chany_top_out[17] ,
    \cby_1__1__4_chany_top_out[18] ,
    \cby_1__1__4_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__4_chany_bottom_out[0] ,
    \sb_1__1__4_chany_bottom_out[1] ,
    \sb_1__1__4_chany_bottom_out[2] ,
    \sb_1__1__4_chany_bottom_out[3] ,
    \sb_1__1__4_chany_bottom_out[4] ,
    \sb_1__1__4_chany_bottom_out[5] ,
    \sb_1__1__4_chany_bottom_out[6] ,
    \sb_1__1__4_chany_bottom_out[7] ,
    \sb_1__1__4_chany_bottom_out[8] ,
    \sb_1__1__4_chany_bottom_out[9] ,
    \sb_1__1__4_chany_bottom_out[10] ,
    \sb_1__1__4_chany_bottom_out[11] ,
    \sb_1__1__4_chany_bottom_out[12] ,
    \sb_1__1__4_chany_bottom_out[13] ,
    \sb_1__1__4_chany_bottom_out[14] ,
    \sb_1__1__4_chany_bottom_out[15] ,
    \sb_1__1__4_chany_bottom_out[16] ,
    \sb_1__1__4_chany_bottom_out[17] ,
    \sb_1__1__4_chany_bottom_out[18] ,
    \sb_1__1__4_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__5_chany_bottom_out[0] ,
    \cby_1__1__5_chany_bottom_out[1] ,
    \cby_1__1__5_chany_bottom_out[2] ,
    \cby_1__1__5_chany_bottom_out[3] ,
    \cby_1__1__5_chany_bottom_out[4] ,
    \cby_1__1__5_chany_bottom_out[5] ,
    \cby_1__1__5_chany_bottom_out[6] ,
    \cby_1__1__5_chany_bottom_out[7] ,
    \cby_1__1__5_chany_bottom_out[8] ,
    \cby_1__1__5_chany_bottom_out[9] ,
    \cby_1__1__5_chany_bottom_out[10] ,
    \cby_1__1__5_chany_bottom_out[11] ,
    \cby_1__1__5_chany_bottom_out[12] ,
    \cby_1__1__5_chany_bottom_out[13] ,
    \cby_1__1__5_chany_bottom_out[14] ,
    \cby_1__1__5_chany_bottom_out[15] ,
    \cby_1__1__5_chany_bottom_out[16] ,
    \cby_1__1__5_chany_bottom_out[17] ,
    \cby_1__1__5_chany_bottom_out[18] ,
    \cby_1__1__5_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__4_chany_top_out[0] ,
    \sb_1__1__4_chany_top_out[1] ,
    \sb_1__1__4_chany_top_out[2] ,
    \sb_1__1__4_chany_top_out[3] ,
    \sb_1__1__4_chany_top_out[4] ,
    \sb_1__1__4_chany_top_out[5] ,
    \sb_1__1__4_chany_top_out[6] ,
    \sb_1__1__4_chany_top_out[7] ,
    \sb_1__1__4_chany_top_out[8] ,
    \sb_1__1__4_chany_top_out[9] ,
    \sb_1__1__4_chany_top_out[10] ,
    \sb_1__1__4_chany_top_out[11] ,
    \sb_1__1__4_chany_top_out[12] ,
    \sb_1__1__4_chany_top_out[13] ,
    \sb_1__1__4_chany_top_out[14] ,
    \sb_1__1__4_chany_top_out[15] ,
    \sb_1__1__4_chany_top_out[16] ,
    \sb_1__1__4_chany_top_out[17] ,
    \sb_1__1__4_chany_top_out[18] ,
    \sb_1__1__4_chany_top_out[19] }));
 sb_1__1_ sb_1__6_ (.bottom_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__12_ccff_tail),
    .ccff_tail(sb_1__1__5_ccff_tail),
    .clk_2_N_in(\clk_2_wires[17] ),
    .clk_2_N_out(\clk_2_wires[18] ),
    .clk_2_S_out(\clk_2_wires[20] ),
    .left_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[33] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[17] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[18] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[20] ),
    .right_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__5_chanx_right_out[0] ,
    \cbx_1__1__5_chanx_right_out[1] ,
    \cbx_1__1__5_chanx_right_out[2] ,
    \cbx_1__1__5_chanx_right_out[3] ,
    \cbx_1__1__5_chanx_right_out[4] ,
    \cbx_1__1__5_chanx_right_out[5] ,
    \cbx_1__1__5_chanx_right_out[6] ,
    \cbx_1__1__5_chanx_right_out[7] ,
    \cbx_1__1__5_chanx_right_out[8] ,
    \cbx_1__1__5_chanx_right_out[9] ,
    \cbx_1__1__5_chanx_right_out[10] ,
    \cbx_1__1__5_chanx_right_out[11] ,
    \cbx_1__1__5_chanx_right_out[12] ,
    \cbx_1__1__5_chanx_right_out[13] ,
    \cbx_1__1__5_chanx_right_out[14] ,
    \cbx_1__1__5_chanx_right_out[15] ,
    \cbx_1__1__5_chanx_right_out[16] ,
    \cbx_1__1__5_chanx_right_out[17] ,
    \cbx_1__1__5_chanx_right_out[18] ,
    \cbx_1__1__5_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__5_chanx_left_out[0] ,
    \sb_1__1__5_chanx_left_out[1] ,
    \sb_1__1__5_chanx_left_out[2] ,
    \sb_1__1__5_chanx_left_out[3] ,
    \sb_1__1__5_chanx_left_out[4] ,
    \sb_1__1__5_chanx_left_out[5] ,
    \sb_1__1__5_chanx_left_out[6] ,
    \sb_1__1__5_chanx_left_out[7] ,
    \sb_1__1__5_chanx_left_out[8] ,
    \sb_1__1__5_chanx_left_out[9] ,
    \sb_1__1__5_chanx_left_out[10] ,
    \sb_1__1__5_chanx_left_out[11] ,
    \sb_1__1__5_chanx_left_out[12] ,
    \sb_1__1__5_chanx_left_out[13] ,
    \sb_1__1__5_chanx_left_out[14] ,
    \sb_1__1__5_chanx_left_out[15] ,
    \sb_1__1__5_chanx_left_out[16] ,
    \sb_1__1__5_chanx_left_out[17] ,
    \sb_1__1__5_chanx_left_out[18] ,
    \sb_1__1__5_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__12_chanx_left_out[0] ,
    \cbx_1__1__12_chanx_left_out[1] ,
    \cbx_1__1__12_chanx_left_out[2] ,
    \cbx_1__1__12_chanx_left_out[3] ,
    \cbx_1__1__12_chanx_left_out[4] ,
    \cbx_1__1__12_chanx_left_out[5] ,
    \cbx_1__1__12_chanx_left_out[6] ,
    \cbx_1__1__12_chanx_left_out[7] ,
    \cbx_1__1__12_chanx_left_out[8] ,
    \cbx_1__1__12_chanx_left_out[9] ,
    \cbx_1__1__12_chanx_left_out[10] ,
    \cbx_1__1__12_chanx_left_out[11] ,
    \cbx_1__1__12_chanx_left_out[12] ,
    \cbx_1__1__12_chanx_left_out[13] ,
    \cbx_1__1__12_chanx_left_out[14] ,
    \cbx_1__1__12_chanx_left_out[15] ,
    \cbx_1__1__12_chanx_left_out[16] ,
    \cbx_1__1__12_chanx_left_out[17] ,
    \cbx_1__1__12_chanx_left_out[18] ,
    \cbx_1__1__12_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__5_chanx_right_out[0] ,
    \sb_1__1__5_chanx_right_out[1] ,
    \sb_1__1__5_chanx_right_out[2] ,
    \sb_1__1__5_chanx_right_out[3] ,
    \sb_1__1__5_chanx_right_out[4] ,
    \sb_1__1__5_chanx_right_out[5] ,
    \sb_1__1__5_chanx_right_out[6] ,
    \sb_1__1__5_chanx_right_out[7] ,
    \sb_1__1__5_chanx_right_out[8] ,
    \sb_1__1__5_chanx_right_out[9] ,
    \sb_1__1__5_chanx_right_out[10] ,
    \sb_1__1__5_chanx_right_out[11] ,
    \sb_1__1__5_chanx_right_out[12] ,
    \sb_1__1__5_chanx_right_out[13] ,
    \sb_1__1__5_chanx_right_out[14] ,
    \sb_1__1__5_chanx_right_out[15] ,
    \sb_1__1__5_chanx_right_out[16] ,
    \sb_1__1__5_chanx_right_out[17] ,
    \sb_1__1__5_chanx_right_out[18] ,
    \sb_1__1__5_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__5_chany_top_out[0] ,
    \cby_1__1__5_chany_top_out[1] ,
    \cby_1__1__5_chany_top_out[2] ,
    \cby_1__1__5_chany_top_out[3] ,
    \cby_1__1__5_chany_top_out[4] ,
    \cby_1__1__5_chany_top_out[5] ,
    \cby_1__1__5_chany_top_out[6] ,
    \cby_1__1__5_chany_top_out[7] ,
    \cby_1__1__5_chany_top_out[8] ,
    \cby_1__1__5_chany_top_out[9] ,
    \cby_1__1__5_chany_top_out[10] ,
    \cby_1__1__5_chany_top_out[11] ,
    \cby_1__1__5_chany_top_out[12] ,
    \cby_1__1__5_chany_top_out[13] ,
    \cby_1__1__5_chany_top_out[14] ,
    \cby_1__1__5_chany_top_out[15] ,
    \cby_1__1__5_chany_top_out[16] ,
    \cby_1__1__5_chany_top_out[17] ,
    \cby_1__1__5_chany_top_out[18] ,
    \cby_1__1__5_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__5_chany_bottom_out[0] ,
    \sb_1__1__5_chany_bottom_out[1] ,
    \sb_1__1__5_chany_bottom_out[2] ,
    \sb_1__1__5_chany_bottom_out[3] ,
    \sb_1__1__5_chany_bottom_out[4] ,
    \sb_1__1__5_chany_bottom_out[5] ,
    \sb_1__1__5_chany_bottom_out[6] ,
    \sb_1__1__5_chany_bottom_out[7] ,
    \sb_1__1__5_chany_bottom_out[8] ,
    \sb_1__1__5_chany_bottom_out[9] ,
    \sb_1__1__5_chany_bottom_out[10] ,
    \sb_1__1__5_chany_bottom_out[11] ,
    \sb_1__1__5_chany_bottom_out[12] ,
    \sb_1__1__5_chany_bottom_out[13] ,
    \sb_1__1__5_chany_bottom_out[14] ,
    \sb_1__1__5_chany_bottom_out[15] ,
    \sb_1__1__5_chany_bottom_out[16] ,
    \sb_1__1__5_chany_bottom_out[17] ,
    \sb_1__1__5_chany_bottom_out[18] ,
    \sb_1__1__5_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__6_chany_bottom_out[0] ,
    \cby_1__1__6_chany_bottom_out[1] ,
    \cby_1__1__6_chany_bottom_out[2] ,
    \cby_1__1__6_chany_bottom_out[3] ,
    \cby_1__1__6_chany_bottom_out[4] ,
    \cby_1__1__6_chany_bottom_out[5] ,
    \cby_1__1__6_chany_bottom_out[6] ,
    \cby_1__1__6_chany_bottom_out[7] ,
    \cby_1__1__6_chany_bottom_out[8] ,
    \cby_1__1__6_chany_bottom_out[9] ,
    \cby_1__1__6_chany_bottom_out[10] ,
    \cby_1__1__6_chany_bottom_out[11] ,
    \cby_1__1__6_chany_bottom_out[12] ,
    \cby_1__1__6_chany_bottom_out[13] ,
    \cby_1__1__6_chany_bottom_out[14] ,
    \cby_1__1__6_chany_bottom_out[15] ,
    \cby_1__1__6_chany_bottom_out[16] ,
    \cby_1__1__6_chany_bottom_out[17] ,
    \cby_1__1__6_chany_bottom_out[18] ,
    \cby_1__1__6_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__5_chany_top_out[0] ,
    \sb_1__1__5_chany_top_out[1] ,
    \sb_1__1__5_chany_top_out[2] ,
    \sb_1__1__5_chany_top_out[3] ,
    \sb_1__1__5_chany_top_out[4] ,
    \sb_1__1__5_chany_top_out[5] ,
    \sb_1__1__5_chany_top_out[6] ,
    \sb_1__1__5_chany_top_out[7] ,
    \sb_1__1__5_chany_top_out[8] ,
    \sb_1__1__5_chany_top_out[9] ,
    \sb_1__1__5_chany_top_out[10] ,
    \sb_1__1__5_chany_top_out[11] ,
    \sb_1__1__5_chany_top_out[12] ,
    \sb_1__1__5_chany_top_out[13] ,
    \sb_1__1__5_chany_top_out[14] ,
    \sb_1__1__5_chany_top_out[15] ,
    \sb_1__1__5_chany_top_out[16] ,
    \sb_1__1__5_chany_top_out[17] ,
    \sb_1__1__5_chany_top_out[18] ,
    \sb_1__1__5_chany_top_out[19] }));
 sb_1__1_ sb_1__7_ (.bottom_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__13_ccff_tail),
    .ccff_tail(sb_1__1__6_ccff_tail),
    .clk_1_E_out(\clk_1_wires[22] ),
    .clk_1_N_in(\clk_2_wires[19] ),
    .clk_1_W_out(\clk_1_wires[23] ),
    .left_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[38] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[22] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[19] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[23] ),
    .right_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__6_chanx_right_out[0] ,
    \cbx_1__1__6_chanx_right_out[1] ,
    \cbx_1__1__6_chanx_right_out[2] ,
    \cbx_1__1__6_chanx_right_out[3] ,
    \cbx_1__1__6_chanx_right_out[4] ,
    \cbx_1__1__6_chanx_right_out[5] ,
    \cbx_1__1__6_chanx_right_out[6] ,
    \cbx_1__1__6_chanx_right_out[7] ,
    \cbx_1__1__6_chanx_right_out[8] ,
    \cbx_1__1__6_chanx_right_out[9] ,
    \cbx_1__1__6_chanx_right_out[10] ,
    \cbx_1__1__6_chanx_right_out[11] ,
    \cbx_1__1__6_chanx_right_out[12] ,
    \cbx_1__1__6_chanx_right_out[13] ,
    \cbx_1__1__6_chanx_right_out[14] ,
    \cbx_1__1__6_chanx_right_out[15] ,
    \cbx_1__1__6_chanx_right_out[16] ,
    \cbx_1__1__6_chanx_right_out[17] ,
    \cbx_1__1__6_chanx_right_out[18] ,
    \cbx_1__1__6_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__6_chanx_left_out[0] ,
    \sb_1__1__6_chanx_left_out[1] ,
    \sb_1__1__6_chanx_left_out[2] ,
    \sb_1__1__6_chanx_left_out[3] ,
    \sb_1__1__6_chanx_left_out[4] ,
    \sb_1__1__6_chanx_left_out[5] ,
    \sb_1__1__6_chanx_left_out[6] ,
    \sb_1__1__6_chanx_left_out[7] ,
    \sb_1__1__6_chanx_left_out[8] ,
    \sb_1__1__6_chanx_left_out[9] ,
    \sb_1__1__6_chanx_left_out[10] ,
    \sb_1__1__6_chanx_left_out[11] ,
    \sb_1__1__6_chanx_left_out[12] ,
    \sb_1__1__6_chanx_left_out[13] ,
    \sb_1__1__6_chanx_left_out[14] ,
    \sb_1__1__6_chanx_left_out[15] ,
    \sb_1__1__6_chanx_left_out[16] ,
    \sb_1__1__6_chanx_left_out[17] ,
    \sb_1__1__6_chanx_left_out[18] ,
    \sb_1__1__6_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__13_chanx_left_out[0] ,
    \cbx_1__1__13_chanx_left_out[1] ,
    \cbx_1__1__13_chanx_left_out[2] ,
    \cbx_1__1__13_chanx_left_out[3] ,
    \cbx_1__1__13_chanx_left_out[4] ,
    \cbx_1__1__13_chanx_left_out[5] ,
    \cbx_1__1__13_chanx_left_out[6] ,
    \cbx_1__1__13_chanx_left_out[7] ,
    \cbx_1__1__13_chanx_left_out[8] ,
    \cbx_1__1__13_chanx_left_out[9] ,
    \cbx_1__1__13_chanx_left_out[10] ,
    \cbx_1__1__13_chanx_left_out[11] ,
    \cbx_1__1__13_chanx_left_out[12] ,
    \cbx_1__1__13_chanx_left_out[13] ,
    \cbx_1__1__13_chanx_left_out[14] ,
    \cbx_1__1__13_chanx_left_out[15] ,
    \cbx_1__1__13_chanx_left_out[16] ,
    \cbx_1__1__13_chanx_left_out[17] ,
    \cbx_1__1__13_chanx_left_out[18] ,
    \cbx_1__1__13_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__6_chanx_right_out[0] ,
    \sb_1__1__6_chanx_right_out[1] ,
    \sb_1__1__6_chanx_right_out[2] ,
    \sb_1__1__6_chanx_right_out[3] ,
    \sb_1__1__6_chanx_right_out[4] ,
    \sb_1__1__6_chanx_right_out[5] ,
    \sb_1__1__6_chanx_right_out[6] ,
    \sb_1__1__6_chanx_right_out[7] ,
    \sb_1__1__6_chanx_right_out[8] ,
    \sb_1__1__6_chanx_right_out[9] ,
    \sb_1__1__6_chanx_right_out[10] ,
    \sb_1__1__6_chanx_right_out[11] ,
    \sb_1__1__6_chanx_right_out[12] ,
    \sb_1__1__6_chanx_right_out[13] ,
    \sb_1__1__6_chanx_right_out[14] ,
    \sb_1__1__6_chanx_right_out[15] ,
    \sb_1__1__6_chanx_right_out[16] ,
    \sb_1__1__6_chanx_right_out[17] ,
    \sb_1__1__6_chanx_right_out[18] ,
    \sb_1__1__6_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__6_chany_top_out[0] ,
    \cby_1__1__6_chany_top_out[1] ,
    \cby_1__1__6_chany_top_out[2] ,
    \cby_1__1__6_chany_top_out[3] ,
    \cby_1__1__6_chany_top_out[4] ,
    \cby_1__1__6_chany_top_out[5] ,
    \cby_1__1__6_chany_top_out[6] ,
    \cby_1__1__6_chany_top_out[7] ,
    \cby_1__1__6_chany_top_out[8] ,
    \cby_1__1__6_chany_top_out[9] ,
    \cby_1__1__6_chany_top_out[10] ,
    \cby_1__1__6_chany_top_out[11] ,
    \cby_1__1__6_chany_top_out[12] ,
    \cby_1__1__6_chany_top_out[13] ,
    \cby_1__1__6_chany_top_out[14] ,
    \cby_1__1__6_chany_top_out[15] ,
    \cby_1__1__6_chany_top_out[16] ,
    \cby_1__1__6_chany_top_out[17] ,
    \cby_1__1__6_chany_top_out[18] ,
    \cby_1__1__6_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__6_chany_bottom_out[0] ,
    \sb_1__1__6_chany_bottom_out[1] ,
    \sb_1__1__6_chany_bottom_out[2] ,
    \sb_1__1__6_chany_bottom_out[3] ,
    \sb_1__1__6_chany_bottom_out[4] ,
    \sb_1__1__6_chany_bottom_out[5] ,
    \sb_1__1__6_chany_bottom_out[6] ,
    \sb_1__1__6_chany_bottom_out[7] ,
    \sb_1__1__6_chany_bottom_out[8] ,
    \sb_1__1__6_chany_bottom_out[9] ,
    \sb_1__1__6_chany_bottom_out[10] ,
    \sb_1__1__6_chany_bottom_out[11] ,
    \sb_1__1__6_chany_bottom_out[12] ,
    \sb_1__1__6_chany_bottom_out[13] ,
    \sb_1__1__6_chany_bottom_out[14] ,
    \sb_1__1__6_chany_bottom_out[15] ,
    \sb_1__1__6_chany_bottom_out[16] ,
    \sb_1__1__6_chany_bottom_out[17] ,
    \sb_1__1__6_chany_bottom_out[18] ,
    \sb_1__1__6_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__7_chany_bottom_out[0] ,
    \cby_1__1__7_chany_bottom_out[1] ,
    \cby_1__1__7_chany_bottom_out[2] ,
    \cby_1__1__7_chany_bottom_out[3] ,
    \cby_1__1__7_chany_bottom_out[4] ,
    \cby_1__1__7_chany_bottom_out[5] ,
    \cby_1__1__7_chany_bottom_out[6] ,
    \cby_1__1__7_chany_bottom_out[7] ,
    \cby_1__1__7_chany_bottom_out[8] ,
    \cby_1__1__7_chany_bottom_out[9] ,
    \cby_1__1__7_chany_bottom_out[10] ,
    \cby_1__1__7_chany_bottom_out[11] ,
    \cby_1__1__7_chany_bottom_out[12] ,
    \cby_1__1__7_chany_bottom_out[13] ,
    \cby_1__1__7_chany_bottom_out[14] ,
    \cby_1__1__7_chany_bottom_out[15] ,
    \cby_1__1__7_chany_bottom_out[16] ,
    \cby_1__1__7_chany_bottom_out[17] ,
    \cby_1__1__7_chany_bottom_out[18] ,
    \cby_1__1__7_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__6_chany_top_out[0] ,
    \sb_1__1__6_chany_top_out[1] ,
    \sb_1__1__6_chany_top_out[2] ,
    \sb_1__1__6_chany_top_out[3] ,
    \sb_1__1__6_chany_top_out[4] ,
    \sb_1__1__6_chany_top_out[5] ,
    \sb_1__1__6_chany_top_out[6] ,
    \sb_1__1__6_chany_top_out[7] ,
    \sb_1__1__6_chany_top_out[8] ,
    \sb_1__1__6_chany_top_out[9] ,
    \sb_1__1__6_chany_top_out[10] ,
    \sb_1__1__6_chany_top_out[11] ,
    \sb_1__1__6_chany_top_out[12] ,
    \sb_1__1__6_chany_top_out[13] ,
    \sb_1__1__6_chany_top_out[14] ,
    \sb_1__1__6_chany_top_out[15] ,
    \sb_1__1__6_chany_top_out[16] ,
    \sb_1__1__6_chany_top_out[17] ,
    \sb_1__1__6_chany_top_out[18] ,
    \sb_1__1__6_chany_top_out[19] }));
 sb_1__2_ sb_1__8_ (.bottom_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_upper),
    .ccff_head(grid_io_top_1_ccff_tail),
    .ccff_tail(sb_1__8__0_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[40] ),
    .right_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__0_chanx_right_out[0] ,
    \cbx_1__8__0_chanx_right_out[1] ,
    \cbx_1__8__0_chanx_right_out[2] ,
    \cbx_1__8__0_chanx_right_out[3] ,
    \cbx_1__8__0_chanx_right_out[4] ,
    \cbx_1__8__0_chanx_right_out[5] ,
    \cbx_1__8__0_chanx_right_out[6] ,
    \cbx_1__8__0_chanx_right_out[7] ,
    \cbx_1__8__0_chanx_right_out[8] ,
    \cbx_1__8__0_chanx_right_out[9] ,
    \cbx_1__8__0_chanx_right_out[10] ,
    \cbx_1__8__0_chanx_right_out[11] ,
    \cbx_1__8__0_chanx_right_out[12] ,
    \cbx_1__8__0_chanx_right_out[13] ,
    \cbx_1__8__0_chanx_right_out[14] ,
    \cbx_1__8__0_chanx_right_out[15] ,
    \cbx_1__8__0_chanx_right_out[16] ,
    \cbx_1__8__0_chanx_right_out[17] ,
    \cbx_1__8__0_chanx_right_out[18] ,
    \cbx_1__8__0_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__8__0_chanx_left_out[0] ,
    \sb_1__8__0_chanx_left_out[1] ,
    \sb_1__8__0_chanx_left_out[2] ,
    \sb_1__8__0_chanx_left_out[3] ,
    \sb_1__8__0_chanx_left_out[4] ,
    \sb_1__8__0_chanx_left_out[5] ,
    \sb_1__8__0_chanx_left_out[6] ,
    \sb_1__8__0_chanx_left_out[7] ,
    \sb_1__8__0_chanx_left_out[8] ,
    \sb_1__8__0_chanx_left_out[9] ,
    \sb_1__8__0_chanx_left_out[10] ,
    \sb_1__8__0_chanx_left_out[11] ,
    \sb_1__8__0_chanx_left_out[12] ,
    \sb_1__8__0_chanx_left_out[13] ,
    \sb_1__8__0_chanx_left_out[14] ,
    \sb_1__8__0_chanx_left_out[15] ,
    \sb_1__8__0_chanx_left_out[16] ,
    \sb_1__8__0_chanx_left_out[17] ,
    \sb_1__8__0_chanx_left_out[18] ,
    \sb_1__8__0_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__8__1_chanx_left_out[0] ,
    \cbx_1__8__1_chanx_left_out[1] ,
    \cbx_1__8__1_chanx_left_out[2] ,
    \cbx_1__8__1_chanx_left_out[3] ,
    \cbx_1__8__1_chanx_left_out[4] ,
    \cbx_1__8__1_chanx_left_out[5] ,
    \cbx_1__8__1_chanx_left_out[6] ,
    \cbx_1__8__1_chanx_left_out[7] ,
    \cbx_1__8__1_chanx_left_out[8] ,
    \cbx_1__8__1_chanx_left_out[9] ,
    \cbx_1__8__1_chanx_left_out[10] ,
    \cbx_1__8__1_chanx_left_out[11] ,
    \cbx_1__8__1_chanx_left_out[12] ,
    \cbx_1__8__1_chanx_left_out[13] ,
    \cbx_1__8__1_chanx_left_out[14] ,
    \cbx_1__8__1_chanx_left_out[15] ,
    \cbx_1__8__1_chanx_left_out[16] ,
    \cbx_1__8__1_chanx_left_out[17] ,
    \cbx_1__8__1_chanx_left_out[18] ,
    \cbx_1__8__1_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__8__0_chanx_right_out[0] ,
    \sb_1__8__0_chanx_right_out[1] ,
    \sb_1__8__0_chanx_right_out[2] ,
    \sb_1__8__0_chanx_right_out[3] ,
    \sb_1__8__0_chanx_right_out[4] ,
    \sb_1__8__0_chanx_right_out[5] ,
    \sb_1__8__0_chanx_right_out[6] ,
    \sb_1__8__0_chanx_right_out[7] ,
    \sb_1__8__0_chanx_right_out[8] ,
    \sb_1__8__0_chanx_right_out[9] ,
    \sb_1__8__0_chanx_right_out[10] ,
    \sb_1__8__0_chanx_right_out[11] ,
    \sb_1__8__0_chanx_right_out[12] ,
    \sb_1__8__0_chanx_right_out[13] ,
    \sb_1__8__0_chanx_right_out[14] ,
    \sb_1__8__0_chanx_right_out[15] ,
    \sb_1__8__0_chanx_right_out[16] ,
    \sb_1__8__0_chanx_right_out[17] ,
    \sb_1__8__0_chanx_right_out[18] ,
    \sb_1__8__0_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__7_chany_top_out[0] ,
    \cby_1__1__7_chany_top_out[1] ,
    \cby_1__1__7_chany_top_out[2] ,
    \cby_1__1__7_chany_top_out[3] ,
    \cby_1__1__7_chany_top_out[4] ,
    \cby_1__1__7_chany_top_out[5] ,
    \cby_1__1__7_chany_top_out[6] ,
    \cby_1__1__7_chany_top_out[7] ,
    \cby_1__1__7_chany_top_out[8] ,
    \cby_1__1__7_chany_top_out[9] ,
    \cby_1__1__7_chany_top_out[10] ,
    \cby_1__1__7_chany_top_out[11] ,
    \cby_1__1__7_chany_top_out[12] ,
    \cby_1__1__7_chany_top_out[13] ,
    \cby_1__1__7_chany_top_out[14] ,
    \cby_1__1__7_chany_top_out[15] ,
    \cby_1__1__7_chany_top_out[16] ,
    \cby_1__1__7_chany_top_out[17] ,
    \cby_1__1__7_chany_top_out[18] ,
    \cby_1__1__7_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__8__0_chany_bottom_out[0] ,
    \sb_1__8__0_chany_bottom_out[1] ,
    \sb_1__8__0_chany_bottom_out[2] ,
    \sb_1__8__0_chany_bottom_out[3] ,
    \sb_1__8__0_chany_bottom_out[4] ,
    \sb_1__8__0_chany_bottom_out[5] ,
    \sb_1__8__0_chany_bottom_out[6] ,
    \sb_1__8__0_chany_bottom_out[7] ,
    \sb_1__8__0_chany_bottom_out[8] ,
    \sb_1__8__0_chany_bottom_out[9] ,
    \sb_1__8__0_chany_bottom_out[10] ,
    \sb_1__8__0_chany_bottom_out[11] ,
    \sb_1__8__0_chany_bottom_out[12] ,
    \sb_1__8__0_chany_bottom_out[13] ,
    \sb_1__8__0_chany_bottom_out[14] ,
    \sb_1__8__0_chany_bottom_out[15] ,
    \sb_1__8__0_chany_bottom_out[16] ,
    \sb_1__8__0_chany_bottom_out[17] ,
    \sb_1__8__0_chany_bottom_out[18] ,
    \sb_1__8__0_chany_bottom_out[19] }));
 sb_1__0_ sb_2__0_ (.ccff_head(grid_io_bottom_5_ccff_tail),
    .ccff_tail(sb_1__0__1_ccff_tail),
    .left_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[45] ),
    .right_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__1_chanx_right_out[0] ,
    \cbx_1__0__1_chanx_right_out[1] ,
    \cbx_1__0__1_chanx_right_out[2] ,
    \cbx_1__0__1_chanx_right_out[3] ,
    \cbx_1__0__1_chanx_right_out[4] ,
    \cbx_1__0__1_chanx_right_out[5] ,
    \cbx_1__0__1_chanx_right_out[6] ,
    \cbx_1__0__1_chanx_right_out[7] ,
    \cbx_1__0__1_chanx_right_out[8] ,
    \cbx_1__0__1_chanx_right_out[9] ,
    \cbx_1__0__1_chanx_right_out[10] ,
    \cbx_1__0__1_chanx_right_out[11] ,
    \cbx_1__0__1_chanx_right_out[12] ,
    \cbx_1__0__1_chanx_right_out[13] ,
    \cbx_1__0__1_chanx_right_out[14] ,
    \cbx_1__0__1_chanx_right_out[15] ,
    \cbx_1__0__1_chanx_right_out[16] ,
    \cbx_1__0__1_chanx_right_out[17] ,
    \cbx_1__0__1_chanx_right_out[18] ,
    \cbx_1__0__1_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__0__1_chanx_left_out[0] ,
    \sb_1__0__1_chanx_left_out[1] ,
    \sb_1__0__1_chanx_left_out[2] ,
    \sb_1__0__1_chanx_left_out[3] ,
    \sb_1__0__1_chanx_left_out[4] ,
    \sb_1__0__1_chanx_left_out[5] ,
    \sb_1__0__1_chanx_left_out[6] ,
    \sb_1__0__1_chanx_left_out[7] ,
    \sb_1__0__1_chanx_left_out[8] ,
    \sb_1__0__1_chanx_left_out[9] ,
    \sb_1__0__1_chanx_left_out[10] ,
    \sb_1__0__1_chanx_left_out[11] ,
    \sb_1__0__1_chanx_left_out[12] ,
    \sb_1__0__1_chanx_left_out[13] ,
    \sb_1__0__1_chanx_left_out[14] ,
    \sb_1__0__1_chanx_left_out[15] ,
    \sb_1__0__1_chanx_left_out[16] ,
    \sb_1__0__1_chanx_left_out[17] ,
    \sb_1__0__1_chanx_left_out[18] ,
    \sb_1__0__1_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__0__2_chanx_left_out[0] ,
    \cbx_1__0__2_chanx_left_out[1] ,
    \cbx_1__0__2_chanx_left_out[2] ,
    \cbx_1__0__2_chanx_left_out[3] ,
    \cbx_1__0__2_chanx_left_out[4] ,
    \cbx_1__0__2_chanx_left_out[5] ,
    \cbx_1__0__2_chanx_left_out[6] ,
    \cbx_1__0__2_chanx_left_out[7] ,
    \cbx_1__0__2_chanx_left_out[8] ,
    \cbx_1__0__2_chanx_left_out[9] ,
    \cbx_1__0__2_chanx_left_out[10] ,
    \cbx_1__0__2_chanx_left_out[11] ,
    \cbx_1__0__2_chanx_left_out[12] ,
    \cbx_1__0__2_chanx_left_out[13] ,
    \cbx_1__0__2_chanx_left_out[14] ,
    \cbx_1__0__2_chanx_left_out[15] ,
    \cbx_1__0__2_chanx_left_out[16] ,
    \cbx_1__0__2_chanx_left_out[17] ,
    \cbx_1__0__2_chanx_left_out[18] ,
    \cbx_1__0__2_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__0__1_chanx_right_out[0] ,
    \sb_1__0__1_chanx_right_out[1] ,
    \sb_1__0__1_chanx_right_out[2] ,
    \sb_1__0__1_chanx_right_out[3] ,
    \sb_1__0__1_chanx_right_out[4] ,
    \sb_1__0__1_chanx_right_out[5] ,
    \sb_1__0__1_chanx_right_out[6] ,
    \sb_1__0__1_chanx_right_out[7] ,
    \sb_1__0__1_chanx_right_out[8] ,
    \sb_1__0__1_chanx_right_out[9] ,
    \sb_1__0__1_chanx_right_out[10] ,
    \sb_1__0__1_chanx_right_out[11] ,
    \sb_1__0__1_chanx_right_out[12] ,
    \sb_1__0__1_chanx_right_out[13] ,
    \sb_1__0__1_chanx_right_out[14] ,
    \sb_1__0__1_chanx_right_out[15] ,
    \sb_1__0__1_chanx_right_out[16] ,
    \sb_1__0__1_chanx_right_out[17] ,
    \sb_1__0__1_chanx_right_out[18] ,
    \sb_1__0__1_chanx_right_out[19] }),
    .chany_top_in({\cby_1__1__8_chany_bottom_out[0] ,
    \cby_1__1__8_chany_bottom_out[1] ,
    \cby_1__1__8_chany_bottom_out[2] ,
    \cby_1__1__8_chany_bottom_out[3] ,
    \cby_1__1__8_chany_bottom_out[4] ,
    \cby_1__1__8_chany_bottom_out[5] ,
    \cby_1__1__8_chany_bottom_out[6] ,
    \cby_1__1__8_chany_bottom_out[7] ,
    \cby_1__1__8_chany_bottom_out[8] ,
    \cby_1__1__8_chany_bottom_out[9] ,
    \cby_1__1__8_chany_bottom_out[10] ,
    \cby_1__1__8_chany_bottom_out[11] ,
    \cby_1__1__8_chany_bottom_out[12] ,
    \cby_1__1__8_chany_bottom_out[13] ,
    \cby_1__1__8_chany_bottom_out[14] ,
    \cby_1__1__8_chany_bottom_out[15] ,
    \cby_1__1__8_chany_bottom_out[16] ,
    \cby_1__1__8_chany_bottom_out[17] ,
    \cby_1__1__8_chany_bottom_out[18] ,
    \cby_1__1__8_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__0__1_chany_top_out[0] ,
    \sb_1__0__1_chany_top_out[1] ,
    \sb_1__0__1_chany_top_out[2] ,
    \sb_1__0__1_chany_top_out[3] ,
    \sb_1__0__1_chany_top_out[4] ,
    \sb_1__0__1_chany_top_out[5] ,
    \sb_1__0__1_chany_top_out[6] ,
    \sb_1__0__1_chany_top_out[7] ,
    \sb_1__0__1_chany_top_out[8] ,
    \sb_1__0__1_chany_top_out[9] ,
    \sb_1__0__1_chany_top_out[10] ,
    \sb_1__0__1_chany_top_out[11] ,
    \sb_1__0__1_chany_top_out[12] ,
    \sb_1__0__1_chany_top_out[13] ,
    \sb_1__0__1_chany_top_out[14] ,
    \sb_1__0__1_chany_top_out[15] ,
    \sb_1__0__1_chany_top_out[16] ,
    \sb_1__0__1_chany_top_out[17] ,
    \sb_1__0__1_chany_top_out[18] ,
    \sb_1__0__1_chany_top_out[19] }));
 sb_1__1_ sb_2__1_ (.bottom_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__14_ccff_tail),
    .ccff_tail(sb_1__1__7_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[48] ),
    .right_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__7_chanx_right_out[0] ,
    \cbx_1__1__7_chanx_right_out[1] ,
    \cbx_1__1__7_chanx_right_out[2] ,
    \cbx_1__1__7_chanx_right_out[3] ,
    \cbx_1__1__7_chanx_right_out[4] ,
    \cbx_1__1__7_chanx_right_out[5] ,
    \cbx_1__1__7_chanx_right_out[6] ,
    \cbx_1__1__7_chanx_right_out[7] ,
    \cbx_1__1__7_chanx_right_out[8] ,
    \cbx_1__1__7_chanx_right_out[9] ,
    \cbx_1__1__7_chanx_right_out[10] ,
    \cbx_1__1__7_chanx_right_out[11] ,
    \cbx_1__1__7_chanx_right_out[12] ,
    \cbx_1__1__7_chanx_right_out[13] ,
    \cbx_1__1__7_chanx_right_out[14] ,
    \cbx_1__1__7_chanx_right_out[15] ,
    \cbx_1__1__7_chanx_right_out[16] ,
    \cbx_1__1__7_chanx_right_out[17] ,
    \cbx_1__1__7_chanx_right_out[18] ,
    \cbx_1__1__7_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__7_chanx_left_out[0] ,
    \sb_1__1__7_chanx_left_out[1] ,
    \sb_1__1__7_chanx_left_out[2] ,
    \sb_1__1__7_chanx_left_out[3] ,
    \sb_1__1__7_chanx_left_out[4] ,
    \sb_1__1__7_chanx_left_out[5] ,
    \sb_1__1__7_chanx_left_out[6] ,
    \sb_1__1__7_chanx_left_out[7] ,
    \sb_1__1__7_chanx_left_out[8] ,
    \sb_1__1__7_chanx_left_out[9] ,
    \sb_1__1__7_chanx_left_out[10] ,
    \sb_1__1__7_chanx_left_out[11] ,
    \sb_1__1__7_chanx_left_out[12] ,
    \sb_1__1__7_chanx_left_out[13] ,
    \sb_1__1__7_chanx_left_out[14] ,
    \sb_1__1__7_chanx_left_out[15] ,
    \sb_1__1__7_chanx_left_out[16] ,
    \sb_1__1__7_chanx_left_out[17] ,
    \sb_1__1__7_chanx_left_out[18] ,
    \sb_1__1__7_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__14_chanx_left_out[0] ,
    \cbx_1__1__14_chanx_left_out[1] ,
    \cbx_1__1__14_chanx_left_out[2] ,
    \cbx_1__1__14_chanx_left_out[3] ,
    \cbx_1__1__14_chanx_left_out[4] ,
    \cbx_1__1__14_chanx_left_out[5] ,
    \cbx_1__1__14_chanx_left_out[6] ,
    \cbx_1__1__14_chanx_left_out[7] ,
    \cbx_1__1__14_chanx_left_out[8] ,
    \cbx_1__1__14_chanx_left_out[9] ,
    \cbx_1__1__14_chanx_left_out[10] ,
    \cbx_1__1__14_chanx_left_out[11] ,
    \cbx_1__1__14_chanx_left_out[12] ,
    \cbx_1__1__14_chanx_left_out[13] ,
    \cbx_1__1__14_chanx_left_out[14] ,
    \cbx_1__1__14_chanx_left_out[15] ,
    \cbx_1__1__14_chanx_left_out[16] ,
    \cbx_1__1__14_chanx_left_out[17] ,
    \cbx_1__1__14_chanx_left_out[18] ,
    \cbx_1__1__14_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__7_chanx_right_out[0] ,
    \sb_1__1__7_chanx_right_out[1] ,
    \sb_1__1__7_chanx_right_out[2] ,
    \sb_1__1__7_chanx_right_out[3] ,
    \sb_1__1__7_chanx_right_out[4] ,
    \sb_1__1__7_chanx_right_out[5] ,
    \sb_1__1__7_chanx_right_out[6] ,
    \sb_1__1__7_chanx_right_out[7] ,
    \sb_1__1__7_chanx_right_out[8] ,
    \sb_1__1__7_chanx_right_out[9] ,
    \sb_1__1__7_chanx_right_out[10] ,
    \sb_1__1__7_chanx_right_out[11] ,
    \sb_1__1__7_chanx_right_out[12] ,
    \sb_1__1__7_chanx_right_out[13] ,
    \sb_1__1__7_chanx_right_out[14] ,
    \sb_1__1__7_chanx_right_out[15] ,
    \sb_1__1__7_chanx_right_out[16] ,
    \sb_1__1__7_chanx_right_out[17] ,
    \sb_1__1__7_chanx_right_out[18] ,
    \sb_1__1__7_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__8_chany_top_out[0] ,
    \cby_1__1__8_chany_top_out[1] ,
    \cby_1__1__8_chany_top_out[2] ,
    \cby_1__1__8_chany_top_out[3] ,
    \cby_1__1__8_chany_top_out[4] ,
    \cby_1__1__8_chany_top_out[5] ,
    \cby_1__1__8_chany_top_out[6] ,
    \cby_1__1__8_chany_top_out[7] ,
    \cby_1__1__8_chany_top_out[8] ,
    \cby_1__1__8_chany_top_out[9] ,
    \cby_1__1__8_chany_top_out[10] ,
    \cby_1__1__8_chany_top_out[11] ,
    \cby_1__1__8_chany_top_out[12] ,
    \cby_1__1__8_chany_top_out[13] ,
    \cby_1__1__8_chany_top_out[14] ,
    \cby_1__1__8_chany_top_out[15] ,
    \cby_1__1__8_chany_top_out[16] ,
    \cby_1__1__8_chany_top_out[17] ,
    \cby_1__1__8_chany_top_out[18] ,
    \cby_1__1__8_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__7_chany_bottom_out[0] ,
    \sb_1__1__7_chany_bottom_out[1] ,
    \sb_1__1__7_chany_bottom_out[2] ,
    \sb_1__1__7_chany_bottom_out[3] ,
    \sb_1__1__7_chany_bottom_out[4] ,
    \sb_1__1__7_chany_bottom_out[5] ,
    \sb_1__1__7_chany_bottom_out[6] ,
    \sb_1__1__7_chany_bottom_out[7] ,
    \sb_1__1__7_chany_bottom_out[8] ,
    \sb_1__1__7_chany_bottom_out[9] ,
    \sb_1__1__7_chany_bottom_out[10] ,
    \sb_1__1__7_chany_bottom_out[11] ,
    \sb_1__1__7_chany_bottom_out[12] ,
    \sb_1__1__7_chany_bottom_out[13] ,
    \sb_1__1__7_chany_bottom_out[14] ,
    \sb_1__1__7_chany_bottom_out[15] ,
    \sb_1__1__7_chany_bottom_out[16] ,
    \sb_1__1__7_chany_bottom_out[17] ,
    \sb_1__1__7_chany_bottom_out[18] ,
    \sb_1__1__7_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__9_chany_bottom_out[0] ,
    \cby_1__1__9_chany_bottom_out[1] ,
    \cby_1__1__9_chany_bottom_out[2] ,
    \cby_1__1__9_chany_bottom_out[3] ,
    \cby_1__1__9_chany_bottom_out[4] ,
    \cby_1__1__9_chany_bottom_out[5] ,
    \cby_1__1__9_chany_bottom_out[6] ,
    \cby_1__1__9_chany_bottom_out[7] ,
    \cby_1__1__9_chany_bottom_out[8] ,
    \cby_1__1__9_chany_bottom_out[9] ,
    \cby_1__1__9_chany_bottom_out[10] ,
    \cby_1__1__9_chany_bottom_out[11] ,
    \cby_1__1__9_chany_bottom_out[12] ,
    \cby_1__1__9_chany_bottom_out[13] ,
    \cby_1__1__9_chany_bottom_out[14] ,
    \cby_1__1__9_chany_bottom_out[15] ,
    \cby_1__1__9_chany_bottom_out[16] ,
    \cby_1__1__9_chany_bottom_out[17] ,
    \cby_1__1__9_chany_bottom_out[18] ,
    \cby_1__1__9_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__7_chany_top_out[0] ,
    \sb_1__1__7_chany_top_out[1] ,
    \sb_1__1__7_chany_top_out[2] ,
    \sb_1__1__7_chany_top_out[3] ,
    \sb_1__1__7_chany_top_out[4] ,
    \sb_1__1__7_chany_top_out[5] ,
    \sb_1__1__7_chany_top_out[6] ,
    \sb_1__1__7_chany_top_out[7] ,
    \sb_1__1__7_chany_top_out[8] ,
    \sb_1__1__7_chany_top_out[9] ,
    \sb_1__1__7_chany_top_out[10] ,
    \sb_1__1__7_chany_top_out[11] ,
    \sb_1__1__7_chany_top_out[12] ,
    \sb_1__1__7_chany_top_out[13] ,
    \sb_1__1__7_chany_top_out[14] ,
    \sb_1__1__7_chany_top_out[15] ,
    \sb_1__1__7_chany_top_out[16] ,
    \sb_1__1__7_chany_top_out[17] ,
    \sb_1__1__7_chany_top_out[18] ,
    \sb_1__1__7_chany_top_out[19] }));
 sb_1__1_ sb_2__2_ (.bottom_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__15_ccff_tail),
    .ccff_tail(sb_1__1__8_ccff_tail),
    .clk_2_E_out(\clk_2_wires[1] ),
    .clk_2_N_in(\clk_3_wires[17] ),
    .clk_2_W_out(\clk_2_wires[3] ),
    .left_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[51] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[1] ),
    .prog_clk_2_N_in(\prog_clk_3_wires[17] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[3] ),
    .right_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__8_chanx_right_out[0] ,
    \cbx_1__1__8_chanx_right_out[1] ,
    \cbx_1__1__8_chanx_right_out[2] ,
    \cbx_1__1__8_chanx_right_out[3] ,
    \cbx_1__1__8_chanx_right_out[4] ,
    \cbx_1__1__8_chanx_right_out[5] ,
    \cbx_1__1__8_chanx_right_out[6] ,
    \cbx_1__1__8_chanx_right_out[7] ,
    \cbx_1__1__8_chanx_right_out[8] ,
    \cbx_1__1__8_chanx_right_out[9] ,
    \cbx_1__1__8_chanx_right_out[10] ,
    \cbx_1__1__8_chanx_right_out[11] ,
    \cbx_1__1__8_chanx_right_out[12] ,
    \cbx_1__1__8_chanx_right_out[13] ,
    \cbx_1__1__8_chanx_right_out[14] ,
    \cbx_1__1__8_chanx_right_out[15] ,
    \cbx_1__1__8_chanx_right_out[16] ,
    \cbx_1__1__8_chanx_right_out[17] ,
    \cbx_1__1__8_chanx_right_out[18] ,
    \cbx_1__1__8_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__8_chanx_left_out[0] ,
    \sb_1__1__8_chanx_left_out[1] ,
    \sb_1__1__8_chanx_left_out[2] ,
    \sb_1__1__8_chanx_left_out[3] ,
    \sb_1__1__8_chanx_left_out[4] ,
    \sb_1__1__8_chanx_left_out[5] ,
    \sb_1__1__8_chanx_left_out[6] ,
    \sb_1__1__8_chanx_left_out[7] ,
    \sb_1__1__8_chanx_left_out[8] ,
    \sb_1__1__8_chanx_left_out[9] ,
    \sb_1__1__8_chanx_left_out[10] ,
    \sb_1__1__8_chanx_left_out[11] ,
    \sb_1__1__8_chanx_left_out[12] ,
    \sb_1__1__8_chanx_left_out[13] ,
    \sb_1__1__8_chanx_left_out[14] ,
    \sb_1__1__8_chanx_left_out[15] ,
    \sb_1__1__8_chanx_left_out[16] ,
    \sb_1__1__8_chanx_left_out[17] ,
    \sb_1__1__8_chanx_left_out[18] ,
    \sb_1__1__8_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__15_chanx_left_out[0] ,
    \cbx_1__1__15_chanx_left_out[1] ,
    \cbx_1__1__15_chanx_left_out[2] ,
    \cbx_1__1__15_chanx_left_out[3] ,
    \cbx_1__1__15_chanx_left_out[4] ,
    \cbx_1__1__15_chanx_left_out[5] ,
    \cbx_1__1__15_chanx_left_out[6] ,
    \cbx_1__1__15_chanx_left_out[7] ,
    \cbx_1__1__15_chanx_left_out[8] ,
    \cbx_1__1__15_chanx_left_out[9] ,
    \cbx_1__1__15_chanx_left_out[10] ,
    \cbx_1__1__15_chanx_left_out[11] ,
    \cbx_1__1__15_chanx_left_out[12] ,
    \cbx_1__1__15_chanx_left_out[13] ,
    \cbx_1__1__15_chanx_left_out[14] ,
    \cbx_1__1__15_chanx_left_out[15] ,
    \cbx_1__1__15_chanx_left_out[16] ,
    \cbx_1__1__15_chanx_left_out[17] ,
    \cbx_1__1__15_chanx_left_out[18] ,
    \cbx_1__1__15_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__8_chanx_right_out[0] ,
    \sb_1__1__8_chanx_right_out[1] ,
    \sb_1__1__8_chanx_right_out[2] ,
    \sb_1__1__8_chanx_right_out[3] ,
    \sb_1__1__8_chanx_right_out[4] ,
    \sb_1__1__8_chanx_right_out[5] ,
    \sb_1__1__8_chanx_right_out[6] ,
    \sb_1__1__8_chanx_right_out[7] ,
    \sb_1__1__8_chanx_right_out[8] ,
    \sb_1__1__8_chanx_right_out[9] ,
    \sb_1__1__8_chanx_right_out[10] ,
    \sb_1__1__8_chanx_right_out[11] ,
    \sb_1__1__8_chanx_right_out[12] ,
    \sb_1__1__8_chanx_right_out[13] ,
    \sb_1__1__8_chanx_right_out[14] ,
    \sb_1__1__8_chanx_right_out[15] ,
    \sb_1__1__8_chanx_right_out[16] ,
    \sb_1__1__8_chanx_right_out[17] ,
    \sb_1__1__8_chanx_right_out[18] ,
    \sb_1__1__8_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__9_chany_top_out[0] ,
    \cby_1__1__9_chany_top_out[1] ,
    \cby_1__1__9_chany_top_out[2] ,
    \cby_1__1__9_chany_top_out[3] ,
    \cby_1__1__9_chany_top_out[4] ,
    \cby_1__1__9_chany_top_out[5] ,
    \cby_1__1__9_chany_top_out[6] ,
    \cby_1__1__9_chany_top_out[7] ,
    \cby_1__1__9_chany_top_out[8] ,
    \cby_1__1__9_chany_top_out[9] ,
    \cby_1__1__9_chany_top_out[10] ,
    \cby_1__1__9_chany_top_out[11] ,
    \cby_1__1__9_chany_top_out[12] ,
    \cby_1__1__9_chany_top_out[13] ,
    \cby_1__1__9_chany_top_out[14] ,
    \cby_1__1__9_chany_top_out[15] ,
    \cby_1__1__9_chany_top_out[16] ,
    \cby_1__1__9_chany_top_out[17] ,
    \cby_1__1__9_chany_top_out[18] ,
    \cby_1__1__9_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__8_chany_bottom_out[0] ,
    \sb_1__1__8_chany_bottom_out[1] ,
    \sb_1__1__8_chany_bottom_out[2] ,
    \sb_1__1__8_chany_bottom_out[3] ,
    \sb_1__1__8_chany_bottom_out[4] ,
    \sb_1__1__8_chany_bottom_out[5] ,
    \sb_1__1__8_chany_bottom_out[6] ,
    \sb_1__1__8_chany_bottom_out[7] ,
    \sb_1__1__8_chany_bottom_out[8] ,
    \sb_1__1__8_chany_bottom_out[9] ,
    \sb_1__1__8_chany_bottom_out[10] ,
    \sb_1__1__8_chany_bottom_out[11] ,
    \sb_1__1__8_chany_bottom_out[12] ,
    \sb_1__1__8_chany_bottom_out[13] ,
    \sb_1__1__8_chany_bottom_out[14] ,
    \sb_1__1__8_chany_bottom_out[15] ,
    \sb_1__1__8_chany_bottom_out[16] ,
    \sb_1__1__8_chany_bottom_out[17] ,
    \sb_1__1__8_chany_bottom_out[18] ,
    \sb_1__1__8_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__10_chany_bottom_out[0] ,
    \cby_1__1__10_chany_bottom_out[1] ,
    \cby_1__1__10_chany_bottom_out[2] ,
    \cby_1__1__10_chany_bottom_out[3] ,
    \cby_1__1__10_chany_bottom_out[4] ,
    \cby_1__1__10_chany_bottom_out[5] ,
    \cby_1__1__10_chany_bottom_out[6] ,
    \cby_1__1__10_chany_bottom_out[7] ,
    \cby_1__1__10_chany_bottom_out[8] ,
    \cby_1__1__10_chany_bottom_out[9] ,
    \cby_1__1__10_chany_bottom_out[10] ,
    \cby_1__1__10_chany_bottom_out[11] ,
    \cby_1__1__10_chany_bottom_out[12] ,
    \cby_1__1__10_chany_bottom_out[13] ,
    \cby_1__1__10_chany_bottom_out[14] ,
    \cby_1__1__10_chany_bottom_out[15] ,
    \cby_1__1__10_chany_bottom_out[16] ,
    \cby_1__1__10_chany_bottom_out[17] ,
    \cby_1__1__10_chany_bottom_out[18] ,
    \cby_1__1__10_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__8_chany_top_out[0] ,
    \sb_1__1__8_chany_top_out[1] ,
    \sb_1__1__8_chany_top_out[2] ,
    \sb_1__1__8_chany_top_out[3] ,
    \sb_1__1__8_chany_top_out[4] ,
    \sb_1__1__8_chany_top_out[5] ,
    \sb_1__1__8_chany_top_out[6] ,
    \sb_1__1__8_chany_top_out[7] ,
    \sb_1__1__8_chany_top_out[8] ,
    \sb_1__1__8_chany_top_out[9] ,
    \sb_1__1__8_chany_top_out[10] ,
    \sb_1__1__8_chany_top_out[11] ,
    \sb_1__1__8_chany_top_out[12] ,
    \sb_1__1__8_chany_top_out[13] ,
    \sb_1__1__8_chany_top_out[14] ,
    \sb_1__1__8_chany_top_out[15] ,
    \sb_1__1__8_chany_top_out[16] ,
    \sb_1__1__8_chany_top_out[17] ,
    \sb_1__1__8_chany_top_out[18] ,
    \sb_1__1__8_chany_top_out[19] }));
 sb_1__1_ sb_2__3_ (.bottom_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__16_ccff_tail),
    .ccff_tail(sb_1__1__9_ccff_tail),
    .clk_3_N_in(\clk_3_wires[13] ),
    .clk_3_S_out(\clk_3_wires[16] ),
    .left_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[54] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[13] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[16] ),
    .right_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__9_chanx_right_out[0] ,
    \cbx_1__1__9_chanx_right_out[1] ,
    \cbx_1__1__9_chanx_right_out[2] ,
    \cbx_1__1__9_chanx_right_out[3] ,
    \cbx_1__1__9_chanx_right_out[4] ,
    \cbx_1__1__9_chanx_right_out[5] ,
    \cbx_1__1__9_chanx_right_out[6] ,
    \cbx_1__1__9_chanx_right_out[7] ,
    \cbx_1__1__9_chanx_right_out[8] ,
    \cbx_1__1__9_chanx_right_out[9] ,
    \cbx_1__1__9_chanx_right_out[10] ,
    \cbx_1__1__9_chanx_right_out[11] ,
    \cbx_1__1__9_chanx_right_out[12] ,
    \cbx_1__1__9_chanx_right_out[13] ,
    \cbx_1__1__9_chanx_right_out[14] ,
    \cbx_1__1__9_chanx_right_out[15] ,
    \cbx_1__1__9_chanx_right_out[16] ,
    \cbx_1__1__9_chanx_right_out[17] ,
    \cbx_1__1__9_chanx_right_out[18] ,
    \cbx_1__1__9_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__9_chanx_left_out[0] ,
    \sb_1__1__9_chanx_left_out[1] ,
    \sb_1__1__9_chanx_left_out[2] ,
    \sb_1__1__9_chanx_left_out[3] ,
    \sb_1__1__9_chanx_left_out[4] ,
    \sb_1__1__9_chanx_left_out[5] ,
    \sb_1__1__9_chanx_left_out[6] ,
    \sb_1__1__9_chanx_left_out[7] ,
    \sb_1__1__9_chanx_left_out[8] ,
    \sb_1__1__9_chanx_left_out[9] ,
    \sb_1__1__9_chanx_left_out[10] ,
    \sb_1__1__9_chanx_left_out[11] ,
    \sb_1__1__9_chanx_left_out[12] ,
    \sb_1__1__9_chanx_left_out[13] ,
    \sb_1__1__9_chanx_left_out[14] ,
    \sb_1__1__9_chanx_left_out[15] ,
    \sb_1__1__9_chanx_left_out[16] ,
    \sb_1__1__9_chanx_left_out[17] ,
    \sb_1__1__9_chanx_left_out[18] ,
    \sb_1__1__9_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__16_chanx_left_out[0] ,
    \cbx_1__1__16_chanx_left_out[1] ,
    \cbx_1__1__16_chanx_left_out[2] ,
    \cbx_1__1__16_chanx_left_out[3] ,
    \cbx_1__1__16_chanx_left_out[4] ,
    \cbx_1__1__16_chanx_left_out[5] ,
    \cbx_1__1__16_chanx_left_out[6] ,
    \cbx_1__1__16_chanx_left_out[7] ,
    \cbx_1__1__16_chanx_left_out[8] ,
    \cbx_1__1__16_chanx_left_out[9] ,
    \cbx_1__1__16_chanx_left_out[10] ,
    \cbx_1__1__16_chanx_left_out[11] ,
    \cbx_1__1__16_chanx_left_out[12] ,
    \cbx_1__1__16_chanx_left_out[13] ,
    \cbx_1__1__16_chanx_left_out[14] ,
    \cbx_1__1__16_chanx_left_out[15] ,
    \cbx_1__1__16_chanx_left_out[16] ,
    \cbx_1__1__16_chanx_left_out[17] ,
    \cbx_1__1__16_chanx_left_out[18] ,
    \cbx_1__1__16_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__9_chanx_right_out[0] ,
    \sb_1__1__9_chanx_right_out[1] ,
    \sb_1__1__9_chanx_right_out[2] ,
    \sb_1__1__9_chanx_right_out[3] ,
    \sb_1__1__9_chanx_right_out[4] ,
    \sb_1__1__9_chanx_right_out[5] ,
    \sb_1__1__9_chanx_right_out[6] ,
    \sb_1__1__9_chanx_right_out[7] ,
    \sb_1__1__9_chanx_right_out[8] ,
    \sb_1__1__9_chanx_right_out[9] ,
    \sb_1__1__9_chanx_right_out[10] ,
    \sb_1__1__9_chanx_right_out[11] ,
    \sb_1__1__9_chanx_right_out[12] ,
    \sb_1__1__9_chanx_right_out[13] ,
    \sb_1__1__9_chanx_right_out[14] ,
    \sb_1__1__9_chanx_right_out[15] ,
    \sb_1__1__9_chanx_right_out[16] ,
    \sb_1__1__9_chanx_right_out[17] ,
    \sb_1__1__9_chanx_right_out[18] ,
    \sb_1__1__9_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__10_chany_top_out[0] ,
    \cby_1__1__10_chany_top_out[1] ,
    \cby_1__1__10_chany_top_out[2] ,
    \cby_1__1__10_chany_top_out[3] ,
    \cby_1__1__10_chany_top_out[4] ,
    \cby_1__1__10_chany_top_out[5] ,
    \cby_1__1__10_chany_top_out[6] ,
    \cby_1__1__10_chany_top_out[7] ,
    \cby_1__1__10_chany_top_out[8] ,
    \cby_1__1__10_chany_top_out[9] ,
    \cby_1__1__10_chany_top_out[10] ,
    \cby_1__1__10_chany_top_out[11] ,
    \cby_1__1__10_chany_top_out[12] ,
    \cby_1__1__10_chany_top_out[13] ,
    \cby_1__1__10_chany_top_out[14] ,
    \cby_1__1__10_chany_top_out[15] ,
    \cby_1__1__10_chany_top_out[16] ,
    \cby_1__1__10_chany_top_out[17] ,
    \cby_1__1__10_chany_top_out[18] ,
    \cby_1__1__10_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__9_chany_bottom_out[0] ,
    \sb_1__1__9_chany_bottom_out[1] ,
    \sb_1__1__9_chany_bottom_out[2] ,
    \sb_1__1__9_chany_bottom_out[3] ,
    \sb_1__1__9_chany_bottom_out[4] ,
    \sb_1__1__9_chany_bottom_out[5] ,
    \sb_1__1__9_chany_bottom_out[6] ,
    \sb_1__1__9_chany_bottom_out[7] ,
    \sb_1__1__9_chany_bottom_out[8] ,
    \sb_1__1__9_chany_bottom_out[9] ,
    \sb_1__1__9_chany_bottom_out[10] ,
    \sb_1__1__9_chany_bottom_out[11] ,
    \sb_1__1__9_chany_bottom_out[12] ,
    \sb_1__1__9_chany_bottom_out[13] ,
    \sb_1__1__9_chany_bottom_out[14] ,
    \sb_1__1__9_chany_bottom_out[15] ,
    \sb_1__1__9_chany_bottom_out[16] ,
    \sb_1__1__9_chany_bottom_out[17] ,
    \sb_1__1__9_chany_bottom_out[18] ,
    \sb_1__1__9_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__11_chany_bottom_out[0] ,
    \cby_1__1__11_chany_bottom_out[1] ,
    \cby_1__1__11_chany_bottom_out[2] ,
    \cby_1__1__11_chany_bottom_out[3] ,
    \cby_1__1__11_chany_bottom_out[4] ,
    \cby_1__1__11_chany_bottom_out[5] ,
    \cby_1__1__11_chany_bottom_out[6] ,
    \cby_1__1__11_chany_bottom_out[7] ,
    \cby_1__1__11_chany_bottom_out[8] ,
    \cby_1__1__11_chany_bottom_out[9] ,
    \cby_1__1__11_chany_bottom_out[10] ,
    \cby_1__1__11_chany_bottom_out[11] ,
    \cby_1__1__11_chany_bottom_out[12] ,
    \cby_1__1__11_chany_bottom_out[13] ,
    \cby_1__1__11_chany_bottom_out[14] ,
    \cby_1__1__11_chany_bottom_out[15] ,
    \cby_1__1__11_chany_bottom_out[16] ,
    \cby_1__1__11_chany_bottom_out[17] ,
    \cby_1__1__11_chany_bottom_out[18] ,
    \cby_1__1__11_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__9_chany_top_out[0] ,
    \sb_1__1__9_chany_top_out[1] ,
    \sb_1__1__9_chany_top_out[2] ,
    \sb_1__1__9_chany_top_out[3] ,
    \sb_1__1__9_chany_top_out[4] ,
    \sb_1__1__9_chany_top_out[5] ,
    \sb_1__1__9_chany_top_out[6] ,
    \sb_1__1__9_chany_top_out[7] ,
    \sb_1__1__9_chany_top_out[8] ,
    \sb_1__1__9_chany_top_out[9] ,
    \sb_1__1__9_chany_top_out[10] ,
    \sb_1__1__9_chany_top_out[11] ,
    \sb_1__1__9_chany_top_out[12] ,
    \sb_1__1__9_chany_top_out[13] ,
    \sb_1__1__9_chany_top_out[14] ,
    \sb_1__1__9_chany_top_out[15] ,
    \sb_1__1__9_chany_top_out[16] ,
    \sb_1__1__9_chany_top_out[17] ,
    \sb_1__1__9_chany_top_out[18] ,
    \sb_1__1__9_chany_top_out[19] }));
 sb_1__1_ sb_2__4_ (.bottom_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__17_ccff_tail),
    .ccff_tail(sb_1__1__10_ccff_tail),
    .clk_3_N_in(\clk_3_wires[9] ),
    .clk_3_N_out(\clk_3_wires[10] ),
    .clk_3_S_out(\clk_3_wires[12] ),
    .left_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[57] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[9] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[10] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[12] ),
    .right_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__10_chanx_right_out[0] ,
    \cbx_1__1__10_chanx_right_out[1] ,
    \cbx_1__1__10_chanx_right_out[2] ,
    \cbx_1__1__10_chanx_right_out[3] ,
    \cbx_1__1__10_chanx_right_out[4] ,
    \cbx_1__1__10_chanx_right_out[5] ,
    \cbx_1__1__10_chanx_right_out[6] ,
    \cbx_1__1__10_chanx_right_out[7] ,
    \cbx_1__1__10_chanx_right_out[8] ,
    \cbx_1__1__10_chanx_right_out[9] ,
    \cbx_1__1__10_chanx_right_out[10] ,
    \cbx_1__1__10_chanx_right_out[11] ,
    \cbx_1__1__10_chanx_right_out[12] ,
    \cbx_1__1__10_chanx_right_out[13] ,
    \cbx_1__1__10_chanx_right_out[14] ,
    \cbx_1__1__10_chanx_right_out[15] ,
    \cbx_1__1__10_chanx_right_out[16] ,
    \cbx_1__1__10_chanx_right_out[17] ,
    \cbx_1__1__10_chanx_right_out[18] ,
    \cbx_1__1__10_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__10_chanx_left_out[0] ,
    \sb_1__1__10_chanx_left_out[1] ,
    \sb_1__1__10_chanx_left_out[2] ,
    \sb_1__1__10_chanx_left_out[3] ,
    \sb_1__1__10_chanx_left_out[4] ,
    \sb_1__1__10_chanx_left_out[5] ,
    \sb_1__1__10_chanx_left_out[6] ,
    \sb_1__1__10_chanx_left_out[7] ,
    \sb_1__1__10_chanx_left_out[8] ,
    \sb_1__1__10_chanx_left_out[9] ,
    \sb_1__1__10_chanx_left_out[10] ,
    \sb_1__1__10_chanx_left_out[11] ,
    \sb_1__1__10_chanx_left_out[12] ,
    \sb_1__1__10_chanx_left_out[13] ,
    \sb_1__1__10_chanx_left_out[14] ,
    \sb_1__1__10_chanx_left_out[15] ,
    \sb_1__1__10_chanx_left_out[16] ,
    \sb_1__1__10_chanx_left_out[17] ,
    \sb_1__1__10_chanx_left_out[18] ,
    \sb_1__1__10_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__17_chanx_left_out[0] ,
    \cbx_1__1__17_chanx_left_out[1] ,
    \cbx_1__1__17_chanx_left_out[2] ,
    \cbx_1__1__17_chanx_left_out[3] ,
    \cbx_1__1__17_chanx_left_out[4] ,
    \cbx_1__1__17_chanx_left_out[5] ,
    \cbx_1__1__17_chanx_left_out[6] ,
    \cbx_1__1__17_chanx_left_out[7] ,
    \cbx_1__1__17_chanx_left_out[8] ,
    \cbx_1__1__17_chanx_left_out[9] ,
    \cbx_1__1__17_chanx_left_out[10] ,
    \cbx_1__1__17_chanx_left_out[11] ,
    \cbx_1__1__17_chanx_left_out[12] ,
    \cbx_1__1__17_chanx_left_out[13] ,
    \cbx_1__1__17_chanx_left_out[14] ,
    \cbx_1__1__17_chanx_left_out[15] ,
    \cbx_1__1__17_chanx_left_out[16] ,
    \cbx_1__1__17_chanx_left_out[17] ,
    \cbx_1__1__17_chanx_left_out[18] ,
    \cbx_1__1__17_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__10_chanx_right_out[0] ,
    \sb_1__1__10_chanx_right_out[1] ,
    \sb_1__1__10_chanx_right_out[2] ,
    \sb_1__1__10_chanx_right_out[3] ,
    \sb_1__1__10_chanx_right_out[4] ,
    \sb_1__1__10_chanx_right_out[5] ,
    \sb_1__1__10_chanx_right_out[6] ,
    \sb_1__1__10_chanx_right_out[7] ,
    \sb_1__1__10_chanx_right_out[8] ,
    \sb_1__1__10_chanx_right_out[9] ,
    \sb_1__1__10_chanx_right_out[10] ,
    \sb_1__1__10_chanx_right_out[11] ,
    \sb_1__1__10_chanx_right_out[12] ,
    \sb_1__1__10_chanx_right_out[13] ,
    \sb_1__1__10_chanx_right_out[14] ,
    \sb_1__1__10_chanx_right_out[15] ,
    \sb_1__1__10_chanx_right_out[16] ,
    \sb_1__1__10_chanx_right_out[17] ,
    \sb_1__1__10_chanx_right_out[18] ,
    \sb_1__1__10_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__11_chany_top_out[0] ,
    \cby_1__1__11_chany_top_out[1] ,
    \cby_1__1__11_chany_top_out[2] ,
    \cby_1__1__11_chany_top_out[3] ,
    \cby_1__1__11_chany_top_out[4] ,
    \cby_1__1__11_chany_top_out[5] ,
    \cby_1__1__11_chany_top_out[6] ,
    \cby_1__1__11_chany_top_out[7] ,
    \cby_1__1__11_chany_top_out[8] ,
    \cby_1__1__11_chany_top_out[9] ,
    \cby_1__1__11_chany_top_out[10] ,
    \cby_1__1__11_chany_top_out[11] ,
    \cby_1__1__11_chany_top_out[12] ,
    \cby_1__1__11_chany_top_out[13] ,
    \cby_1__1__11_chany_top_out[14] ,
    \cby_1__1__11_chany_top_out[15] ,
    \cby_1__1__11_chany_top_out[16] ,
    \cby_1__1__11_chany_top_out[17] ,
    \cby_1__1__11_chany_top_out[18] ,
    \cby_1__1__11_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__10_chany_bottom_out[0] ,
    \sb_1__1__10_chany_bottom_out[1] ,
    \sb_1__1__10_chany_bottom_out[2] ,
    \sb_1__1__10_chany_bottom_out[3] ,
    \sb_1__1__10_chany_bottom_out[4] ,
    \sb_1__1__10_chany_bottom_out[5] ,
    \sb_1__1__10_chany_bottom_out[6] ,
    \sb_1__1__10_chany_bottom_out[7] ,
    \sb_1__1__10_chany_bottom_out[8] ,
    \sb_1__1__10_chany_bottom_out[9] ,
    \sb_1__1__10_chany_bottom_out[10] ,
    \sb_1__1__10_chany_bottom_out[11] ,
    \sb_1__1__10_chany_bottom_out[12] ,
    \sb_1__1__10_chany_bottom_out[13] ,
    \sb_1__1__10_chany_bottom_out[14] ,
    \sb_1__1__10_chany_bottom_out[15] ,
    \sb_1__1__10_chany_bottom_out[16] ,
    \sb_1__1__10_chany_bottom_out[17] ,
    \sb_1__1__10_chany_bottom_out[18] ,
    \sb_1__1__10_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__12_chany_bottom_out[0] ,
    \cby_1__1__12_chany_bottom_out[1] ,
    \cby_1__1__12_chany_bottom_out[2] ,
    \cby_1__1__12_chany_bottom_out[3] ,
    \cby_1__1__12_chany_bottom_out[4] ,
    \cby_1__1__12_chany_bottom_out[5] ,
    \cby_1__1__12_chany_bottom_out[6] ,
    \cby_1__1__12_chany_bottom_out[7] ,
    \cby_1__1__12_chany_bottom_out[8] ,
    \cby_1__1__12_chany_bottom_out[9] ,
    \cby_1__1__12_chany_bottom_out[10] ,
    \cby_1__1__12_chany_bottom_out[11] ,
    \cby_1__1__12_chany_bottom_out[12] ,
    \cby_1__1__12_chany_bottom_out[13] ,
    \cby_1__1__12_chany_bottom_out[14] ,
    \cby_1__1__12_chany_bottom_out[15] ,
    \cby_1__1__12_chany_bottom_out[16] ,
    \cby_1__1__12_chany_bottom_out[17] ,
    \cby_1__1__12_chany_bottom_out[18] ,
    \cby_1__1__12_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__10_chany_top_out[0] ,
    \sb_1__1__10_chany_top_out[1] ,
    \sb_1__1__10_chany_top_out[2] ,
    \sb_1__1__10_chany_top_out[3] ,
    \sb_1__1__10_chany_top_out[4] ,
    \sb_1__1__10_chany_top_out[5] ,
    \sb_1__1__10_chany_top_out[6] ,
    \sb_1__1__10_chany_top_out[7] ,
    \sb_1__1__10_chany_top_out[8] ,
    \sb_1__1__10_chany_top_out[9] ,
    \sb_1__1__10_chany_top_out[10] ,
    \sb_1__1__10_chany_top_out[11] ,
    \sb_1__1__10_chany_top_out[12] ,
    \sb_1__1__10_chany_top_out[13] ,
    \sb_1__1__10_chany_top_out[14] ,
    \sb_1__1__10_chany_top_out[15] ,
    \sb_1__1__10_chany_top_out[16] ,
    \sb_1__1__10_chany_top_out[17] ,
    \sb_1__1__10_chany_top_out[18] ,
    \sb_1__1__10_chany_top_out[19] }));
 sb_1__1_ sb_2__5_ (.bottom_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__18_ccff_tail),
    .ccff_tail(sb_1__1__11_ccff_tail),
    .clk_3_N_in(\clk_3_wires[11] ),
    .clk_3_N_out(\clk_3_wires[14] ),
    .left_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[60] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[11] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[14] ),
    .right_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__11_chanx_right_out[0] ,
    \cbx_1__1__11_chanx_right_out[1] ,
    \cbx_1__1__11_chanx_right_out[2] ,
    \cbx_1__1__11_chanx_right_out[3] ,
    \cbx_1__1__11_chanx_right_out[4] ,
    \cbx_1__1__11_chanx_right_out[5] ,
    \cbx_1__1__11_chanx_right_out[6] ,
    \cbx_1__1__11_chanx_right_out[7] ,
    \cbx_1__1__11_chanx_right_out[8] ,
    \cbx_1__1__11_chanx_right_out[9] ,
    \cbx_1__1__11_chanx_right_out[10] ,
    \cbx_1__1__11_chanx_right_out[11] ,
    \cbx_1__1__11_chanx_right_out[12] ,
    \cbx_1__1__11_chanx_right_out[13] ,
    \cbx_1__1__11_chanx_right_out[14] ,
    \cbx_1__1__11_chanx_right_out[15] ,
    \cbx_1__1__11_chanx_right_out[16] ,
    \cbx_1__1__11_chanx_right_out[17] ,
    \cbx_1__1__11_chanx_right_out[18] ,
    \cbx_1__1__11_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__11_chanx_left_out[0] ,
    \sb_1__1__11_chanx_left_out[1] ,
    \sb_1__1__11_chanx_left_out[2] ,
    \sb_1__1__11_chanx_left_out[3] ,
    \sb_1__1__11_chanx_left_out[4] ,
    \sb_1__1__11_chanx_left_out[5] ,
    \sb_1__1__11_chanx_left_out[6] ,
    \sb_1__1__11_chanx_left_out[7] ,
    \sb_1__1__11_chanx_left_out[8] ,
    \sb_1__1__11_chanx_left_out[9] ,
    \sb_1__1__11_chanx_left_out[10] ,
    \sb_1__1__11_chanx_left_out[11] ,
    \sb_1__1__11_chanx_left_out[12] ,
    \sb_1__1__11_chanx_left_out[13] ,
    \sb_1__1__11_chanx_left_out[14] ,
    \sb_1__1__11_chanx_left_out[15] ,
    \sb_1__1__11_chanx_left_out[16] ,
    \sb_1__1__11_chanx_left_out[17] ,
    \sb_1__1__11_chanx_left_out[18] ,
    \sb_1__1__11_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__18_chanx_left_out[0] ,
    \cbx_1__1__18_chanx_left_out[1] ,
    \cbx_1__1__18_chanx_left_out[2] ,
    \cbx_1__1__18_chanx_left_out[3] ,
    \cbx_1__1__18_chanx_left_out[4] ,
    \cbx_1__1__18_chanx_left_out[5] ,
    \cbx_1__1__18_chanx_left_out[6] ,
    \cbx_1__1__18_chanx_left_out[7] ,
    \cbx_1__1__18_chanx_left_out[8] ,
    \cbx_1__1__18_chanx_left_out[9] ,
    \cbx_1__1__18_chanx_left_out[10] ,
    \cbx_1__1__18_chanx_left_out[11] ,
    \cbx_1__1__18_chanx_left_out[12] ,
    \cbx_1__1__18_chanx_left_out[13] ,
    \cbx_1__1__18_chanx_left_out[14] ,
    \cbx_1__1__18_chanx_left_out[15] ,
    \cbx_1__1__18_chanx_left_out[16] ,
    \cbx_1__1__18_chanx_left_out[17] ,
    \cbx_1__1__18_chanx_left_out[18] ,
    \cbx_1__1__18_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__11_chanx_right_out[0] ,
    \sb_1__1__11_chanx_right_out[1] ,
    \sb_1__1__11_chanx_right_out[2] ,
    \sb_1__1__11_chanx_right_out[3] ,
    \sb_1__1__11_chanx_right_out[4] ,
    \sb_1__1__11_chanx_right_out[5] ,
    \sb_1__1__11_chanx_right_out[6] ,
    \sb_1__1__11_chanx_right_out[7] ,
    \sb_1__1__11_chanx_right_out[8] ,
    \sb_1__1__11_chanx_right_out[9] ,
    \sb_1__1__11_chanx_right_out[10] ,
    \sb_1__1__11_chanx_right_out[11] ,
    \sb_1__1__11_chanx_right_out[12] ,
    \sb_1__1__11_chanx_right_out[13] ,
    \sb_1__1__11_chanx_right_out[14] ,
    \sb_1__1__11_chanx_right_out[15] ,
    \sb_1__1__11_chanx_right_out[16] ,
    \sb_1__1__11_chanx_right_out[17] ,
    \sb_1__1__11_chanx_right_out[18] ,
    \sb_1__1__11_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__12_chany_top_out[0] ,
    \cby_1__1__12_chany_top_out[1] ,
    \cby_1__1__12_chany_top_out[2] ,
    \cby_1__1__12_chany_top_out[3] ,
    \cby_1__1__12_chany_top_out[4] ,
    \cby_1__1__12_chany_top_out[5] ,
    \cby_1__1__12_chany_top_out[6] ,
    \cby_1__1__12_chany_top_out[7] ,
    \cby_1__1__12_chany_top_out[8] ,
    \cby_1__1__12_chany_top_out[9] ,
    \cby_1__1__12_chany_top_out[10] ,
    \cby_1__1__12_chany_top_out[11] ,
    \cby_1__1__12_chany_top_out[12] ,
    \cby_1__1__12_chany_top_out[13] ,
    \cby_1__1__12_chany_top_out[14] ,
    \cby_1__1__12_chany_top_out[15] ,
    \cby_1__1__12_chany_top_out[16] ,
    \cby_1__1__12_chany_top_out[17] ,
    \cby_1__1__12_chany_top_out[18] ,
    \cby_1__1__12_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__11_chany_bottom_out[0] ,
    \sb_1__1__11_chany_bottom_out[1] ,
    \sb_1__1__11_chany_bottom_out[2] ,
    \sb_1__1__11_chany_bottom_out[3] ,
    \sb_1__1__11_chany_bottom_out[4] ,
    \sb_1__1__11_chany_bottom_out[5] ,
    \sb_1__1__11_chany_bottom_out[6] ,
    \sb_1__1__11_chany_bottom_out[7] ,
    \sb_1__1__11_chany_bottom_out[8] ,
    \sb_1__1__11_chany_bottom_out[9] ,
    \sb_1__1__11_chany_bottom_out[10] ,
    \sb_1__1__11_chany_bottom_out[11] ,
    \sb_1__1__11_chany_bottom_out[12] ,
    \sb_1__1__11_chany_bottom_out[13] ,
    \sb_1__1__11_chany_bottom_out[14] ,
    \sb_1__1__11_chany_bottom_out[15] ,
    \sb_1__1__11_chany_bottom_out[16] ,
    \sb_1__1__11_chany_bottom_out[17] ,
    \sb_1__1__11_chany_bottom_out[18] ,
    \sb_1__1__11_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__13_chany_bottom_out[0] ,
    \cby_1__1__13_chany_bottom_out[1] ,
    \cby_1__1__13_chany_bottom_out[2] ,
    \cby_1__1__13_chany_bottom_out[3] ,
    \cby_1__1__13_chany_bottom_out[4] ,
    \cby_1__1__13_chany_bottom_out[5] ,
    \cby_1__1__13_chany_bottom_out[6] ,
    \cby_1__1__13_chany_bottom_out[7] ,
    \cby_1__1__13_chany_bottom_out[8] ,
    \cby_1__1__13_chany_bottom_out[9] ,
    \cby_1__1__13_chany_bottom_out[10] ,
    \cby_1__1__13_chany_bottom_out[11] ,
    \cby_1__1__13_chany_bottom_out[12] ,
    \cby_1__1__13_chany_bottom_out[13] ,
    \cby_1__1__13_chany_bottom_out[14] ,
    \cby_1__1__13_chany_bottom_out[15] ,
    \cby_1__1__13_chany_bottom_out[16] ,
    \cby_1__1__13_chany_bottom_out[17] ,
    \cby_1__1__13_chany_bottom_out[18] ,
    \cby_1__1__13_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__11_chany_top_out[0] ,
    \sb_1__1__11_chany_top_out[1] ,
    \sb_1__1__11_chany_top_out[2] ,
    \sb_1__1__11_chany_top_out[3] ,
    \sb_1__1__11_chany_top_out[4] ,
    \sb_1__1__11_chany_top_out[5] ,
    \sb_1__1__11_chany_top_out[6] ,
    \sb_1__1__11_chany_top_out[7] ,
    \sb_1__1__11_chany_top_out[8] ,
    \sb_1__1__11_chany_top_out[9] ,
    \sb_1__1__11_chany_top_out[10] ,
    \sb_1__1__11_chany_top_out[11] ,
    \sb_1__1__11_chany_top_out[12] ,
    \sb_1__1__11_chany_top_out[13] ,
    \sb_1__1__11_chany_top_out[14] ,
    \sb_1__1__11_chany_top_out[15] ,
    \sb_1__1__11_chany_top_out[16] ,
    \sb_1__1__11_chany_top_out[17] ,
    \sb_1__1__11_chany_top_out[18] ,
    \sb_1__1__11_chany_top_out[19] }));
 sb_1__1_ sb_2__6_ (.bottom_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__19_ccff_tail),
    .ccff_tail(sb_1__1__12_ccff_tail),
    .clk_2_E_out(\clk_2_wires[14] ),
    .clk_2_N_in(\clk_3_wires[15] ),
    .clk_2_W_out(\clk_2_wires[16] ),
    .left_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[63] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[14] ),
    .prog_clk_2_N_in(\prog_clk_3_wires[15] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[16] ),
    .right_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__12_chanx_right_out[0] ,
    \cbx_1__1__12_chanx_right_out[1] ,
    \cbx_1__1__12_chanx_right_out[2] ,
    \cbx_1__1__12_chanx_right_out[3] ,
    \cbx_1__1__12_chanx_right_out[4] ,
    \cbx_1__1__12_chanx_right_out[5] ,
    \cbx_1__1__12_chanx_right_out[6] ,
    \cbx_1__1__12_chanx_right_out[7] ,
    \cbx_1__1__12_chanx_right_out[8] ,
    \cbx_1__1__12_chanx_right_out[9] ,
    \cbx_1__1__12_chanx_right_out[10] ,
    \cbx_1__1__12_chanx_right_out[11] ,
    \cbx_1__1__12_chanx_right_out[12] ,
    \cbx_1__1__12_chanx_right_out[13] ,
    \cbx_1__1__12_chanx_right_out[14] ,
    \cbx_1__1__12_chanx_right_out[15] ,
    \cbx_1__1__12_chanx_right_out[16] ,
    \cbx_1__1__12_chanx_right_out[17] ,
    \cbx_1__1__12_chanx_right_out[18] ,
    \cbx_1__1__12_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__12_chanx_left_out[0] ,
    \sb_1__1__12_chanx_left_out[1] ,
    \sb_1__1__12_chanx_left_out[2] ,
    \sb_1__1__12_chanx_left_out[3] ,
    \sb_1__1__12_chanx_left_out[4] ,
    \sb_1__1__12_chanx_left_out[5] ,
    \sb_1__1__12_chanx_left_out[6] ,
    \sb_1__1__12_chanx_left_out[7] ,
    \sb_1__1__12_chanx_left_out[8] ,
    \sb_1__1__12_chanx_left_out[9] ,
    \sb_1__1__12_chanx_left_out[10] ,
    \sb_1__1__12_chanx_left_out[11] ,
    \sb_1__1__12_chanx_left_out[12] ,
    \sb_1__1__12_chanx_left_out[13] ,
    \sb_1__1__12_chanx_left_out[14] ,
    \sb_1__1__12_chanx_left_out[15] ,
    \sb_1__1__12_chanx_left_out[16] ,
    \sb_1__1__12_chanx_left_out[17] ,
    \sb_1__1__12_chanx_left_out[18] ,
    \sb_1__1__12_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__19_chanx_left_out[0] ,
    \cbx_1__1__19_chanx_left_out[1] ,
    \cbx_1__1__19_chanx_left_out[2] ,
    \cbx_1__1__19_chanx_left_out[3] ,
    \cbx_1__1__19_chanx_left_out[4] ,
    \cbx_1__1__19_chanx_left_out[5] ,
    \cbx_1__1__19_chanx_left_out[6] ,
    \cbx_1__1__19_chanx_left_out[7] ,
    \cbx_1__1__19_chanx_left_out[8] ,
    \cbx_1__1__19_chanx_left_out[9] ,
    \cbx_1__1__19_chanx_left_out[10] ,
    \cbx_1__1__19_chanx_left_out[11] ,
    \cbx_1__1__19_chanx_left_out[12] ,
    \cbx_1__1__19_chanx_left_out[13] ,
    \cbx_1__1__19_chanx_left_out[14] ,
    \cbx_1__1__19_chanx_left_out[15] ,
    \cbx_1__1__19_chanx_left_out[16] ,
    \cbx_1__1__19_chanx_left_out[17] ,
    \cbx_1__1__19_chanx_left_out[18] ,
    \cbx_1__1__19_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__12_chanx_right_out[0] ,
    \sb_1__1__12_chanx_right_out[1] ,
    \sb_1__1__12_chanx_right_out[2] ,
    \sb_1__1__12_chanx_right_out[3] ,
    \sb_1__1__12_chanx_right_out[4] ,
    \sb_1__1__12_chanx_right_out[5] ,
    \sb_1__1__12_chanx_right_out[6] ,
    \sb_1__1__12_chanx_right_out[7] ,
    \sb_1__1__12_chanx_right_out[8] ,
    \sb_1__1__12_chanx_right_out[9] ,
    \sb_1__1__12_chanx_right_out[10] ,
    \sb_1__1__12_chanx_right_out[11] ,
    \sb_1__1__12_chanx_right_out[12] ,
    \sb_1__1__12_chanx_right_out[13] ,
    \sb_1__1__12_chanx_right_out[14] ,
    \sb_1__1__12_chanx_right_out[15] ,
    \sb_1__1__12_chanx_right_out[16] ,
    \sb_1__1__12_chanx_right_out[17] ,
    \sb_1__1__12_chanx_right_out[18] ,
    \sb_1__1__12_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__13_chany_top_out[0] ,
    \cby_1__1__13_chany_top_out[1] ,
    \cby_1__1__13_chany_top_out[2] ,
    \cby_1__1__13_chany_top_out[3] ,
    \cby_1__1__13_chany_top_out[4] ,
    \cby_1__1__13_chany_top_out[5] ,
    \cby_1__1__13_chany_top_out[6] ,
    \cby_1__1__13_chany_top_out[7] ,
    \cby_1__1__13_chany_top_out[8] ,
    \cby_1__1__13_chany_top_out[9] ,
    \cby_1__1__13_chany_top_out[10] ,
    \cby_1__1__13_chany_top_out[11] ,
    \cby_1__1__13_chany_top_out[12] ,
    \cby_1__1__13_chany_top_out[13] ,
    \cby_1__1__13_chany_top_out[14] ,
    \cby_1__1__13_chany_top_out[15] ,
    \cby_1__1__13_chany_top_out[16] ,
    \cby_1__1__13_chany_top_out[17] ,
    \cby_1__1__13_chany_top_out[18] ,
    \cby_1__1__13_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__12_chany_bottom_out[0] ,
    \sb_1__1__12_chany_bottom_out[1] ,
    \sb_1__1__12_chany_bottom_out[2] ,
    \sb_1__1__12_chany_bottom_out[3] ,
    \sb_1__1__12_chany_bottom_out[4] ,
    \sb_1__1__12_chany_bottom_out[5] ,
    \sb_1__1__12_chany_bottom_out[6] ,
    \sb_1__1__12_chany_bottom_out[7] ,
    \sb_1__1__12_chany_bottom_out[8] ,
    \sb_1__1__12_chany_bottom_out[9] ,
    \sb_1__1__12_chany_bottom_out[10] ,
    \sb_1__1__12_chany_bottom_out[11] ,
    \sb_1__1__12_chany_bottom_out[12] ,
    \sb_1__1__12_chany_bottom_out[13] ,
    \sb_1__1__12_chany_bottom_out[14] ,
    \sb_1__1__12_chany_bottom_out[15] ,
    \sb_1__1__12_chany_bottom_out[16] ,
    \sb_1__1__12_chany_bottom_out[17] ,
    \sb_1__1__12_chany_bottom_out[18] ,
    \sb_1__1__12_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__14_chany_bottom_out[0] ,
    \cby_1__1__14_chany_bottom_out[1] ,
    \cby_1__1__14_chany_bottom_out[2] ,
    \cby_1__1__14_chany_bottom_out[3] ,
    \cby_1__1__14_chany_bottom_out[4] ,
    \cby_1__1__14_chany_bottom_out[5] ,
    \cby_1__1__14_chany_bottom_out[6] ,
    \cby_1__1__14_chany_bottom_out[7] ,
    \cby_1__1__14_chany_bottom_out[8] ,
    \cby_1__1__14_chany_bottom_out[9] ,
    \cby_1__1__14_chany_bottom_out[10] ,
    \cby_1__1__14_chany_bottom_out[11] ,
    \cby_1__1__14_chany_bottom_out[12] ,
    \cby_1__1__14_chany_bottom_out[13] ,
    \cby_1__1__14_chany_bottom_out[14] ,
    \cby_1__1__14_chany_bottom_out[15] ,
    \cby_1__1__14_chany_bottom_out[16] ,
    \cby_1__1__14_chany_bottom_out[17] ,
    \cby_1__1__14_chany_bottom_out[18] ,
    \cby_1__1__14_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__12_chany_top_out[0] ,
    \sb_1__1__12_chany_top_out[1] ,
    \sb_1__1__12_chany_top_out[2] ,
    \sb_1__1__12_chany_top_out[3] ,
    \sb_1__1__12_chany_top_out[4] ,
    \sb_1__1__12_chany_top_out[5] ,
    \sb_1__1__12_chany_top_out[6] ,
    \sb_1__1__12_chany_top_out[7] ,
    \sb_1__1__12_chany_top_out[8] ,
    \sb_1__1__12_chany_top_out[9] ,
    \sb_1__1__12_chany_top_out[10] ,
    \sb_1__1__12_chany_top_out[11] ,
    \sb_1__1__12_chany_top_out[12] ,
    \sb_1__1__12_chany_top_out[13] ,
    \sb_1__1__12_chany_top_out[14] ,
    \sb_1__1__12_chany_top_out[15] ,
    \sb_1__1__12_chany_top_out[16] ,
    \sb_1__1__12_chany_top_out[17] ,
    \sb_1__1__12_chany_top_out[18] ,
    \sb_1__1__12_chany_top_out[19] }));
 sb_1__1_ sb_2__7_ (.bottom_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__20_ccff_tail),
    .ccff_tail(sb_1__1__13_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[66] ),
    .right_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__13_chanx_right_out[0] ,
    \cbx_1__1__13_chanx_right_out[1] ,
    \cbx_1__1__13_chanx_right_out[2] ,
    \cbx_1__1__13_chanx_right_out[3] ,
    \cbx_1__1__13_chanx_right_out[4] ,
    \cbx_1__1__13_chanx_right_out[5] ,
    \cbx_1__1__13_chanx_right_out[6] ,
    \cbx_1__1__13_chanx_right_out[7] ,
    \cbx_1__1__13_chanx_right_out[8] ,
    \cbx_1__1__13_chanx_right_out[9] ,
    \cbx_1__1__13_chanx_right_out[10] ,
    \cbx_1__1__13_chanx_right_out[11] ,
    \cbx_1__1__13_chanx_right_out[12] ,
    \cbx_1__1__13_chanx_right_out[13] ,
    \cbx_1__1__13_chanx_right_out[14] ,
    \cbx_1__1__13_chanx_right_out[15] ,
    \cbx_1__1__13_chanx_right_out[16] ,
    \cbx_1__1__13_chanx_right_out[17] ,
    \cbx_1__1__13_chanx_right_out[18] ,
    \cbx_1__1__13_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__13_chanx_left_out[0] ,
    \sb_1__1__13_chanx_left_out[1] ,
    \sb_1__1__13_chanx_left_out[2] ,
    \sb_1__1__13_chanx_left_out[3] ,
    \sb_1__1__13_chanx_left_out[4] ,
    \sb_1__1__13_chanx_left_out[5] ,
    \sb_1__1__13_chanx_left_out[6] ,
    \sb_1__1__13_chanx_left_out[7] ,
    \sb_1__1__13_chanx_left_out[8] ,
    \sb_1__1__13_chanx_left_out[9] ,
    \sb_1__1__13_chanx_left_out[10] ,
    \sb_1__1__13_chanx_left_out[11] ,
    \sb_1__1__13_chanx_left_out[12] ,
    \sb_1__1__13_chanx_left_out[13] ,
    \sb_1__1__13_chanx_left_out[14] ,
    \sb_1__1__13_chanx_left_out[15] ,
    \sb_1__1__13_chanx_left_out[16] ,
    \sb_1__1__13_chanx_left_out[17] ,
    \sb_1__1__13_chanx_left_out[18] ,
    \sb_1__1__13_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__20_chanx_left_out[0] ,
    \cbx_1__1__20_chanx_left_out[1] ,
    \cbx_1__1__20_chanx_left_out[2] ,
    \cbx_1__1__20_chanx_left_out[3] ,
    \cbx_1__1__20_chanx_left_out[4] ,
    \cbx_1__1__20_chanx_left_out[5] ,
    \cbx_1__1__20_chanx_left_out[6] ,
    \cbx_1__1__20_chanx_left_out[7] ,
    \cbx_1__1__20_chanx_left_out[8] ,
    \cbx_1__1__20_chanx_left_out[9] ,
    \cbx_1__1__20_chanx_left_out[10] ,
    \cbx_1__1__20_chanx_left_out[11] ,
    \cbx_1__1__20_chanx_left_out[12] ,
    \cbx_1__1__20_chanx_left_out[13] ,
    \cbx_1__1__20_chanx_left_out[14] ,
    \cbx_1__1__20_chanx_left_out[15] ,
    \cbx_1__1__20_chanx_left_out[16] ,
    \cbx_1__1__20_chanx_left_out[17] ,
    \cbx_1__1__20_chanx_left_out[18] ,
    \cbx_1__1__20_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__13_chanx_right_out[0] ,
    \sb_1__1__13_chanx_right_out[1] ,
    \sb_1__1__13_chanx_right_out[2] ,
    \sb_1__1__13_chanx_right_out[3] ,
    \sb_1__1__13_chanx_right_out[4] ,
    \sb_1__1__13_chanx_right_out[5] ,
    \sb_1__1__13_chanx_right_out[6] ,
    \sb_1__1__13_chanx_right_out[7] ,
    \sb_1__1__13_chanx_right_out[8] ,
    \sb_1__1__13_chanx_right_out[9] ,
    \sb_1__1__13_chanx_right_out[10] ,
    \sb_1__1__13_chanx_right_out[11] ,
    \sb_1__1__13_chanx_right_out[12] ,
    \sb_1__1__13_chanx_right_out[13] ,
    \sb_1__1__13_chanx_right_out[14] ,
    \sb_1__1__13_chanx_right_out[15] ,
    \sb_1__1__13_chanx_right_out[16] ,
    \sb_1__1__13_chanx_right_out[17] ,
    \sb_1__1__13_chanx_right_out[18] ,
    \sb_1__1__13_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__14_chany_top_out[0] ,
    \cby_1__1__14_chany_top_out[1] ,
    \cby_1__1__14_chany_top_out[2] ,
    \cby_1__1__14_chany_top_out[3] ,
    \cby_1__1__14_chany_top_out[4] ,
    \cby_1__1__14_chany_top_out[5] ,
    \cby_1__1__14_chany_top_out[6] ,
    \cby_1__1__14_chany_top_out[7] ,
    \cby_1__1__14_chany_top_out[8] ,
    \cby_1__1__14_chany_top_out[9] ,
    \cby_1__1__14_chany_top_out[10] ,
    \cby_1__1__14_chany_top_out[11] ,
    \cby_1__1__14_chany_top_out[12] ,
    \cby_1__1__14_chany_top_out[13] ,
    \cby_1__1__14_chany_top_out[14] ,
    \cby_1__1__14_chany_top_out[15] ,
    \cby_1__1__14_chany_top_out[16] ,
    \cby_1__1__14_chany_top_out[17] ,
    \cby_1__1__14_chany_top_out[18] ,
    \cby_1__1__14_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__13_chany_bottom_out[0] ,
    \sb_1__1__13_chany_bottom_out[1] ,
    \sb_1__1__13_chany_bottom_out[2] ,
    \sb_1__1__13_chany_bottom_out[3] ,
    \sb_1__1__13_chany_bottom_out[4] ,
    \sb_1__1__13_chany_bottom_out[5] ,
    \sb_1__1__13_chany_bottom_out[6] ,
    \sb_1__1__13_chany_bottom_out[7] ,
    \sb_1__1__13_chany_bottom_out[8] ,
    \sb_1__1__13_chany_bottom_out[9] ,
    \sb_1__1__13_chany_bottom_out[10] ,
    \sb_1__1__13_chany_bottom_out[11] ,
    \sb_1__1__13_chany_bottom_out[12] ,
    \sb_1__1__13_chany_bottom_out[13] ,
    \sb_1__1__13_chany_bottom_out[14] ,
    \sb_1__1__13_chany_bottom_out[15] ,
    \sb_1__1__13_chany_bottom_out[16] ,
    \sb_1__1__13_chany_bottom_out[17] ,
    \sb_1__1__13_chany_bottom_out[18] ,
    \sb_1__1__13_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__15_chany_bottom_out[0] ,
    \cby_1__1__15_chany_bottom_out[1] ,
    \cby_1__1__15_chany_bottom_out[2] ,
    \cby_1__1__15_chany_bottom_out[3] ,
    \cby_1__1__15_chany_bottom_out[4] ,
    \cby_1__1__15_chany_bottom_out[5] ,
    \cby_1__1__15_chany_bottom_out[6] ,
    \cby_1__1__15_chany_bottom_out[7] ,
    \cby_1__1__15_chany_bottom_out[8] ,
    \cby_1__1__15_chany_bottom_out[9] ,
    \cby_1__1__15_chany_bottom_out[10] ,
    \cby_1__1__15_chany_bottom_out[11] ,
    \cby_1__1__15_chany_bottom_out[12] ,
    \cby_1__1__15_chany_bottom_out[13] ,
    \cby_1__1__15_chany_bottom_out[14] ,
    \cby_1__1__15_chany_bottom_out[15] ,
    \cby_1__1__15_chany_bottom_out[16] ,
    \cby_1__1__15_chany_bottom_out[17] ,
    \cby_1__1__15_chany_bottom_out[18] ,
    \cby_1__1__15_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__13_chany_top_out[0] ,
    \sb_1__1__13_chany_top_out[1] ,
    \sb_1__1__13_chany_top_out[2] ,
    \sb_1__1__13_chany_top_out[3] ,
    \sb_1__1__13_chany_top_out[4] ,
    \sb_1__1__13_chany_top_out[5] ,
    \sb_1__1__13_chany_top_out[6] ,
    \sb_1__1__13_chany_top_out[7] ,
    \sb_1__1__13_chany_top_out[8] ,
    \sb_1__1__13_chany_top_out[9] ,
    \sb_1__1__13_chany_top_out[10] ,
    \sb_1__1__13_chany_top_out[11] ,
    \sb_1__1__13_chany_top_out[12] ,
    \sb_1__1__13_chany_top_out[13] ,
    \sb_1__1__13_chany_top_out[14] ,
    \sb_1__1__13_chany_top_out[15] ,
    \sb_1__1__13_chany_top_out[16] ,
    \sb_1__1__13_chany_top_out[17] ,
    \sb_1__1__13_chany_top_out[18] ,
    \sb_1__1__13_chany_top_out[19] }));
 sb_1__2_ sb_2__8_ (.SC_IN_BOT(\scff_Wires[36] ),
    .SC_OUT_BOT(\scff_Wires[37] ),
    .bottom_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_upper),
    .ccff_head(grid_io_top_2_ccff_tail),
    .ccff_tail(sb_1__8__1_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[68] ),
    .right_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__1_chanx_right_out[0] ,
    \cbx_1__8__1_chanx_right_out[1] ,
    \cbx_1__8__1_chanx_right_out[2] ,
    \cbx_1__8__1_chanx_right_out[3] ,
    \cbx_1__8__1_chanx_right_out[4] ,
    \cbx_1__8__1_chanx_right_out[5] ,
    \cbx_1__8__1_chanx_right_out[6] ,
    \cbx_1__8__1_chanx_right_out[7] ,
    \cbx_1__8__1_chanx_right_out[8] ,
    \cbx_1__8__1_chanx_right_out[9] ,
    \cbx_1__8__1_chanx_right_out[10] ,
    \cbx_1__8__1_chanx_right_out[11] ,
    \cbx_1__8__1_chanx_right_out[12] ,
    \cbx_1__8__1_chanx_right_out[13] ,
    \cbx_1__8__1_chanx_right_out[14] ,
    \cbx_1__8__1_chanx_right_out[15] ,
    \cbx_1__8__1_chanx_right_out[16] ,
    \cbx_1__8__1_chanx_right_out[17] ,
    \cbx_1__8__1_chanx_right_out[18] ,
    \cbx_1__8__1_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__8__1_chanx_left_out[0] ,
    \sb_1__8__1_chanx_left_out[1] ,
    \sb_1__8__1_chanx_left_out[2] ,
    \sb_1__8__1_chanx_left_out[3] ,
    \sb_1__8__1_chanx_left_out[4] ,
    \sb_1__8__1_chanx_left_out[5] ,
    \sb_1__8__1_chanx_left_out[6] ,
    \sb_1__8__1_chanx_left_out[7] ,
    \sb_1__8__1_chanx_left_out[8] ,
    \sb_1__8__1_chanx_left_out[9] ,
    \sb_1__8__1_chanx_left_out[10] ,
    \sb_1__8__1_chanx_left_out[11] ,
    \sb_1__8__1_chanx_left_out[12] ,
    \sb_1__8__1_chanx_left_out[13] ,
    \sb_1__8__1_chanx_left_out[14] ,
    \sb_1__8__1_chanx_left_out[15] ,
    \sb_1__8__1_chanx_left_out[16] ,
    \sb_1__8__1_chanx_left_out[17] ,
    \sb_1__8__1_chanx_left_out[18] ,
    \sb_1__8__1_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__8__2_chanx_left_out[0] ,
    \cbx_1__8__2_chanx_left_out[1] ,
    \cbx_1__8__2_chanx_left_out[2] ,
    \cbx_1__8__2_chanx_left_out[3] ,
    \cbx_1__8__2_chanx_left_out[4] ,
    \cbx_1__8__2_chanx_left_out[5] ,
    \cbx_1__8__2_chanx_left_out[6] ,
    \cbx_1__8__2_chanx_left_out[7] ,
    \cbx_1__8__2_chanx_left_out[8] ,
    \cbx_1__8__2_chanx_left_out[9] ,
    \cbx_1__8__2_chanx_left_out[10] ,
    \cbx_1__8__2_chanx_left_out[11] ,
    \cbx_1__8__2_chanx_left_out[12] ,
    \cbx_1__8__2_chanx_left_out[13] ,
    \cbx_1__8__2_chanx_left_out[14] ,
    \cbx_1__8__2_chanx_left_out[15] ,
    \cbx_1__8__2_chanx_left_out[16] ,
    \cbx_1__8__2_chanx_left_out[17] ,
    \cbx_1__8__2_chanx_left_out[18] ,
    \cbx_1__8__2_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__8__1_chanx_right_out[0] ,
    \sb_1__8__1_chanx_right_out[1] ,
    \sb_1__8__1_chanx_right_out[2] ,
    \sb_1__8__1_chanx_right_out[3] ,
    \sb_1__8__1_chanx_right_out[4] ,
    \sb_1__8__1_chanx_right_out[5] ,
    \sb_1__8__1_chanx_right_out[6] ,
    \sb_1__8__1_chanx_right_out[7] ,
    \sb_1__8__1_chanx_right_out[8] ,
    \sb_1__8__1_chanx_right_out[9] ,
    \sb_1__8__1_chanx_right_out[10] ,
    \sb_1__8__1_chanx_right_out[11] ,
    \sb_1__8__1_chanx_right_out[12] ,
    \sb_1__8__1_chanx_right_out[13] ,
    \sb_1__8__1_chanx_right_out[14] ,
    \sb_1__8__1_chanx_right_out[15] ,
    \sb_1__8__1_chanx_right_out[16] ,
    \sb_1__8__1_chanx_right_out[17] ,
    \sb_1__8__1_chanx_right_out[18] ,
    \sb_1__8__1_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__15_chany_top_out[0] ,
    \cby_1__1__15_chany_top_out[1] ,
    \cby_1__1__15_chany_top_out[2] ,
    \cby_1__1__15_chany_top_out[3] ,
    \cby_1__1__15_chany_top_out[4] ,
    \cby_1__1__15_chany_top_out[5] ,
    \cby_1__1__15_chany_top_out[6] ,
    \cby_1__1__15_chany_top_out[7] ,
    \cby_1__1__15_chany_top_out[8] ,
    \cby_1__1__15_chany_top_out[9] ,
    \cby_1__1__15_chany_top_out[10] ,
    \cby_1__1__15_chany_top_out[11] ,
    \cby_1__1__15_chany_top_out[12] ,
    \cby_1__1__15_chany_top_out[13] ,
    \cby_1__1__15_chany_top_out[14] ,
    \cby_1__1__15_chany_top_out[15] ,
    \cby_1__1__15_chany_top_out[16] ,
    \cby_1__1__15_chany_top_out[17] ,
    \cby_1__1__15_chany_top_out[18] ,
    \cby_1__1__15_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__8__1_chany_bottom_out[0] ,
    \sb_1__8__1_chany_bottom_out[1] ,
    \sb_1__8__1_chany_bottom_out[2] ,
    \sb_1__8__1_chany_bottom_out[3] ,
    \sb_1__8__1_chany_bottom_out[4] ,
    \sb_1__8__1_chany_bottom_out[5] ,
    \sb_1__8__1_chany_bottom_out[6] ,
    \sb_1__8__1_chany_bottom_out[7] ,
    \sb_1__8__1_chany_bottom_out[8] ,
    \sb_1__8__1_chany_bottom_out[9] ,
    \sb_1__8__1_chany_bottom_out[10] ,
    \sb_1__8__1_chany_bottom_out[11] ,
    \sb_1__8__1_chany_bottom_out[12] ,
    \sb_1__8__1_chany_bottom_out[13] ,
    \sb_1__8__1_chany_bottom_out[14] ,
    \sb_1__8__1_chany_bottom_out[15] ,
    \sb_1__8__1_chany_bottom_out[16] ,
    \sb_1__8__1_chany_bottom_out[17] ,
    \sb_1__8__1_chany_bottom_out[18] ,
    \sb_1__8__1_chany_bottom_out[19] }));
 sb_1__0_ sb_3__0_ (.SC_IN_TOP(\scff_Wires[55] ),
    .SC_OUT_TOP(\scff_Wires[56] ),
    .ccff_head(grid_io_bottom_4_ccff_tail),
    .ccff_tail(sb_1__0__2_ccff_tail),
    .left_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[71] ),
    .right_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__2_chanx_right_out[0] ,
    \cbx_1__0__2_chanx_right_out[1] ,
    \cbx_1__0__2_chanx_right_out[2] ,
    \cbx_1__0__2_chanx_right_out[3] ,
    \cbx_1__0__2_chanx_right_out[4] ,
    \cbx_1__0__2_chanx_right_out[5] ,
    \cbx_1__0__2_chanx_right_out[6] ,
    \cbx_1__0__2_chanx_right_out[7] ,
    \cbx_1__0__2_chanx_right_out[8] ,
    \cbx_1__0__2_chanx_right_out[9] ,
    \cbx_1__0__2_chanx_right_out[10] ,
    \cbx_1__0__2_chanx_right_out[11] ,
    \cbx_1__0__2_chanx_right_out[12] ,
    \cbx_1__0__2_chanx_right_out[13] ,
    \cbx_1__0__2_chanx_right_out[14] ,
    \cbx_1__0__2_chanx_right_out[15] ,
    \cbx_1__0__2_chanx_right_out[16] ,
    \cbx_1__0__2_chanx_right_out[17] ,
    \cbx_1__0__2_chanx_right_out[18] ,
    \cbx_1__0__2_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__0__2_chanx_left_out[0] ,
    \sb_1__0__2_chanx_left_out[1] ,
    \sb_1__0__2_chanx_left_out[2] ,
    \sb_1__0__2_chanx_left_out[3] ,
    \sb_1__0__2_chanx_left_out[4] ,
    \sb_1__0__2_chanx_left_out[5] ,
    \sb_1__0__2_chanx_left_out[6] ,
    \sb_1__0__2_chanx_left_out[7] ,
    \sb_1__0__2_chanx_left_out[8] ,
    \sb_1__0__2_chanx_left_out[9] ,
    \sb_1__0__2_chanx_left_out[10] ,
    \sb_1__0__2_chanx_left_out[11] ,
    \sb_1__0__2_chanx_left_out[12] ,
    \sb_1__0__2_chanx_left_out[13] ,
    \sb_1__0__2_chanx_left_out[14] ,
    \sb_1__0__2_chanx_left_out[15] ,
    \sb_1__0__2_chanx_left_out[16] ,
    \sb_1__0__2_chanx_left_out[17] ,
    \sb_1__0__2_chanx_left_out[18] ,
    \sb_1__0__2_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__0__3_chanx_left_out[0] ,
    \cbx_1__0__3_chanx_left_out[1] ,
    \cbx_1__0__3_chanx_left_out[2] ,
    \cbx_1__0__3_chanx_left_out[3] ,
    \cbx_1__0__3_chanx_left_out[4] ,
    \cbx_1__0__3_chanx_left_out[5] ,
    \cbx_1__0__3_chanx_left_out[6] ,
    \cbx_1__0__3_chanx_left_out[7] ,
    \cbx_1__0__3_chanx_left_out[8] ,
    \cbx_1__0__3_chanx_left_out[9] ,
    \cbx_1__0__3_chanx_left_out[10] ,
    \cbx_1__0__3_chanx_left_out[11] ,
    \cbx_1__0__3_chanx_left_out[12] ,
    \cbx_1__0__3_chanx_left_out[13] ,
    \cbx_1__0__3_chanx_left_out[14] ,
    \cbx_1__0__3_chanx_left_out[15] ,
    \cbx_1__0__3_chanx_left_out[16] ,
    \cbx_1__0__3_chanx_left_out[17] ,
    \cbx_1__0__3_chanx_left_out[18] ,
    \cbx_1__0__3_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__0__2_chanx_right_out[0] ,
    \sb_1__0__2_chanx_right_out[1] ,
    \sb_1__0__2_chanx_right_out[2] ,
    \sb_1__0__2_chanx_right_out[3] ,
    \sb_1__0__2_chanx_right_out[4] ,
    \sb_1__0__2_chanx_right_out[5] ,
    \sb_1__0__2_chanx_right_out[6] ,
    \sb_1__0__2_chanx_right_out[7] ,
    \sb_1__0__2_chanx_right_out[8] ,
    \sb_1__0__2_chanx_right_out[9] ,
    \sb_1__0__2_chanx_right_out[10] ,
    \sb_1__0__2_chanx_right_out[11] ,
    \sb_1__0__2_chanx_right_out[12] ,
    \sb_1__0__2_chanx_right_out[13] ,
    \sb_1__0__2_chanx_right_out[14] ,
    \sb_1__0__2_chanx_right_out[15] ,
    \sb_1__0__2_chanx_right_out[16] ,
    \sb_1__0__2_chanx_right_out[17] ,
    \sb_1__0__2_chanx_right_out[18] ,
    \sb_1__0__2_chanx_right_out[19] }),
    .chany_top_in({\cby_1__1__16_chany_bottom_out[0] ,
    \cby_1__1__16_chany_bottom_out[1] ,
    \cby_1__1__16_chany_bottom_out[2] ,
    \cby_1__1__16_chany_bottom_out[3] ,
    \cby_1__1__16_chany_bottom_out[4] ,
    \cby_1__1__16_chany_bottom_out[5] ,
    \cby_1__1__16_chany_bottom_out[6] ,
    \cby_1__1__16_chany_bottom_out[7] ,
    \cby_1__1__16_chany_bottom_out[8] ,
    \cby_1__1__16_chany_bottom_out[9] ,
    \cby_1__1__16_chany_bottom_out[10] ,
    \cby_1__1__16_chany_bottom_out[11] ,
    \cby_1__1__16_chany_bottom_out[12] ,
    \cby_1__1__16_chany_bottom_out[13] ,
    \cby_1__1__16_chany_bottom_out[14] ,
    \cby_1__1__16_chany_bottom_out[15] ,
    \cby_1__1__16_chany_bottom_out[16] ,
    \cby_1__1__16_chany_bottom_out[17] ,
    \cby_1__1__16_chany_bottom_out[18] ,
    \cby_1__1__16_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__0__2_chany_top_out[0] ,
    \sb_1__0__2_chany_top_out[1] ,
    \sb_1__0__2_chany_top_out[2] ,
    \sb_1__0__2_chany_top_out[3] ,
    \sb_1__0__2_chany_top_out[4] ,
    \sb_1__0__2_chany_top_out[5] ,
    \sb_1__0__2_chany_top_out[6] ,
    \sb_1__0__2_chany_top_out[7] ,
    \sb_1__0__2_chany_top_out[8] ,
    \sb_1__0__2_chany_top_out[9] ,
    \sb_1__0__2_chany_top_out[10] ,
    \sb_1__0__2_chany_top_out[11] ,
    \sb_1__0__2_chany_top_out[12] ,
    \sb_1__0__2_chany_top_out[13] ,
    \sb_1__0__2_chany_top_out[14] ,
    \sb_1__0__2_chany_top_out[15] ,
    \sb_1__0__2_chany_top_out[16] ,
    \sb_1__0__2_chany_top_out[17] ,
    \sb_1__0__2_chany_top_out[18] ,
    \sb_1__0__2_chany_top_out[19] }));
 sb_1__1_ sb_3__1_ (.bottom_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__21_ccff_tail),
    .ccff_tail(sb_1__1__14_ccff_tail),
    .clk_1_E_out(\clk_1_wires[29] ),
    .clk_1_N_in(\clk_2_wires[12] ),
    .clk_1_W_out(\clk_1_wires[30] ),
    .left_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[74] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[29] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[12] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[30] ),
    .right_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__14_chanx_right_out[0] ,
    \cbx_1__1__14_chanx_right_out[1] ,
    \cbx_1__1__14_chanx_right_out[2] ,
    \cbx_1__1__14_chanx_right_out[3] ,
    \cbx_1__1__14_chanx_right_out[4] ,
    \cbx_1__1__14_chanx_right_out[5] ,
    \cbx_1__1__14_chanx_right_out[6] ,
    \cbx_1__1__14_chanx_right_out[7] ,
    \cbx_1__1__14_chanx_right_out[8] ,
    \cbx_1__1__14_chanx_right_out[9] ,
    \cbx_1__1__14_chanx_right_out[10] ,
    \cbx_1__1__14_chanx_right_out[11] ,
    \cbx_1__1__14_chanx_right_out[12] ,
    \cbx_1__1__14_chanx_right_out[13] ,
    \cbx_1__1__14_chanx_right_out[14] ,
    \cbx_1__1__14_chanx_right_out[15] ,
    \cbx_1__1__14_chanx_right_out[16] ,
    \cbx_1__1__14_chanx_right_out[17] ,
    \cbx_1__1__14_chanx_right_out[18] ,
    \cbx_1__1__14_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__14_chanx_left_out[0] ,
    \sb_1__1__14_chanx_left_out[1] ,
    \sb_1__1__14_chanx_left_out[2] ,
    \sb_1__1__14_chanx_left_out[3] ,
    \sb_1__1__14_chanx_left_out[4] ,
    \sb_1__1__14_chanx_left_out[5] ,
    \sb_1__1__14_chanx_left_out[6] ,
    \sb_1__1__14_chanx_left_out[7] ,
    \sb_1__1__14_chanx_left_out[8] ,
    \sb_1__1__14_chanx_left_out[9] ,
    \sb_1__1__14_chanx_left_out[10] ,
    \sb_1__1__14_chanx_left_out[11] ,
    \sb_1__1__14_chanx_left_out[12] ,
    \sb_1__1__14_chanx_left_out[13] ,
    \sb_1__1__14_chanx_left_out[14] ,
    \sb_1__1__14_chanx_left_out[15] ,
    \sb_1__1__14_chanx_left_out[16] ,
    \sb_1__1__14_chanx_left_out[17] ,
    \sb_1__1__14_chanx_left_out[18] ,
    \sb_1__1__14_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__21_chanx_left_out[0] ,
    \cbx_1__1__21_chanx_left_out[1] ,
    \cbx_1__1__21_chanx_left_out[2] ,
    \cbx_1__1__21_chanx_left_out[3] ,
    \cbx_1__1__21_chanx_left_out[4] ,
    \cbx_1__1__21_chanx_left_out[5] ,
    \cbx_1__1__21_chanx_left_out[6] ,
    \cbx_1__1__21_chanx_left_out[7] ,
    \cbx_1__1__21_chanx_left_out[8] ,
    \cbx_1__1__21_chanx_left_out[9] ,
    \cbx_1__1__21_chanx_left_out[10] ,
    \cbx_1__1__21_chanx_left_out[11] ,
    \cbx_1__1__21_chanx_left_out[12] ,
    \cbx_1__1__21_chanx_left_out[13] ,
    \cbx_1__1__21_chanx_left_out[14] ,
    \cbx_1__1__21_chanx_left_out[15] ,
    \cbx_1__1__21_chanx_left_out[16] ,
    \cbx_1__1__21_chanx_left_out[17] ,
    \cbx_1__1__21_chanx_left_out[18] ,
    \cbx_1__1__21_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__14_chanx_right_out[0] ,
    \sb_1__1__14_chanx_right_out[1] ,
    \sb_1__1__14_chanx_right_out[2] ,
    \sb_1__1__14_chanx_right_out[3] ,
    \sb_1__1__14_chanx_right_out[4] ,
    \sb_1__1__14_chanx_right_out[5] ,
    \sb_1__1__14_chanx_right_out[6] ,
    \sb_1__1__14_chanx_right_out[7] ,
    \sb_1__1__14_chanx_right_out[8] ,
    \sb_1__1__14_chanx_right_out[9] ,
    \sb_1__1__14_chanx_right_out[10] ,
    \sb_1__1__14_chanx_right_out[11] ,
    \sb_1__1__14_chanx_right_out[12] ,
    \sb_1__1__14_chanx_right_out[13] ,
    \sb_1__1__14_chanx_right_out[14] ,
    \sb_1__1__14_chanx_right_out[15] ,
    \sb_1__1__14_chanx_right_out[16] ,
    \sb_1__1__14_chanx_right_out[17] ,
    \sb_1__1__14_chanx_right_out[18] ,
    \sb_1__1__14_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__16_chany_top_out[0] ,
    \cby_1__1__16_chany_top_out[1] ,
    \cby_1__1__16_chany_top_out[2] ,
    \cby_1__1__16_chany_top_out[3] ,
    \cby_1__1__16_chany_top_out[4] ,
    \cby_1__1__16_chany_top_out[5] ,
    \cby_1__1__16_chany_top_out[6] ,
    \cby_1__1__16_chany_top_out[7] ,
    \cby_1__1__16_chany_top_out[8] ,
    \cby_1__1__16_chany_top_out[9] ,
    \cby_1__1__16_chany_top_out[10] ,
    \cby_1__1__16_chany_top_out[11] ,
    \cby_1__1__16_chany_top_out[12] ,
    \cby_1__1__16_chany_top_out[13] ,
    \cby_1__1__16_chany_top_out[14] ,
    \cby_1__1__16_chany_top_out[15] ,
    \cby_1__1__16_chany_top_out[16] ,
    \cby_1__1__16_chany_top_out[17] ,
    \cby_1__1__16_chany_top_out[18] ,
    \cby_1__1__16_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__14_chany_bottom_out[0] ,
    \sb_1__1__14_chany_bottom_out[1] ,
    \sb_1__1__14_chany_bottom_out[2] ,
    \sb_1__1__14_chany_bottom_out[3] ,
    \sb_1__1__14_chany_bottom_out[4] ,
    \sb_1__1__14_chany_bottom_out[5] ,
    \sb_1__1__14_chany_bottom_out[6] ,
    \sb_1__1__14_chany_bottom_out[7] ,
    \sb_1__1__14_chany_bottom_out[8] ,
    \sb_1__1__14_chany_bottom_out[9] ,
    \sb_1__1__14_chany_bottom_out[10] ,
    \sb_1__1__14_chany_bottom_out[11] ,
    \sb_1__1__14_chany_bottom_out[12] ,
    \sb_1__1__14_chany_bottom_out[13] ,
    \sb_1__1__14_chany_bottom_out[14] ,
    \sb_1__1__14_chany_bottom_out[15] ,
    \sb_1__1__14_chany_bottom_out[16] ,
    \sb_1__1__14_chany_bottom_out[17] ,
    \sb_1__1__14_chany_bottom_out[18] ,
    \sb_1__1__14_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__17_chany_bottom_out[0] ,
    \cby_1__1__17_chany_bottom_out[1] ,
    \cby_1__1__17_chany_bottom_out[2] ,
    \cby_1__1__17_chany_bottom_out[3] ,
    \cby_1__1__17_chany_bottom_out[4] ,
    \cby_1__1__17_chany_bottom_out[5] ,
    \cby_1__1__17_chany_bottom_out[6] ,
    \cby_1__1__17_chany_bottom_out[7] ,
    \cby_1__1__17_chany_bottom_out[8] ,
    \cby_1__1__17_chany_bottom_out[9] ,
    \cby_1__1__17_chany_bottom_out[10] ,
    \cby_1__1__17_chany_bottom_out[11] ,
    \cby_1__1__17_chany_bottom_out[12] ,
    \cby_1__1__17_chany_bottom_out[13] ,
    \cby_1__1__17_chany_bottom_out[14] ,
    \cby_1__1__17_chany_bottom_out[15] ,
    \cby_1__1__17_chany_bottom_out[16] ,
    \cby_1__1__17_chany_bottom_out[17] ,
    \cby_1__1__17_chany_bottom_out[18] ,
    \cby_1__1__17_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__14_chany_top_out[0] ,
    \sb_1__1__14_chany_top_out[1] ,
    \sb_1__1__14_chany_top_out[2] ,
    \sb_1__1__14_chany_top_out[3] ,
    \sb_1__1__14_chany_top_out[4] ,
    \sb_1__1__14_chany_top_out[5] ,
    \sb_1__1__14_chany_top_out[6] ,
    \sb_1__1__14_chany_top_out[7] ,
    \sb_1__1__14_chany_top_out[8] ,
    \sb_1__1__14_chany_top_out[9] ,
    \sb_1__1__14_chany_top_out[10] ,
    \sb_1__1__14_chany_top_out[11] ,
    \sb_1__1__14_chany_top_out[12] ,
    \sb_1__1__14_chany_top_out[13] ,
    \sb_1__1__14_chany_top_out[14] ,
    \sb_1__1__14_chany_top_out[15] ,
    \sb_1__1__14_chany_top_out[16] ,
    \sb_1__1__14_chany_top_out[17] ,
    \sb_1__1__14_chany_top_out[18] ,
    \sb_1__1__14_chany_top_out[19] }));
 sb_1__1_ sb_3__2_ (.bottom_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__22_ccff_tail),
    .ccff_tail(sb_1__1__15_ccff_tail),
    .clk_2_N_in(\clk_2_wires[2] ),
    .clk_2_N_out(\clk_2_wires[9] ),
    .clk_2_S_out(\clk_2_wires[11] ),
    .left_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[77] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[2] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[9] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[11] ),
    .right_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__15_chanx_right_out[0] ,
    \cbx_1__1__15_chanx_right_out[1] ,
    \cbx_1__1__15_chanx_right_out[2] ,
    \cbx_1__1__15_chanx_right_out[3] ,
    \cbx_1__1__15_chanx_right_out[4] ,
    \cbx_1__1__15_chanx_right_out[5] ,
    \cbx_1__1__15_chanx_right_out[6] ,
    \cbx_1__1__15_chanx_right_out[7] ,
    \cbx_1__1__15_chanx_right_out[8] ,
    \cbx_1__1__15_chanx_right_out[9] ,
    \cbx_1__1__15_chanx_right_out[10] ,
    \cbx_1__1__15_chanx_right_out[11] ,
    \cbx_1__1__15_chanx_right_out[12] ,
    \cbx_1__1__15_chanx_right_out[13] ,
    \cbx_1__1__15_chanx_right_out[14] ,
    \cbx_1__1__15_chanx_right_out[15] ,
    \cbx_1__1__15_chanx_right_out[16] ,
    \cbx_1__1__15_chanx_right_out[17] ,
    \cbx_1__1__15_chanx_right_out[18] ,
    \cbx_1__1__15_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__15_chanx_left_out[0] ,
    \sb_1__1__15_chanx_left_out[1] ,
    \sb_1__1__15_chanx_left_out[2] ,
    \sb_1__1__15_chanx_left_out[3] ,
    \sb_1__1__15_chanx_left_out[4] ,
    \sb_1__1__15_chanx_left_out[5] ,
    \sb_1__1__15_chanx_left_out[6] ,
    \sb_1__1__15_chanx_left_out[7] ,
    \sb_1__1__15_chanx_left_out[8] ,
    \sb_1__1__15_chanx_left_out[9] ,
    \sb_1__1__15_chanx_left_out[10] ,
    \sb_1__1__15_chanx_left_out[11] ,
    \sb_1__1__15_chanx_left_out[12] ,
    \sb_1__1__15_chanx_left_out[13] ,
    \sb_1__1__15_chanx_left_out[14] ,
    \sb_1__1__15_chanx_left_out[15] ,
    \sb_1__1__15_chanx_left_out[16] ,
    \sb_1__1__15_chanx_left_out[17] ,
    \sb_1__1__15_chanx_left_out[18] ,
    \sb_1__1__15_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__22_chanx_left_out[0] ,
    \cbx_1__1__22_chanx_left_out[1] ,
    \cbx_1__1__22_chanx_left_out[2] ,
    \cbx_1__1__22_chanx_left_out[3] ,
    \cbx_1__1__22_chanx_left_out[4] ,
    \cbx_1__1__22_chanx_left_out[5] ,
    \cbx_1__1__22_chanx_left_out[6] ,
    \cbx_1__1__22_chanx_left_out[7] ,
    \cbx_1__1__22_chanx_left_out[8] ,
    \cbx_1__1__22_chanx_left_out[9] ,
    \cbx_1__1__22_chanx_left_out[10] ,
    \cbx_1__1__22_chanx_left_out[11] ,
    \cbx_1__1__22_chanx_left_out[12] ,
    \cbx_1__1__22_chanx_left_out[13] ,
    \cbx_1__1__22_chanx_left_out[14] ,
    \cbx_1__1__22_chanx_left_out[15] ,
    \cbx_1__1__22_chanx_left_out[16] ,
    \cbx_1__1__22_chanx_left_out[17] ,
    \cbx_1__1__22_chanx_left_out[18] ,
    \cbx_1__1__22_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__15_chanx_right_out[0] ,
    \sb_1__1__15_chanx_right_out[1] ,
    \sb_1__1__15_chanx_right_out[2] ,
    \sb_1__1__15_chanx_right_out[3] ,
    \sb_1__1__15_chanx_right_out[4] ,
    \sb_1__1__15_chanx_right_out[5] ,
    \sb_1__1__15_chanx_right_out[6] ,
    \sb_1__1__15_chanx_right_out[7] ,
    \sb_1__1__15_chanx_right_out[8] ,
    \sb_1__1__15_chanx_right_out[9] ,
    \sb_1__1__15_chanx_right_out[10] ,
    \sb_1__1__15_chanx_right_out[11] ,
    \sb_1__1__15_chanx_right_out[12] ,
    \sb_1__1__15_chanx_right_out[13] ,
    \sb_1__1__15_chanx_right_out[14] ,
    \sb_1__1__15_chanx_right_out[15] ,
    \sb_1__1__15_chanx_right_out[16] ,
    \sb_1__1__15_chanx_right_out[17] ,
    \sb_1__1__15_chanx_right_out[18] ,
    \sb_1__1__15_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__17_chany_top_out[0] ,
    \cby_1__1__17_chany_top_out[1] ,
    \cby_1__1__17_chany_top_out[2] ,
    \cby_1__1__17_chany_top_out[3] ,
    \cby_1__1__17_chany_top_out[4] ,
    \cby_1__1__17_chany_top_out[5] ,
    \cby_1__1__17_chany_top_out[6] ,
    \cby_1__1__17_chany_top_out[7] ,
    \cby_1__1__17_chany_top_out[8] ,
    \cby_1__1__17_chany_top_out[9] ,
    \cby_1__1__17_chany_top_out[10] ,
    \cby_1__1__17_chany_top_out[11] ,
    \cby_1__1__17_chany_top_out[12] ,
    \cby_1__1__17_chany_top_out[13] ,
    \cby_1__1__17_chany_top_out[14] ,
    \cby_1__1__17_chany_top_out[15] ,
    \cby_1__1__17_chany_top_out[16] ,
    \cby_1__1__17_chany_top_out[17] ,
    \cby_1__1__17_chany_top_out[18] ,
    \cby_1__1__17_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__15_chany_bottom_out[0] ,
    \sb_1__1__15_chany_bottom_out[1] ,
    \sb_1__1__15_chany_bottom_out[2] ,
    \sb_1__1__15_chany_bottom_out[3] ,
    \sb_1__1__15_chany_bottom_out[4] ,
    \sb_1__1__15_chany_bottom_out[5] ,
    \sb_1__1__15_chany_bottom_out[6] ,
    \sb_1__1__15_chany_bottom_out[7] ,
    \sb_1__1__15_chany_bottom_out[8] ,
    \sb_1__1__15_chany_bottom_out[9] ,
    \sb_1__1__15_chany_bottom_out[10] ,
    \sb_1__1__15_chany_bottom_out[11] ,
    \sb_1__1__15_chany_bottom_out[12] ,
    \sb_1__1__15_chany_bottom_out[13] ,
    \sb_1__1__15_chany_bottom_out[14] ,
    \sb_1__1__15_chany_bottom_out[15] ,
    \sb_1__1__15_chany_bottom_out[16] ,
    \sb_1__1__15_chany_bottom_out[17] ,
    \sb_1__1__15_chany_bottom_out[18] ,
    \sb_1__1__15_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__18_chany_bottom_out[0] ,
    \cby_1__1__18_chany_bottom_out[1] ,
    \cby_1__1__18_chany_bottom_out[2] ,
    \cby_1__1__18_chany_bottom_out[3] ,
    \cby_1__1__18_chany_bottom_out[4] ,
    \cby_1__1__18_chany_bottom_out[5] ,
    \cby_1__1__18_chany_bottom_out[6] ,
    \cby_1__1__18_chany_bottom_out[7] ,
    \cby_1__1__18_chany_bottom_out[8] ,
    \cby_1__1__18_chany_bottom_out[9] ,
    \cby_1__1__18_chany_bottom_out[10] ,
    \cby_1__1__18_chany_bottom_out[11] ,
    \cby_1__1__18_chany_bottom_out[12] ,
    \cby_1__1__18_chany_bottom_out[13] ,
    \cby_1__1__18_chany_bottom_out[14] ,
    \cby_1__1__18_chany_bottom_out[15] ,
    \cby_1__1__18_chany_bottom_out[16] ,
    \cby_1__1__18_chany_bottom_out[17] ,
    \cby_1__1__18_chany_bottom_out[18] ,
    \cby_1__1__18_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__15_chany_top_out[0] ,
    \sb_1__1__15_chany_top_out[1] ,
    \sb_1__1__15_chany_top_out[2] ,
    \sb_1__1__15_chany_top_out[3] ,
    \sb_1__1__15_chany_top_out[4] ,
    \sb_1__1__15_chany_top_out[5] ,
    \sb_1__1__15_chany_top_out[6] ,
    \sb_1__1__15_chany_top_out[7] ,
    \sb_1__1__15_chany_top_out[8] ,
    \sb_1__1__15_chany_top_out[9] ,
    \sb_1__1__15_chany_top_out[10] ,
    \sb_1__1__15_chany_top_out[11] ,
    \sb_1__1__15_chany_top_out[12] ,
    \sb_1__1__15_chany_top_out[13] ,
    \sb_1__1__15_chany_top_out[14] ,
    \sb_1__1__15_chany_top_out[15] ,
    \sb_1__1__15_chany_top_out[16] ,
    \sb_1__1__15_chany_top_out[17] ,
    \sb_1__1__15_chany_top_out[18] ,
    \sb_1__1__15_chany_top_out[19] }));
 sb_1__1_ sb_3__3_ (.bottom_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__23_ccff_tail),
    .ccff_tail(sb_1__1__16_ccff_tail),
    .clk_1_E_out(\clk_1_wires[36] ),
    .clk_1_N_in(\clk_2_wires[10] ),
    .clk_1_W_out(\clk_1_wires[37] ),
    .left_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[80] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[36] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[10] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[37] ),
    .right_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__16_chanx_right_out[0] ,
    \cbx_1__1__16_chanx_right_out[1] ,
    \cbx_1__1__16_chanx_right_out[2] ,
    \cbx_1__1__16_chanx_right_out[3] ,
    \cbx_1__1__16_chanx_right_out[4] ,
    \cbx_1__1__16_chanx_right_out[5] ,
    \cbx_1__1__16_chanx_right_out[6] ,
    \cbx_1__1__16_chanx_right_out[7] ,
    \cbx_1__1__16_chanx_right_out[8] ,
    \cbx_1__1__16_chanx_right_out[9] ,
    \cbx_1__1__16_chanx_right_out[10] ,
    \cbx_1__1__16_chanx_right_out[11] ,
    \cbx_1__1__16_chanx_right_out[12] ,
    \cbx_1__1__16_chanx_right_out[13] ,
    \cbx_1__1__16_chanx_right_out[14] ,
    \cbx_1__1__16_chanx_right_out[15] ,
    \cbx_1__1__16_chanx_right_out[16] ,
    \cbx_1__1__16_chanx_right_out[17] ,
    \cbx_1__1__16_chanx_right_out[18] ,
    \cbx_1__1__16_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__16_chanx_left_out[0] ,
    \sb_1__1__16_chanx_left_out[1] ,
    \sb_1__1__16_chanx_left_out[2] ,
    \sb_1__1__16_chanx_left_out[3] ,
    \sb_1__1__16_chanx_left_out[4] ,
    \sb_1__1__16_chanx_left_out[5] ,
    \sb_1__1__16_chanx_left_out[6] ,
    \sb_1__1__16_chanx_left_out[7] ,
    \sb_1__1__16_chanx_left_out[8] ,
    \sb_1__1__16_chanx_left_out[9] ,
    \sb_1__1__16_chanx_left_out[10] ,
    \sb_1__1__16_chanx_left_out[11] ,
    \sb_1__1__16_chanx_left_out[12] ,
    \sb_1__1__16_chanx_left_out[13] ,
    \sb_1__1__16_chanx_left_out[14] ,
    \sb_1__1__16_chanx_left_out[15] ,
    \sb_1__1__16_chanx_left_out[16] ,
    \sb_1__1__16_chanx_left_out[17] ,
    \sb_1__1__16_chanx_left_out[18] ,
    \sb_1__1__16_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__23_chanx_left_out[0] ,
    \cbx_1__1__23_chanx_left_out[1] ,
    \cbx_1__1__23_chanx_left_out[2] ,
    \cbx_1__1__23_chanx_left_out[3] ,
    \cbx_1__1__23_chanx_left_out[4] ,
    \cbx_1__1__23_chanx_left_out[5] ,
    \cbx_1__1__23_chanx_left_out[6] ,
    \cbx_1__1__23_chanx_left_out[7] ,
    \cbx_1__1__23_chanx_left_out[8] ,
    \cbx_1__1__23_chanx_left_out[9] ,
    \cbx_1__1__23_chanx_left_out[10] ,
    \cbx_1__1__23_chanx_left_out[11] ,
    \cbx_1__1__23_chanx_left_out[12] ,
    \cbx_1__1__23_chanx_left_out[13] ,
    \cbx_1__1__23_chanx_left_out[14] ,
    \cbx_1__1__23_chanx_left_out[15] ,
    \cbx_1__1__23_chanx_left_out[16] ,
    \cbx_1__1__23_chanx_left_out[17] ,
    \cbx_1__1__23_chanx_left_out[18] ,
    \cbx_1__1__23_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__16_chanx_right_out[0] ,
    \sb_1__1__16_chanx_right_out[1] ,
    \sb_1__1__16_chanx_right_out[2] ,
    \sb_1__1__16_chanx_right_out[3] ,
    \sb_1__1__16_chanx_right_out[4] ,
    \sb_1__1__16_chanx_right_out[5] ,
    \sb_1__1__16_chanx_right_out[6] ,
    \sb_1__1__16_chanx_right_out[7] ,
    \sb_1__1__16_chanx_right_out[8] ,
    \sb_1__1__16_chanx_right_out[9] ,
    \sb_1__1__16_chanx_right_out[10] ,
    \sb_1__1__16_chanx_right_out[11] ,
    \sb_1__1__16_chanx_right_out[12] ,
    \sb_1__1__16_chanx_right_out[13] ,
    \sb_1__1__16_chanx_right_out[14] ,
    \sb_1__1__16_chanx_right_out[15] ,
    \sb_1__1__16_chanx_right_out[16] ,
    \sb_1__1__16_chanx_right_out[17] ,
    \sb_1__1__16_chanx_right_out[18] ,
    \sb_1__1__16_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__18_chany_top_out[0] ,
    \cby_1__1__18_chany_top_out[1] ,
    \cby_1__1__18_chany_top_out[2] ,
    \cby_1__1__18_chany_top_out[3] ,
    \cby_1__1__18_chany_top_out[4] ,
    \cby_1__1__18_chany_top_out[5] ,
    \cby_1__1__18_chany_top_out[6] ,
    \cby_1__1__18_chany_top_out[7] ,
    \cby_1__1__18_chany_top_out[8] ,
    \cby_1__1__18_chany_top_out[9] ,
    \cby_1__1__18_chany_top_out[10] ,
    \cby_1__1__18_chany_top_out[11] ,
    \cby_1__1__18_chany_top_out[12] ,
    \cby_1__1__18_chany_top_out[13] ,
    \cby_1__1__18_chany_top_out[14] ,
    \cby_1__1__18_chany_top_out[15] ,
    \cby_1__1__18_chany_top_out[16] ,
    \cby_1__1__18_chany_top_out[17] ,
    \cby_1__1__18_chany_top_out[18] ,
    \cby_1__1__18_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__16_chany_bottom_out[0] ,
    \sb_1__1__16_chany_bottom_out[1] ,
    \sb_1__1__16_chany_bottom_out[2] ,
    \sb_1__1__16_chany_bottom_out[3] ,
    \sb_1__1__16_chany_bottom_out[4] ,
    \sb_1__1__16_chany_bottom_out[5] ,
    \sb_1__1__16_chany_bottom_out[6] ,
    \sb_1__1__16_chany_bottom_out[7] ,
    \sb_1__1__16_chany_bottom_out[8] ,
    \sb_1__1__16_chany_bottom_out[9] ,
    \sb_1__1__16_chany_bottom_out[10] ,
    \sb_1__1__16_chany_bottom_out[11] ,
    \sb_1__1__16_chany_bottom_out[12] ,
    \sb_1__1__16_chany_bottom_out[13] ,
    \sb_1__1__16_chany_bottom_out[14] ,
    \sb_1__1__16_chany_bottom_out[15] ,
    \sb_1__1__16_chany_bottom_out[16] ,
    \sb_1__1__16_chany_bottom_out[17] ,
    \sb_1__1__16_chany_bottom_out[18] ,
    \sb_1__1__16_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__19_chany_bottom_out[0] ,
    \cby_1__1__19_chany_bottom_out[1] ,
    \cby_1__1__19_chany_bottom_out[2] ,
    \cby_1__1__19_chany_bottom_out[3] ,
    \cby_1__1__19_chany_bottom_out[4] ,
    \cby_1__1__19_chany_bottom_out[5] ,
    \cby_1__1__19_chany_bottom_out[6] ,
    \cby_1__1__19_chany_bottom_out[7] ,
    \cby_1__1__19_chany_bottom_out[8] ,
    \cby_1__1__19_chany_bottom_out[9] ,
    \cby_1__1__19_chany_bottom_out[10] ,
    \cby_1__1__19_chany_bottom_out[11] ,
    \cby_1__1__19_chany_bottom_out[12] ,
    \cby_1__1__19_chany_bottom_out[13] ,
    \cby_1__1__19_chany_bottom_out[14] ,
    \cby_1__1__19_chany_bottom_out[15] ,
    \cby_1__1__19_chany_bottom_out[16] ,
    \cby_1__1__19_chany_bottom_out[17] ,
    \cby_1__1__19_chany_bottom_out[18] ,
    \cby_1__1__19_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__16_chany_top_out[0] ,
    \sb_1__1__16_chany_top_out[1] ,
    \sb_1__1__16_chany_top_out[2] ,
    \sb_1__1__16_chany_top_out[3] ,
    \sb_1__1__16_chany_top_out[4] ,
    \sb_1__1__16_chany_top_out[5] ,
    \sb_1__1__16_chany_top_out[6] ,
    \sb_1__1__16_chany_top_out[7] ,
    \sb_1__1__16_chany_top_out[8] ,
    \sb_1__1__16_chany_top_out[9] ,
    \sb_1__1__16_chany_top_out[10] ,
    \sb_1__1__16_chany_top_out[11] ,
    \sb_1__1__16_chany_top_out[12] ,
    \sb_1__1__16_chany_top_out[13] ,
    \sb_1__1__16_chany_top_out[14] ,
    \sb_1__1__16_chany_top_out[15] ,
    \sb_1__1__16_chany_top_out[16] ,
    \sb_1__1__16_chany_top_out[17] ,
    \sb_1__1__16_chany_top_out[18] ,
    \sb_1__1__16_chany_top_out[19] }));
 sb_1__1_ sb_3__4_ (.bottom_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__24_ccff_tail),
    .ccff_tail(sb_1__1__17_ccff_tail),
    .clk_3_N_in(\clk_3_wires[4] ),
    .clk_3_W_out(\clk_3_wires[8] ),
    .left_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[83] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[4] ),
    .prog_clk_3_W_out(\prog_clk_3_wires[8] ),
    .right_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__17_chanx_right_out[0] ,
    \cbx_1__1__17_chanx_right_out[1] ,
    \cbx_1__1__17_chanx_right_out[2] ,
    \cbx_1__1__17_chanx_right_out[3] ,
    \cbx_1__1__17_chanx_right_out[4] ,
    \cbx_1__1__17_chanx_right_out[5] ,
    \cbx_1__1__17_chanx_right_out[6] ,
    \cbx_1__1__17_chanx_right_out[7] ,
    \cbx_1__1__17_chanx_right_out[8] ,
    \cbx_1__1__17_chanx_right_out[9] ,
    \cbx_1__1__17_chanx_right_out[10] ,
    \cbx_1__1__17_chanx_right_out[11] ,
    \cbx_1__1__17_chanx_right_out[12] ,
    \cbx_1__1__17_chanx_right_out[13] ,
    \cbx_1__1__17_chanx_right_out[14] ,
    \cbx_1__1__17_chanx_right_out[15] ,
    \cbx_1__1__17_chanx_right_out[16] ,
    \cbx_1__1__17_chanx_right_out[17] ,
    \cbx_1__1__17_chanx_right_out[18] ,
    \cbx_1__1__17_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__17_chanx_left_out[0] ,
    \sb_1__1__17_chanx_left_out[1] ,
    \sb_1__1__17_chanx_left_out[2] ,
    \sb_1__1__17_chanx_left_out[3] ,
    \sb_1__1__17_chanx_left_out[4] ,
    \sb_1__1__17_chanx_left_out[5] ,
    \sb_1__1__17_chanx_left_out[6] ,
    \sb_1__1__17_chanx_left_out[7] ,
    \sb_1__1__17_chanx_left_out[8] ,
    \sb_1__1__17_chanx_left_out[9] ,
    \sb_1__1__17_chanx_left_out[10] ,
    \sb_1__1__17_chanx_left_out[11] ,
    \sb_1__1__17_chanx_left_out[12] ,
    \sb_1__1__17_chanx_left_out[13] ,
    \sb_1__1__17_chanx_left_out[14] ,
    \sb_1__1__17_chanx_left_out[15] ,
    \sb_1__1__17_chanx_left_out[16] ,
    \sb_1__1__17_chanx_left_out[17] ,
    \sb_1__1__17_chanx_left_out[18] ,
    \sb_1__1__17_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__24_chanx_left_out[0] ,
    \cbx_1__1__24_chanx_left_out[1] ,
    \cbx_1__1__24_chanx_left_out[2] ,
    \cbx_1__1__24_chanx_left_out[3] ,
    \cbx_1__1__24_chanx_left_out[4] ,
    \cbx_1__1__24_chanx_left_out[5] ,
    \cbx_1__1__24_chanx_left_out[6] ,
    \cbx_1__1__24_chanx_left_out[7] ,
    \cbx_1__1__24_chanx_left_out[8] ,
    \cbx_1__1__24_chanx_left_out[9] ,
    \cbx_1__1__24_chanx_left_out[10] ,
    \cbx_1__1__24_chanx_left_out[11] ,
    \cbx_1__1__24_chanx_left_out[12] ,
    \cbx_1__1__24_chanx_left_out[13] ,
    \cbx_1__1__24_chanx_left_out[14] ,
    \cbx_1__1__24_chanx_left_out[15] ,
    \cbx_1__1__24_chanx_left_out[16] ,
    \cbx_1__1__24_chanx_left_out[17] ,
    \cbx_1__1__24_chanx_left_out[18] ,
    \cbx_1__1__24_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__17_chanx_right_out[0] ,
    \sb_1__1__17_chanx_right_out[1] ,
    \sb_1__1__17_chanx_right_out[2] ,
    \sb_1__1__17_chanx_right_out[3] ,
    \sb_1__1__17_chanx_right_out[4] ,
    \sb_1__1__17_chanx_right_out[5] ,
    \sb_1__1__17_chanx_right_out[6] ,
    \sb_1__1__17_chanx_right_out[7] ,
    \sb_1__1__17_chanx_right_out[8] ,
    \sb_1__1__17_chanx_right_out[9] ,
    \sb_1__1__17_chanx_right_out[10] ,
    \sb_1__1__17_chanx_right_out[11] ,
    \sb_1__1__17_chanx_right_out[12] ,
    \sb_1__1__17_chanx_right_out[13] ,
    \sb_1__1__17_chanx_right_out[14] ,
    \sb_1__1__17_chanx_right_out[15] ,
    \sb_1__1__17_chanx_right_out[16] ,
    \sb_1__1__17_chanx_right_out[17] ,
    \sb_1__1__17_chanx_right_out[18] ,
    \sb_1__1__17_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__19_chany_top_out[0] ,
    \cby_1__1__19_chany_top_out[1] ,
    \cby_1__1__19_chany_top_out[2] ,
    \cby_1__1__19_chany_top_out[3] ,
    \cby_1__1__19_chany_top_out[4] ,
    \cby_1__1__19_chany_top_out[5] ,
    \cby_1__1__19_chany_top_out[6] ,
    \cby_1__1__19_chany_top_out[7] ,
    \cby_1__1__19_chany_top_out[8] ,
    \cby_1__1__19_chany_top_out[9] ,
    \cby_1__1__19_chany_top_out[10] ,
    \cby_1__1__19_chany_top_out[11] ,
    \cby_1__1__19_chany_top_out[12] ,
    \cby_1__1__19_chany_top_out[13] ,
    \cby_1__1__19_chany_top_out[14] ,
    \cby_1__1__19_chany_top_out[15] ,
    \cby_1__1__19_chany_top_out[16] ,
    \cby_1__1__19_chany_top_out[17] ,
    \cby_1__1__19_chany_top_out[18] ,
    \cby_1__1__19_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__17_chany_bottom_out[0] ,
    \sb_1__1__17_chany_bottom_out[1] ,
    \sb_1__1__17_chany_bottom_out[2] ,
    \sb_1__1__17_chany_bottom_out[3] ,
    \sb_1__1__17_chany_bottom_out[4] ,
    \sb_1__1__17_chany_bottom_out[5] ,
    \sb_1__1__17_chany_bottom_out[6] ,
    \sb_1__1__17_chany_bottom_out[7] ,
    \sb_1__1__17_chany_bottom_out[8] ,
    \sb_1__1__17_chany_bottom_out[9] ,
    \sb_1__1__17_chany_bottom_out[10] ,
    \sb_1__1__17_chany_bottom_out[11] ,
    \sb_1__1__17_chany_bottom_out[12] ,
    \sb_1__1__17_chany_bottom_out[13] ,
    \sb_1__1__17_chany_bottom_out[14] ,
    \sb_1__1__17_chany_bottom_out[15] ,
    \sb_1__1__17_chany_bottom_out[16] ,
    \sb_1__1__17_chany_bottom_out[17] ,
    \sb_1__1__17_chany_bottom_out[18] ,
    \sb_1__1__17_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__20_chany_bottom_out[0] ,
    \cby_1__1__20_chany_bottom_out[1] ,
    \cby_1__1__20_chany_bottom_out[2] ,
    \cby_1__1__20_chany_bottom_out[3] ,
    \cby_1__1__20_chany_bottom_out[4] ,
    \cby_1__1__20_chany_bottom_out[5] ,
    \cby_1__1__20_chany_bottom_out[6] ,
    \cby_1__1__20_chany_bottom_out[7] ,
    \cby_1__1__20_chany_bottom_out[8] ,
    \cby_1__1__20_chany_bottom_out[9] ,
    \cby_1__1__20_chany_bottom_out[10] ,
    \cby_1__1__20_chany_bottom_out[11] ,
    \cby_1__1__20_chany_bottom_out[12] ,
    \cby_1__1__20_chany_bottom_out[13] ,
    \cby_1__1__20_chany_bottom_out[14] ,
    \cby_1__1__20_chany_bottom_out[15] ,
    \cby_1__1__20_chany_bottom_out[16] ,
    \cby_1__1__20_chany_bottom_out[17] ,
    \cby_1__1__20_chany_bottom_out[18] ,
    \cby_1__1__20_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__17_chany_top_out[0] ,
    \sb_1__1__17_chany_top_out[1] ,
    \sb_1__1__17_chany_top_out[2] ,
    \sb_1__1__17_chany_top_out[3] ,
    \sb_1__1__17_chany_top_out[4] ,
    \sb_1__1__17_chany_top_out[5] ,
    \sb_1__1__17_chany_top_out[6] ,
    \sb_1__1__17_chany_top_out[7] ,
    \sb_1__1__17_chany_top_out[8] ,
    \sb_1__1__17_chany_top_out[9] ,
    \sb_1__1__17_chany_top_out[10] ,
    \sb_1__1__17_chany_top_out[11] ,
    \sb_1__1__17_chany_top_out[12] ,
    \sb_1__1__17_chany_top_out[13] ,
    \sb_1__1__17_chany_top_out[14] ,
    \sb_1__1__17_chany_top_out[15] ,
    \sb_1__1__17_chany_top_out[16] ,
    \sb_1__1__17_chany_top_out[17] ,
    \sb_1__1__17_chany_top_out[18] ,
    \sb_1__1__17_chany_top_out[19] }));
 sb_1__1_ sb_3__5_ (.bottom_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__25_ccff_tail),
    .ccff_tail(sb_1__1__18_ccff_tail),
    .clk_1_E_out(\clk_1_wires[43] ),
    .clk_1_N_in(\clk_2_wires[25] ),
    .clk_1_W_out(\clk_1_wires[44] ),
    .left_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[86] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[43] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[25] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[44] ),
    .right_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__18_chanx_right_out[0] ,
    \cbx_1__1__18_chanx_right_out[1] ,
    \cbx_1__1__18_chanx_right_out[2] ,
    \cbx_1__1__18_chanx_right_out[3] ,
    \cbx_1__1__18_chanx_right_out[4] ,
    \cbx_1__1__18_chanx_right_out[5] ,
    \cbx_1__1__18_chanx_right_out[6] ,
    \cbx_1__1__18_chanx_right_out[7] ,
    \cbx_1__1__18_chanx_right_out[8] ,
    \cbx_1__1__18_chanx_right_out[9] ,
    \cbx_1__1__18_chanx_right_out[10] ,
    \cbx_1__1__18_chanx_right_out[11] ,
    \cbx_1__1__18_chanx_right_out[12] ,
    \cbx_1__1__18_chanx_right_out[13] ,
    \cbx_1__1__18_chanx_right_out[14] ,
    \cbx_1__1__18_chanx_right_out[15] ,
    \cbx_1__1__18_chanx_right_out[16] ,
    \cbx_1__1__18_chanx_right_out[17] ,
    \cbx_1__1__18_chanx_right_out[18] ,
    \cbx_1__1__18_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__18_chanx_left_out[0] ,
    \sb_1__1__18_chanx_left_out[1] ,
    \sb_1__1__18_chanx_left_out[2] ,
    \sb_1__1__18_chanx_left_out[3] ,
    \sb_1__1__18_chanx_left_out[4] ,
    \sb_1__1__18_chanx_left_out[5] ,
    \sb_1__1__18_chanx_left_out[6] ,
    \sb_1__1__18_chanx_left_out[7] ,
    \sb_1__1__18_chanx_left_out[8] ,
    \sb_1__1__18_chanx_left_out[9] ,
    \sb_1__1__18_chanx_left_out[10] ,
    \sb_1__1__18_chanx_left_out[11] ,
    \sb_1__1__18_chanx_left_out[12] ,
    \sb_1__1__18_chanx_left_out[13] ,
    \sb_1__1__18_chanx_left_out[14] ,
    \sb_1__1__18_chanx_left_out[15] ,
    \sb_1__1__18_chanx_left_out[16] ,
    \sb_1__1__18_chanx_left_out[17] ,
    \sb_1__1__18_chanx_left_out[18] ,
    \sb_1__1__18_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__25_chanx_left_out[0] ,
    \cbx_1__1__25_chanx_left_out[1] ,
    \cbx_1__1__25_chanx_left_out[2] ,
    \cbx_1__1__25_chanx_left_out[3] ,
    \cbx_1__1__25_chanx_left_out[4] ,
    \cbx_1__1__25_chanx_left_out[5] ,
    \cbx_1__1__25_chanx_left_out[6] ,
    \cbx_1__1__25_chanx_left_out[7] ,
    \cbx_1__1__25_chanx_left_out[8] ,
    \cbx_1__1__25_chanx_left_out[9] ,
    \cbx_1__1__25_chanx_left_out[10] ,
    \cbx_1__1__25_chanx_left_out[11] ,
    \cbx_1__1__25_chanx_left_out[12] ,
    \cbx_1__1__25_chanx_left_out[13] ,
    \cbx_1__1__25_chanx_left_out[14] ,
    \cbx_1__1__25_chanx_left_out[15] ,
    \cbx_1__1__25_chanx_left_out[16] ,
    \cbx_1__1__25_chanx_left_out[17] ,
    \cbx_1__1__25_chanx_left_out[18] ,
    \cbx_1__1__25_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__18_chanx_right_out[0] ,
    \sb_1__1__18_chanx_right_out[1] ,
    \sb_1__1__18_chanx_right_out[2] ,
    \sb_1__1__18_chanx_right_out[3] ,
    \sb_1__1__18_chanx_right_out[4] ,
    \sb_1__1__18_chanx_right_out[5] ,
    \sb_1__1__18_chanx_right_out[6] ,
    \sb_1__1__18_chanx_right_out[7] ,
    \sb_1__1__18_chanx_right_out[8] ,
    \sb_1__1__18_chanx_right_out[9] ,
    \sb_1__1__18_chanx_right_out[10] ,
    \sb_1__1__18_chanx_right_out[11] ,
    \sb_1__1__18_chanx_right_out[12] ,
    \sb_1__1__18_chanx_right_out[13] ,
    \sb_1__1__18_chanx_right_out[14] ,
    \sb_1__1__18_chanx_right_out[15] ,
    \sb_1__1__18_chanx_right_out[16] ,
    \sb_1__1__18_chanx_right_out[17] ,
    \sb_1__1__18_chanx_right_out[18] ,
    \sb_1__1__18_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__20_chany_top_out[0] ,
    \cby_1__1__20_chany_top_out[1] ,
    \cby_1__1__20_chany_top_out[2] ,
    \cby_1__1__20_chany_top_out[3] ,
    \cby_1__1__20_chany_top_out[4] ,
    \cby_1__1__20_chany_top_out[5] ,
    \cby_1__1__20_chany_top_out[6] ,
    \cby_1__1__20_chany_top_out[7] ,
    \cby_1__1__20_chany_top_out[8] ,
    \cby_1__1__20_chany_top_out[9] ,
    \cby_1__1__20_chany_top_out[10] ,
    \cby_1__1__20_chany_top_out[11] ,
    \cby_1__1__20_chany_top_out[12] ,
    \cby_1__1__20_chany_top_out[13] ,
    \cby_1__1__20_chany_top_out[14] ,
    \cby_1__1__20_chany_top_out[15] ,
    \cby_1__1__20_chany_top_out[16] ,
    \cby_1__1__20_chany_top_out[17] ,
    \cby_1__1__20_chany_top_out[18] ,
    \cby_1__1__20_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__18_chany_bottom_out[0] ,
    \sb_1__1__18_chany_bottom_out[1] ,
    \sb_1__1__18_chany_bottom_out[2] ,
    \sb_1__1__18_chany_bottom_out[3] ,
    \sb_1__1__18_chany_bottom_out[4] ,
    \sb_1__1__18_chany_bottom_out[5] ,
    \sb_1__1__18_chany_bottom_out[6] ,
    \sb_1__1__18_chany_bottom_out[7] ,
    \sb_1__1__18_chany_bottom_out[8] ,
    \sb_1__1__18_chany_bottom_out[9] ,
    \sb_1__1__18_chany_bottom_out[10] ,
    \sb_1__1__18_chany_bottom_out[11] ,
    \sb_1__1__18_chany_bottom_out[12] ,
    \sb_1__1__18_chany_bottom_out[13] ,
    \sb_1__1__18_chany_bottom_out[14] ,
    \sb_1__1__18_chany_bottom_out[15] ,
    \sb_1__1__18_chany_bottom_out[16] ,
    \sb_1__1__18_chany_bottom_out[17] ,
    \sb_1__1__18_chany_bottom_out[18] ,
    \sb_1__1__18_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__21_chany_bottom_out[0] ,
    \cby_1__1__21_chany_bottom_out[1] ,
    \cby_1__1__21_chany_bottom_out[2] ,
    \cby_1__1__21_chany_bottom_out[3] ,
    \cby_1__1__21_chany_bottom_out[4] ,
    \cby_1__1__21_chany_bottom_out[5] ,
    \cby_1__1__21_chany_bottom_out[6] ,
    \cby_1__1__21_chany_bottom_out[7] ,
    \cby_1__1__21_chany_bottom_out[8] ,
    \cby_1__1__21_chany_bottom_out[9] ,
    \cby_1__1__21_chany_bottom_out[10] ,
    \cby_1__1__21_chany_bottom_out[11] ,
    \cby_1__1__21_chany_bottom_out[12] ,
    \cby_1__1__21_chany_bottom_out[13] ,
    \cby_1__1__21_chany_bottom_out[14] ,
    \cby_1__1__21_chany_bottom_out[15] ,
    \cby_1__1__21_chany_bottom_out[16] ,
    \cby_1__1__21_chany_bottom_out[17] ,
    \cby_1__1__21_chany_bottom_out[18] ,
    \cby_1__1__21_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__18_chany_top_out[0] ,
    \sb_1__1__18_chany_top_out[1] ,
    \sb_1__1__18_chany_top_out[2] ,
    \sb_1__1__18_chany_top_out[3] ,
    \sb_1__1__18_chany_top_out[4] ,
    \sb_1__1__18_chany_top_out[5] ,
    \sb_1__1__18_chany_top_out[6] ,
    \sb_1__1__18_chany_top_out[7] ,
    \sb_1__1__18_chany_top_out[8] ,
    \sb_1__1__18_chany_top_out[9] ,
    \sb_1__1__18_chany_top_out[10] ,
    \sb_1__1__18_chany_top_out[11] ,
    \sb_1__1__18_chany_top_out[12] ,
    \sb_1__1__18_chany_top_out[13] ,
    \sb_1__1__18_chany_top_out[14] ,
    \sb_1__1__18_chany_top_out[15] ,
    \sb_1__1__18_chany_top_out[16] ,
    \sb_1__1__18_chany_top_out[17] ,
    \sb_1__1__18_chany_top_out[18] ,
    \sb_1__1__18_chany_top_out[19] }));
 sb_1__1_ sb_3__6_ (.bottom_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__26_ccff_tail),
    .ccff_tail(sb_1__1__19_ccff_tail),
    .clk_2_N_in(\clk_2_wires[15] ),
    .clk_2_N_out(\clk_2_wires[22] ),
    .clk_2_S_out(\clk_2_wires[24] ),
    .left_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[89] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[15] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[22] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[24] ),
    .right_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__19_chanx_right_out[0] ,
    \cbx_1__1__19_chanx_right_out[1] ,
    \cbx_1__1__19_chanx_right_out[2] ,
    \cbx_1__1__19_chanx_right_out[3] ,
    \cbx_1__1__19_chanx_right_out[4] ,
    \cbx_1__1__19_chanx_right_out[5] ,
    \cbx_1__1__19_chanx_right_out[6] ,
    \cbx_1__1__19_chanx_right_out[7] ,
    \cbx_1__1__19_chanx_right_out[8] ,
    \cbx_1__1__19_chanx_right_out[9] ,
    \cbx_1__1__19_chanx_right_out[10] ,
    \cbx_1__1__19_chanx_right_out[11] ,
    \cbx_1__1__19_chanx_right_out[12] ,
    \cbx_1__1__19_chanx_right_out[13] ,
    \cbx_1__1__19_chanx_right_out[14] ,
    \cbx_1__1__19_chanx_right_out[15] ,
    \cbx_1__1__19_chanx_right_out[16] ,
    \cbx_1__1__19_chanx_right_out[17] ,
    \cbx_1__1__19_chanx_right_out[18] ,
    \cbx_1__1__19_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__19_chanx_left_out[0] ,
    \sb_1__1__19_chanx_left_out[1] ,
    \sb_1__1__19_chanx_left_out[2] ,
    \sb_1__1__19_chanx_left_out[3] ,
    \sb_1__1__19_chanx_left_out[4] ,
    \sb_1__1__19_chanx_left_out[5] ,
    \sb_1__1__19_chanx_left_out[6] ,
    \sb_1__1__19_chanx_left_out[7] ,
    \sb_1__1__19_chanx_left_out[8] ,
    \sb_1__1__19_chanx_left_out[9] ,
    \sb_1__1__19_chanx_left_out[10] ,
    \sb_1__1__19_chanx_left_out[11] ,
    \sb_1__1__19_chanx_left_out[12] ,
    \sb_1__1__19_chanx_left_out[13] ,
    \sb_1__1__19_chanx_left_out[14] ,
    \sb_1__1__19_chanx_left_out[15] ,
    \sb_1__1__19_chanx_left_out[16] ,
    \sb_1__1__19_chanx_left_out[17] ,
    \sb_1__1__19_chanx_left_out[18] ,
    \sb_1__1__19_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__26_chanx_left_out[0] ,
    \cbx_1__1__26_chanx_left_out[1] ,
    \cbx_1__1__26_chanx_left_out[2] ,
    \cbx_1__1__26_chanx_left_out[3] ,
    \cbx_1__1__26_chanx_left_out[4] ,
    \cbx_1__1__26_chanx_left_out[5] ,
    \cbx_1__1__26_chanx_left_out[6] ,
    \cbx_1__1__26_chanx_left_out[7] ,
    \cbx_1__1__26_chanx_left_out[8] ,
    \cbx_1__1__26_chanx_left_out[9] ,
    \cbx_1__1__26_chanx_left_out[10] ,
    \cbx_1__1__26_chanx_left_out[11] ,
    \cbx_1__1__26_chanx_left_out[12] ,
    \cbx_1__1__26_chanx_left_out[13] ,
    \cbx_1__1__26_chanx_left_out[14] ,
    \cbx_1__1__26_chanx_left_out[15] ,
    \cbx_1__1__26_chanx_left_out[16] ,
    \cbx_1__1__26_chanx_left_out[17] ,
    \cbx_1__1__26_chanx_left_out[18] ,
    \cbx_1__1__26_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__19_chanx_right_out[0] ,
    \sb_1__1__19_chanx_right_out[1] ,
    \sb_1__1__19_chanx_right_out[2] ,
    \sb_1__1__19_chanx_right_out[3] ,
    \sb_1__1__19_chanx_right_out[4] ,
    \sb_1__1__19_chanx_right_out[5] ,
    \sb_1__1__19_chanx_right_out[6] ,
    \sb_1__1__19_chanx_right_out[7] ,
    \sb_1__1__19_chanx_right_out[8] ,
    \sb_1__1__19_chanx_right_out[9] ,
    \sb_1__1__19_chanx_right_out[10] ,
    \sb_1__1__19_chanx_right_out[11] ,
    \sb_1__1__19_chanx_right_out[12] ,
    \sb_1__1__19_chanx_right_out[13] ,
    \sb_1__1__19_chanx_right_out[14] ,
    \sb_1__1__19_chanx_right_out[15] ,
    \sb_1__1__19_chanx_right_out[16] ,
    \sb_1__1__19_chanx_right_out[17] ,
    \sb_1__1__19_chanx_right_out[18] ,
    \sb_1__1__19_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__21_chany_top_out[0] ,
    \cby_1__1__21_chany_top_out[1] ,
    \cby_1__1__21_chany_top_out[2] ,
    \cby_1__1__21_chany_top_out[3] ,
    \cby_1__1__21_chany_top_out[4] ,
    \cby_1__1__21_chany_top_out[5] ,
    \cby_1__1__21_chany_top_out[6] ,
    \cby_1__1__21_chany_top_out[7] ,
    \cby_1__1__21_chany_top_out[8] ,
    \cby_1__1__21_chany_top_out[9] ,
    \cby_1__1__21_chany_top_out[10] ,
    \cby_1__1__21_chany_top_out[11] ,
    \cby_1__1__21_chany_top_out[12] ,
    \cby_1__1__21_chany_top_out[13] ,
    \cby_1__1__21_chany_top_out[14] ,
    \cby_1__1__21_chany_top_out[15] ,
    \cby_1__1__21_chany_top_out[16] ,
    \cby_1__1__21_chany_top_out[17] ,
    \cby_1__1__21_chany_top_out[18] ,
    \cby_1__1__21_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__19_chany_bottom_out[0] ,
    \sb_1__1__19_chany_bottom_out[1] ,
    \sb_1__1__19_chany_bottom_out[2] ,
    \sb_1__1__19_chany_bottom_out[3] ,
    \sb_1__1__19_chany_bottom_out[4] ,
    \sb_1__1__19_chany_bottom_out[5] ,
    \sb_1__1__19_chany_bottom_out[6] ,
    \sb_1__1__19_chany_bottom_out[7] ,
    \sb_1__1__19_chany_bottom_out[8] ,
    \sb_1__1__19_chany_bottom_out[9] ,
    \sb_1__1__19_chany_bottom_out[10] ,
    \sb_1__1__19_chany_bottom_out[11] ,
    \sb_1__1__19_chany_bottom_out[12] ,
    \sb_1__1__19_chany_bottom_out[13] ,
    \sb_1__1__19_chany_bottom_out[14] ,
    \sb_1__1__19_chany_bottom_out[15] ,
    \sb_1__1__19_chany_bottom_out[16] ,
    \sb_1__1__19_chany_bottom_out[17] ,
    \sb_1__1__19_chany_bottom_out[18] ,
    \sb_1__1__19_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__22_chany_bottom_out[0] ,
    \cby_1__1__22_chany_bottom_out[1] ,
    \cby_1__1__22_chany_bottom_out[2] ,
    \cby_1__1__22_chany_bottom_out[3] ,
    \cby_1__1__22_chany_bottom_out[4] ,
    \cby_1__1__22_chany_bottom_out[5] ,
    \cby_1__1__22_chany_bottom_out[6] ,
    \cby_1__1__22_chany_bottom_out[7] ,
    \cby_1__1__22_chany_bottom_out[8] ,
    \cby_1__1__22_chany_bottom_out[9] ,
    \cby_1__1__22_chany_bottom_out[10] ,
    \cby_1__1__22_chany_bottom_out[11] ,
    \cby_1__1__22_chany_bottom_out[12] ,
    \cby_1__1__22_chany_bottom_out[13] ,
    \cby_1__1__22_chany_bottom_out[14] ,
    \cby_1__1__22_chany_bottom_out[15] ,
    \cby_1__1__22_chany_bottom_out[16] ,
    \cby_1__1__22_chany_bottom_out[17] ,
    \cby_1__1__22_chany_bottom_out[18] ,
    \cby_1__1__22_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__19_chany_top_out[0] ,
    \sb_1__1__19_chany_top_out[1] ,
    \sb_1__1__19_chany_top_out[2] ,
    \sb_1__1__19_chany_top_out[3] ,
    \sb_1__1__19_chany_top_out[4] ,
    \sb_1__1__19_chany_top_out[5] ,
    \sb_1__1__19_chany_top_out[6] ,
    \sb_1__1__19_chany_top_out[7] ,
    \sb_1__1__19_chany_top_out[8] ,
    \sb_1__1__19_chany_top_out[9] ,
    \sb_1__1__19_chany_top_out[10] ,
    \sb_1__1__19_chany_top_out[11] ,
    \sb_1__1__19_chany_top_out[12] ,
    \sb_1__1__19_chany_top_out[13] ,
    \sb_1__1__19_chany_top_out[14] ,
    \sb_1__1__19_chany_top_out[15] ,
    \sb_1__1__19_chany_top_out[16] ,
    \sb_1__1__19_chany_top_out[17] ,
    \sb_1__1__19_chany_top_out[18] ,
    \sb_1__1__19_chany_top_out[19] }));
 sb_1__1_ sb_3__7_ (.bottom_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__27_ccff_tail),
    .ccff_tail(sb_1__1__20_ccff_tail),
    .clk_1_E_out(\clk_1_wires[50] ),
    .clk_1_N_in(\clk_2_wires[23] ),
    .clk_1_W_out(\clk_1_wires[51] ),
    .left_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[92] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[50] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[23] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[51] ),
    .right_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__20_chanx_right_out[0] ,
    \cbx_1__1__20_chanx_right_out[1] ,
    \cbx_1__1__20_chanx_right_out[2] ,
    \cbx_1__1__20_chanx_right_out[3] ,
    \cbx_1__1__20_chanx_right_out[4] ,
    \cbx_1__1__20_chanx_right_out[5] ,
    \cbx_1__1__20_chanx_right_out[6] ,
    \cbx_1__1__20_chanx_right_out[7] ,
    \cbx_1__1__20_chanx_right_out[8] ,
    \cbx_1__1__20_chanx_right_out[9] ,
    \cbx_1__1__20_chanx_right_out[10] ,
    \cbx_1__1__20_chanx_right_out[11] ,
    \cbx_1__1__20_chanx_right_out[12] ,
    \cbx_1__1__20_chanx_right_out[13] ,
    \cbx_1__1__20_chanx_right_out[14] ,
    \cbx_1__1__20_chanx_right_out[15] ,
    \cbx_1__1__20_chanx_right_out[16] ,
    \cbx_1__1__20_chanx_right_out[17] ,
    \cbx_1__1__20_chanx_right_out[18] ,
    \cbx_1__1__20_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__20_chanx_left_out[0] ,
    \sb_1__1__20_chanx_left_out[1] ,
    \sb_1__1__20_chanx_left_out[2] ,
    \sb_1__1__20_chanx_left_out[3] ,
    \sb_1__1__20_chanx_left_out[4] ,
    \sb_1__1__20_chanx_left_out[5] ,
    \sb_1__1__20_chanx_left_out[6] ,
    \sb_1__1__20_chanx_left_out[7] ,
    \sb_1__1__20_chanx_left_out[8] ,
    \sb_1__1__20_chanx_left_out[9] ,
    \sb_1__1__20_chanx_left_out[10] ,
    \sb_1__1__20_chanx_left_out[11] ,
    \sb_1__1__20_chanx_left_out[12] ,
    \sb_1__1__20_chanx_left_out[13] ,
    \sb_1__1__20_chanx_left_out[14] ,
    \sb_1__1__20_chanx_left_out[15] ,
    \sb_1__1__20_chanx_left_out[16] ,
    \sb_1__1__20_chanx_left_out[17] ,
    \sb_1__1__20_chanx_left_out[18] ,
    \sb_1__1__20_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__27_chanx_left_out[0] ,
    \cbx_1__1__27_chanx_left_out[1] ,
    \cbx_1__1__27_chanx_left_out[2] ,
    \cbx_1__1__27_chanx_left_out[3] ,
    \cbx_1__1__27_chanx_left_out[4] ,
    \cbx_1__1__27_chanx_left_out[5] ,
    \cbx_1__1__27_chanx_left_out[6] ,
    \cbx_1__1__27_chanx_left_out[7] ,
    \cbx_1__1__27_chanx_left_out[8] ,
    \cbx_1__1__27_chanx_left_out[9] ,
    \cbx_1__1__27_chanx_left_out[10] ,
    \cbx_1__1__27_chanx_left_out[11] ,
    \cbx_1__1__27_chanx_left_out[12] ,
    \cbx_1__1__27_chanx_left_out[13] ,
    \cbx_1__1__27_chanx_left_out[14] ,
    \cbx_1__1__27_chanx_left_out[15] ,
    \cbx_1__1__27_chanx_left_out[16] ,
    \cbx_1__1__27_chanx_left_out[17] ,
    \cbx_1__1__27_chanx_left_out[18] ,
    \cbx_1__1__27_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__20_chanx_right_out[0] ,
    \sb_1__1__20_chanx_right_out[1] ,
    \sb_1__1__20_chanx_right_out[2] ,
    \sb_1__1__20_chanx_right_out[3] ,
    \sb_1__1__20_chanx_right_out[4] ,
    \sb_1__1__20_chanx_right_out[5] ,
    \sb_1__1__20_chanx_right_out[6] ,
    \sb_1__1__20_chanx_right_out[7] ,
    \sb_1__1__20_chanx_right_out[8] ,
    \sb_1__1__20_chanx_right_out[9] ,
    \sb_1__1__20_chanx_right_out[10] ,
    \sb_1__1__20_chanx_right_out[11] ,
    \sb_1__1__20_chanx_right_out[12] ,
    \sb_1__1__20_chanx_right_out[13] ,
    \sb_1__1__20_chanx_right_out[14] ,
    \sb_1__1__20_chanx_right_out[15] ,
    \sb_1__1__20_chanx_right_out[16] ,
    \sb_1__1__20_chanx_right_out[17] ,
    \sb_1__1__20_chanx_right_out[18] ,
    \sb_1__1__20_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__22_chany_top_out[0] ,
    \cby_1__1__22_chany_top_out[1] ,
    \cby_1__1__22_chany_top_out[2] ,
    \cby_1__1__22_chany_top_out[3] ,
    \cby_1__1__22_chany_top_out[4] ,
    \cby_1__1__22_chany_top_out[5] ,
    \cby_1__1__22_chany_top_out[6] ,
    \cby_1__1__22_chany_top_out[7] ,
    \cby_1__1__22_chany_top_out[8] ,
    \cby_1__1__22_chany_top_out[9] ,
    \cby_1__1__22_chany_top_out[10] ,
    \cby_1__1__22_chany_top_out[11] ,
    \cby_1__1__22_chany_top_out[12] ,
    \cby_1__1__22_chany_top_out[13] ,
    \cby_1__1__22_chany_top_out[14] ,
    \cby_1__1__22_chany_top_out[15] ,
    \cby_1__1__22_chany_top_out[16] ,
    \cby_1__1__22_chany_top_out[17] ,
    \cby_1__1__22_chany_top_out[18] ,
    \cby_1__1__22_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__20_chany_bottom_out[0] ,
    \sb_1__1__20_chany_bottom_out[1] ,
    \sb_1__1__20_chany_bottom_out[2] ,
    \sb_1__1__20_chany_bottom_out[3] ,
    \sb_1__1__20_chany_bottom_out[4] ,
    \sb_1__1__20_chany_bottom_out[5] ,
    \sb_1__1__20_chany_bottom_out[6] ,
    \sb_1__1__20_chany_bottom_out[7] ,
    \sb_1__1__20_chany_bottom_out[8] ,
    \sb_1__1__20_chany_bottom_out[9] ,
    \sb_1__1__20_chany_bottom_out[10] ,
    \sb_1__1__20_chany_bottom_out[11] ,
    \sb_1__1__20_chany_bottom_out[12] ,
    \sb_1__1__20_chany_bottom_out[13] ,
    \sb_1__1__20_chany_bottom_out[14] ,
    \sb_1__1__20_chany_bottom_out[15] ,
    \sb_1__1__20_chany_bottom_out[16] ,
    \sb_1__1__20_chany_bottom_out[17] ,
    \sb_1__1__20_chany_bottom_out[18] ,
    \sb_1__1__20_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__23_chany_bottom_out[0] ,
    \cby_1__1__23_chany_bottom_out[1] ,
    \cby_1__1__23_chany_bottom_out[2] ,
    \cby_1__1__23_chany_bottom_out[3] ,
    \cby_1__1__23_chany_bottom_out[4] ,
    \cby_1__1__23_chany_bottom_out[5] ,
    \cby_1__1__23_chany_bottom_out[6] ,
    \cby_1__1__23_chany_bottom_out[7] ,
    \cby_1__1__23_chany_bottom_out[8] ,
    \cby_1__1__23_chany_bottom_out[9] ,
    \cby_1__1__23_chany_bottom_out[10] ,
    \cby_1__1__23_chany_bottom_out[11] ,
    \cby_1__1__23_chany_bottom_out[12] ,
    \cby_1__1__23_chany_bottom_out[13] ,
    \cby_1__1__23_chany_bottom_out[14] ,
    \cby_1__1__23_chany_bottom_out[15] ,
    \cby_1__1__23_chany_bottom_out[16] ,
    \cby_1__1__23_chany_bottom_out[17] ,
    \cby_1__1__23_chany_bottom_out[18] ,
    \cby_1__1__23_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__20_chany_top_out[0] ,
    \sb_1__1__20_chany_top_out[1] ,
    \sb_1__1__20_chany_top_out[2] ,
    \sb_1__1__20_chany_top_out[3] ,
    \sb_1__1__20_chany_top_out[4] ,
    \sb_1__1__20_chany_top_out[5] ,
    \sb_1__1__20_chany_top_out[6] ,
    \sb_1__1__20_chany_top_out[7] ,
    \sb_1__1__20_chany_top_out[8] ,
    \sb_1__1__20_chany_top_out[9] ,
    \sb_1__1__20_chany_top_out[10] ,
    \sb_1__1__20_chany_top_out[11] ,
    \sb_1__1__20_chany_top_out[12] ,
    \sb_1__1__20_chany_top_out[13] ,
    \sb_1__1__20_chany_top_out[14] ,
    \sb_1__1__20_chany_top_out[15] ,
    \sb_1__1__20_chany_top_out[16] ,
    \sb_1__1__20_chany_top_out[17] ,
    \sb_1__1__20_chany_top_out[18] ,
    \sb_1__1__20_chany_top_out[19] }));
 sb_1__2_ sb_3__8_ (.bottom_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_upper),
    .ccff_head(grid_io_top_3_ccff_tail),
    .ccff_tail(sb_1__8__2_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[94] ),
    .right_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__2_chanx_right_out[0] ,
    \cbx_1__8__2_chanx_right_out[1] ,
    \cbx_1__8__2_chanx_right_out[2] ,
    \cbx_1__8__2_chanx_right_out[3] ,
    \cbx_1__8__2_chanx_right_out[4] ,
    \cbx_1__8__2_chanx_right_out[5] ,
    \cbx_1__8__2_chanx_right_out[6] ,
    \cbx_1__8__2_chanx_right_out[7] ,
    \cbx_1__8__2_chanx_right_out[8] ,
    \cbx_1__8__2_chanx_right_out[9] ,
    \cbx_1__8__2_chanx_right_out[10] ,
    \cbx_1__8__2_chanx_right_out[11] ,
    \cbx_1__8__2_chanx_right_out[12] ,
    \cbx_1__8__2_chanx_right_out[13] ,
    \cbx_1__8__2_chanx_right_out[14] ,
    \cbx_1__8__2_chanx_right_out[15] ,
    \cbx_1__8__2_chanx_right_out[16] ,
    \cbx_1__8__2_chanx_right_out[17] ,
    \cbx_1__8__2_chanx_right_out[18] ,
    \cbx_1__8__2_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__8__2_chanx_left_out[0] ,
    \sb_1__8__2_chanx_left_out[1] ,
    \sb_1__8__2_chanx_left_out[2] ,
    \sb_1__8__2_chanx_left_out[3] ,
    \sb_1__8__2_chanx_left_out[4] ,
    \sb_1__8__2_chanx_left_out[5] ,
    \sb_1__8__2_chanx_left_out[6] ,
    \sb_1__8__2_chanx_left_out[7] ,
    \sb_1__8__2_chanx_left_out[8] ,
    \sb_1__8__2_chanx_left_out[9] ,
    \sb_1__8__2_chanx_left_out[10] ,
    \sb_1__8__2_chanx_left_out[11] ,
    \sb_1__8__2_chanx_left_out[12] ,
    \sb_1__8__2_chanx_left_out[13] ,
    \sb_1__8__2_chanx_left_out[14] ,
    \sb_1__8__2_chanx_left_out[15] ,
    \sb_1__8__2_chanx_left_out[16] ,
    \sb_1__8__2_chanx_left_out[17] ,
    \sb_1__8__2_chanx_left_out[18] ,
    \sb_1__8__2_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__8__3_chanx_left_out[0] ,
    \cbx_1__8__3_chanx_left_out[1] ,
    \cbx_1__8__3_chanx_left_out[2] ,
    \cbx_1__8__3_chanx_left_out[3] ,
    \cbx_1__8__3_chanx_left_out[4] ,
    \cbx_1__8__3_chanx_left_out[5] ,
    \cbx_1__8__3_chanx_left_out[6] ,
    \cbx_1__8__3_chanx_left_out[7] ,
    \cbx_1__8__3_chanx_left_out[8] ,
    \cbx_1__8__3_chanx_left_out[9] ,
    \cbx_1__8__3_chanx_left_out[10] ,
    \cbx_1__8__3_chanx_left_out[11] ,
    \cbx_1__8__3_chanx_left_out[12] ,
    \cbx_1__8__3_chanx_left_out[13] ,
    \cbx_1__8__3_chanx_left_out[14] ,
    \cbx_1__8__3_chanx_left_out[15] ,
    \cbx_1__8__3_chanx_left_out[16] ,
    \cbx_1__8__3_chanx_left_out[17] ,
    \cbx_1__8__3_chanx_left_out[18] ,
    \cbx_1__8__3_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__8__2_chanx_right_out[0] ,
    \sb_1__8__2_chanx_right_out[1] ,
    \sb_1__8__2_chanx_right_out[2] ,
    \sb_1__8__2_chanx_right_out[3] ,
    \sb_1__8__2_chanx_right_out[4] ,
    \sb_1__8__2_chanx_right_out[5] ,
    \sb_1__8__2_chanx_right_out[6] ,
    \sb_1__8__2_chanx_right_out[7] ,
    \sb_1__8__2_chanx_right_out[8] ,
    \sb_1__8__2_chanx_right_out[9] ,
    \sb_1__8__2_chanx_right_out[10] ,
    \sb_1__8__2_chanx_right_out[11] ,
    \sb_1__8__2_chanx_right_out[12] ,
    \sb_1__8__2_chanx_right_out[13] ,
    \sb_1__8__2_chanx_right_out[14] ,
    \sb_1__8__2_chanx_right_out[15] ,
    \sb_1__8__2_chanx_right_out[16] ,
    \sb_1__8__2_chanx_right_out[17] ,
    \sb_1__8__2_chanx_right_out[18] ,
    \sb_1__8__2_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__23_chany_top_out[0] ,
    \cby_1__1__23_chany_top_out[1] ,
    \cby_1__1__23_chany_top_out[2] ,
    \cby_1__1__23_chany_top_out[3] ,
    \cby_1__1__23_chany_top_out[4] ,
    \cby_1__1__23_chany_top_out[5] ,
    \cby_1__1__23_chany_top_out[6] ,
    \cby_1__1__23_chany_top_out[7] ,
    \cby_1__1__23_chany_top_out[8] ,
    \cby_1__1__23_chany_top_out[9] ,
    \cby_1__1__23_chany_top_out[10] ,
    \cby_1__1__23_chany_top_out[11] ,
    \cby_1__1__23_chany_top_out[12] ,
    \cby_1__1__23_chany_top_out[13] ,
    \cby_1__1__23_chany_top_out[14] ,
    \cby_1__1__23_chany_top_out[15] ,
    \cby_1__1__23_chany_top_out[16] ,
    \cby_1__1__23_chany_top_out[17] ,
    \cby_1__1__23_chany_top_out[18] ,
    \cby_1__1__23_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__8__2_chany_bottom_out[0] ,
    \sb_1__8__2_chany_bottom_out[1] ,
    \sb_1__8__2_chany_bottom_out[2] ,
    \sb_1__8__2_chany_bottom_out[3] ,
    \sb_1__8__2_chany_bottom_out[4] ,
    \sb_1__8__2_chany_bottom_out[5] ,
    \sb_1__8__2_chany_bottom_out[6] ,
    \sb_1__8__2_chany_bottom_out[7] ,
    \sb_1__8__2_chany_bottom_out[8] ,
    \sb_1__8__2_chany_bottom_out[9] ,
    \sb_1__8__2_chany_bottom_out[10] ,
    \sb_1__8__2_chany_bottom_out[11] ,
    \sb_1__8__2_chany_bottom_out[12] ,
    \sb_1__8__2_chany_bottom_out[13] ,
    \sb_1__8__2_chany_bottom_out[14] ,
    \sb_1__8__2_chany_bottom_out[15] ,
    \sb_1__8__2_chany_bottom_out[16] ,
    \sb_1__8__2_chany_bottom_out[17] ,
    \sb_1__8__2_chany_bottom_out[18] ,
    \sb_1__8__2_chany_bottom_out[19] }));
 sb_1__0_ sb_4__0_ (.Test_en_N_out(\Test_enWires[1] ),
    .Test_en_S_in(Test_en),
    .ccff_head(grid_io_bottom_3_ccff_tail),
    .ccff_tail(sb_1__0__3_ccff_tail),
    .clk_3_N_out(\clk_3_wires[28] ),
    .clk_3_S_in(clk),
    .left_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[97] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[28] ),
    .prog_clk_3_S_in(prog_clk),
    .right_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__3_chanx_right_out[0] ,
    \cbx_1__0__3_chanx_right_out[1] ,
    \cbx_1__0__3_chanx_right_out[2] ,
    \cbx_1__0__3_chanx_right_out[3] ,
    \cbx_1__0__3_chanx_right_out[4] ,
    \cbx_1__0__3_chanx_right_out[5] ,
    \cbx_1__0__3_chanx_right_out[6] ,
    \cbx_1__0__3_chanx_right_out[7] ,
    \cbx_1__0__3_chanx_right_out[8] ,
    \cbx_1__0__3_chanx_right_out[9] ,
    \cbx_1__0__3_chanx_right_out[10] ,
    \cbx_1__0__3_chanx_right_out[11] ,
    \cbx_1__0__3_chanx_right_out[12] ,
    \cbx_1__0__3_chanx_right_out[13] ,
    \cbx_1__0__3_chanx_right_out[14] ,
    \cbx_1__0__3_chanx_right_out[15] ,
    \cbx_1__0__3_chanx_right_out[16] ,
    \cbx_1__0__3_chanx_right_out[17] ,
    \cbx_1__0__3_chanx_right_out[18] ,
    \cbx_1__0__3_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__0__3_chanx_left_out[0] ,
    \sb_1__0__3_chanx_left_out[1] ,
    \sb_1__0__3_chanx_left_out[2] ,
    \sb_1__0__3_chanx_left_out[3] ,
    \sb_1__0__3_chanx_left_out[4] ,
    \sb_1__0__3_chanx_left_out[5] ,
    \sb_1__0__3_chanx_left_out[6] ,
    \sb_1__0__3_chanx_left_out[7] ,
    \sb_1__0__3_chanx_left_out[8] ,
    \sb_1__0__3_chanx_left_out[9] ,
    \sb_1__0__3_chanx_left_out[10] ,
    \sb_1__0__3_chanx_left_out[11] ,
    \sb_1__0__3_chanx_left_out[12] ,
    \sb_1__0__3_chanx_left_out[13] ,
    \sb_1__0__3_chanx_left_out[14] ,
    \sb_1__0__3_chanx_left_out[15] ,
    \sb_1__0__3_chanx_left_out[16] ,
    \sb_1__0__3_chanx_left_out[17] ,
    \sb_1__0__3_chanx_left_out[18] ,
    \sb_1__0__3_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__0__4_chanx_left_out[0] ,
    \cbx_1__0__4_chanx_left_out[1] ,
    \cbx_1__0__4_chanx_left_out[2] ,
    \cbx_1__0__4_chanx_left_out[3] ,
    \cbx_1__0__4_chanx_left_out[4] ,
    \cbx_1__0__4_chanx_left_out[5] ,
    \cbx_1__0__4_chanx_left_out[6] ,
    \cbx_1__0__4_chanx_left_out[7] ,
    \cbx_1__0__4_chanx_left_out[8] ,
    \cbx_1__0__4_chanx_left_out[9] ,
    \cbx_1__0__4_chanx_left_out[10] ,
    \cbx_1__0__4_chanx_left_out[11] ,
    \cbx_1__0__4_chanx_left_out[12] ,
    \cbx_1__0__4_chanx_left_out[13] ,
    \cbx_1__0__4_chanx_left_out[14] ,
    \cbx_1__0__4_chanx_left_out[15] ,
    \cbx_1__0__4_chanx_left_out[16] ,
    \cbx_1__0__4_chanx_left_out[17] ,
    \cbx_1__0__4_chanx_left_out[18] ,
    \cbx_1__0__4_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__0__3_chanx_right_out[0] ,
    \sb_1__0__3_chanx_right_out[1] ,
    \sb_1__0__3_chanx_right_out[2] ,
    \sb_1__0__3_chanx_right_out[3] ,
    \sb_1__0__3_chanx_right_out[4] ,
    \sb_1__0__3_chanx_right_out[5] ,
    \sb_1__0__3_chanx_right_out[6] ,
    \sb_1__0__3_chanx_right_out[7] ,
    \sb_1__0__3_chanx_right_out[8] ,
    \sb_1__0__3_chanx_right_out[9] ,
    \sb_1__0__3_chanx_right_out[10] ,
    \sb_1__0__3_chanx_right_out[11] ,
    \sb_1__0__3_chanx_right_out[12] ,
    \sb_1__0__3_chanx_right_out[13] ,
    \sb_1__0__3_chanx_right_out[14] ,
    \sb_1__0__3_chanx_right_out[15] ,
    \sb_1__0__3_chanx_right_out[16] ,
    \sb_1__0__3_chanx_right_out[17] ,
    \sb_1__0__3_chanx_right_out[18] ,
    \sb_1__0__3_chanx_right_out[19] }),
    .chany_top_in({\cby_1__1__24_chany_bottom_out[0] ,
    \cby_1__1__24_chany_bottom_out[1] ,
    \cby_1__1__24_chany_bottom_out[2] ,
    \cby_1__1__24_chany_bottom_out[3] ,
    \cby_1__1__24_chany_bottom_out[4] ,
    \cby_1__1__24_chany_bottom_out[5] ,
    \cby_1__1__24_chany_bottom_out[6] ,
    \cby_1__1__24_chany_bottom_out[7] ,
    \cby_1__1__24_chany_bottom_out[8] ,
    \cby_1__1__24_chany_bottom_out[9] ,
    \cby_1__1__24_chany_bottom_out[10] ,
    \cby_1__1__24_chany_bottom_out[11] ,
    \cby_1__1__24_chany_bottom_out[12] ,
    \cby_1__1__24_chany_bottom_out[13] ,
    \cby_1__1__24_chany_bottom_out[14] ,
    \cby_1__1__24_chany_bottom_out[15] ,
    \cby_1__1__24_chany_bottom_out[16] ,
    \cby_1__1__24_chany_bottom_out[17] ,
    \cby_1__1__24_chany_bottom_out[18] ,
    \cby_1__1__24_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__0__3_chany_top_out[0] ,
    \sb_1__0__3_chany_top_out[1] ,
    \sb_1__0__3_chany_top_out[2] ,
    \sb_1__0__3_chany_top_out[3] ,
    \sb_1__0__3_chany_top_out[4] ,
    \sb_1__0__3_chany_top_out[5] ,
    \sb_1__0__3_chany_top_out[6] ,
    \sb_1__0__3_chany_top_out[7] ,
    \sb_1__0__3_chany_top_out[8] ,
    \sb_1__0__3_chany_top_out[9] ,
    \sb_1__0__3_chany_top_out[10] ,
    \sb_1__0__3_chany_top_out[11] ,
    \sb_1__0__3_chany_top_out[12] ,
    \sb_1__0__3_chany_top_out[13] ,
    \sb_1__0__3_chany_top_out[14] ,
    \sb_1__0__3_chany_top_out[15] ,
    \sb_1__0__3_chany_top_out[16] ,
    \sb_1__0__3_chany_top_out[17] ,
    \sb_1__0__3_chany_top_out[18] ,
    \sb_1__0__3_chany_top_out[19] }));
 sb_1__1_ sb_4__1_ (.Test_en_N_out(\Test_enWires[3] ),
    .Test_en_S_in(\Test_enWires[2] ),
    .bottom_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__28_ccff_tail),
    .ccff_tail(sb_1__1__21_ccff_tail),
    .clk_3_N_in(\clk_3_wires[27] ),
    .clk_3_N_out(\clk_3_wires[30] ),
    .left_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[100] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[27] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[30] ),
    .right_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__21_chanx_right_out[0] ,
    \cbx_1__1__21_chanx_right_out[1] ,
    \cbx_1__1__21_chanx_right_out[2] ,
    \cbx_1__1__21_chanx_right_out[3] ,
    \cbx_1__1__21_chanx_right_out[4] ,
    \cbx_1__1__21_chanx_right_out[5] ,
    \cbx_1__1__21_chanx_right_out[6] ,
    \cbx_1__1__21_chanx_right_out[7] ,
    \cbx_1__1__21_chanx_right_out[8] ,
    \cbx_1__1__21_chanx_right_out[9] ,
    \cbx_1__1__21_chanx_right_out[10] ,
    \cbx_1__1__21_chanx_right_out[11] ,
    \cbx_1__1__21_chanx_right_out[12] ,
    \cbx_1__1__21_chanx_right_out[13] ,
    \cbx_1__1__21_chanx_right_out[14] ,
    \cbx_1__1__21_chanx_right_out[15] ,
    \cbx_1__1__21_chanx_right_out[16] ,
    \cbx_1__1__21_chanx_right_out[17] ,
    \cbx_1__1__21_chanx_right_out[18] ,
    \cbx_1__1__21_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__21_chanx_left_out[0] ,
    \sb_1__1__21_chanx_left_out[1] ,
    \sb_1__1__21_chanx_left_out[2] ,
    \sb_1__1__21_chanx_left_out[3] ,
    \sb_1__1__21_chanx_left_out[4] ,
    \sb_1__1__21_chanx_left_out[5] ,
    \sb_1__1__21_chanx_left_out[6] ,
    \sb_1__1__21_chanx_left_out[7] ,
    \sb_1__1__21_chanx_left_out[8] ,
    \sb_1__1__21_chanx_left_out[9] ,
    \sb_1__1__21_chanx_left_out[10] ,
    \sb_1__1__21_chanx_left_out[11] ,
    \sb_1__1__21_chanx_left_out[12] ,
    \sb_1__1__21_chanx_left_out[13] ,
    \sb_1__1__21_chanx_left_out[14] ,
    \sb_1__1__21_chanx_left_out[15] ,
    \sb_1__1__21_chanx_left_out[16] ,
    \sb_1__1__21_chanx_left_out[17] ,
    \sb_1__1__21_chanx_left_out[18] ,
    \sb_1__1__21_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__28_chanx_left_out[0] ,
    \cbx_1__1__28_chanx_left_out[1] ,
    \cbx_1__1__28_chanx_left_out[2] ,
    \cbx_1__1__28_chanx_left_out[3] ,
    \cbx_1__1__28_chanx_left_out[4] ,
    \cbx_1__1__28_chanx_left_out[5] ,
    \cbx_1__1__28_chanx_left_out[6] ,
    \cbx_1__1__28_chanx_left_out[7] ,
    \cbx_1__1__28_chanx_left_out[8] ,
    \cbx_1__1__28_chanx_left_out[9] ,
    \cbx_1__1__28_chanx_left_out[10] ,
    \cbx_1__1__28_chanx_left_out[11] ,
    \cbx_1__1__28_chanx_left_out[12] ,
    \cbx_1__1__28_chanx_left_out[13] ,
    \cbx_1__1__28_chanx_left_out[14] ,
    \cbx_1__1__28_chanx_left_out[15] ,
    \cbx_1__1__28_chanx_left_out[16] ,
    \cbx_1__1__28_chanx_left_out[17] ,
    \cbx_1__1__28_chanx_left_out[18] ,
    \cbx_1__1__28_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__21_chanx_right_out[0] ,
    \sb_1__1__21_chanx_right_out[1] ,
    \sb_1__1__21_chanx_right_out[2] ,
    \sb_1__1__21_chanx_right_out[3] ,
    \sb_1__1__21_chanx_right_out[4] ,
    \sb_1__1__21_chanx_right_out[5] ,
    \sb_1__1__21_chanx_right_out[6] ,
    \sb_1__1__21_chanx_right_out[7] ,
    \sb_1__1__21_chanx_right_out[8] ,
    \sb_1__1__21_chanx_right_out[9] ,
    \sb_1__1__21_chanx_right_out[10] ,
    \sb_1__1__21_chanx_right_out[11] ,
    \sb_1__1__21_chanx_right_out[12] ,
    \sb_1__1__21_chanx_right_out[13] ,
    \sb_1__1__21_chanx_right_out[14] ,
    \sb_1__1__21_chanx_right_out[15] ,
    \sb_1__1__21_chanx_right_out[16] ,
    \sb_1__1__21_chanx_right_out[17] ,
    \sb_1__1__21_chanx_right_out[18] ,
    \sb_1__1__21_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__24_chany_top_out[0] ,
    \cby_1__1__24_chany_top_out[1] ,
    \cby_1__1__24_chany_top_out[2] ,
    \cby_1__1__24_chany_top_out[3] ,
    \cby_1__1__24_chany_top_out[4] ,
    \cby_1__1__24_chany_top_out[5] ,
    \cby_1__1__24_chany_top_out[6] ,
    \cby_1__1__24_chany_top_out[7] ,
    \cby_1__1__24_chany_top_out[8] ,
    \cby_1__1__24_chany_top_out[9] ,
    \cby_1__1__24_chany_top_out[10] ,
    \cby_1__1__24_chany_top_out[11] ,
    \cby_1__1__24_chany_top_out[12] ,
    \cby_1__1__24_chany_top_out[13] ,
    \cby_1__1__24_chany_top_out[14] ,
    \cby_1__1__24_chany_top_out[15] ,
    \cby_1__1__24_chany_top_out[16] ,
    \cby_1__1__24_chany_top_out[17] ,
    \cby_1__1__24_chany_top_out[18] ,
    \cby_1__1__24_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__21_chany_bottom_out[0] ,
    \sb_1__1__21_chany_bottom_out[1] ,
    \sb_1__1__21_chany_bottom_out[2] ,
    \sb_1__1__21_chany_bottom_out[3] ,
    \sb_1__1__21_chany_bottom_out[4] ,
    \sb_1__1__21_chany_bottom_out[5] ,
    \sb_1__1__21_chany_bottom_out[6] ,
    \sb_1__1__21_chany_bottom_out[7] ,
    \sb_1__1__21_chany_bottom_out[8] ,
    \sb_1__1__21_chany_bottom_out[9] ,
    \sb_1__1__21_chany_bottom_out[10] ,
    \sb_1__1__21_chany_bottom_out[11] ,
    \sb_1__1__21_chany_bottom_out[12] ,
    \sb_1__1__21_chany_bottom_out[13] ,
    \sb_1__1__21_chany_bottom_out[14] ,
    \sb_1__1__21_chany_bottom_out[15] ,
    \sb_1__1__21_chany_bottom_out[16] ,
    \sb_1__1__21_chany_bottom_out[17] ,
    \sb_1__1__21_chany_bottom_out[18] ,
    \sb_1__1__21_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__25_chany_bottom_out[0] ,
    \cby_1__1__25_chany_bottom_out[1] ,
    \cby_1__1__25_chany_bottom_out[2] ,
    \cby_1__1__25_chany_bottom_out[3] ,
    \cby_1__1__25_chany_bottom_out[4] ,
    \cby_1__1__25_chany_bottom_out[5] ,
    \cby_1__1__25_chany_bottom_out[6] ,
    \cby_1__1__25_chany_bottom_out[7] ,
    \cby_1__1__25_chany_bottom_out[8] ,
    \cby_1__1__25_chany_bottom_out[9] ,
    \cby_1__1__25_chany_bottom_out[10] ,
    \cby_1__1__25_chany_bottom_out[11] ,
    \cby_1__1__25_chany_bottom_out[12] ,
    \cby_1__1__25_chany_bottom_out[13] ,
    \cby_1__1__25_chany_bottom_out[14] ,
    \cby_1__1__25_chany_bottom_out[15] ,
    \cby_1__1__25_chany_bottom_out[16] ,
    \cby_1__1__25_chany_bottom_out[17] ,
    \cby_1__1__25_chany_bottom_out[18] ,
    \cby_1__1__25_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__21_chany_top_out[0] ,
    \sb_1__1__21_chany_top_out[1] ,
    \sb_1__1__21_chany_top_out[2] ,
    \sb_1__1__21_chany_top_out[3] ,
    \sb_1__1__21_chany_top_out[4] ,
    \sb_1__1__21_chany_top_out[5] ,
    \sb_1__1__21_chany_top_out[6] ,
    \sb_1__1__21_chany_top_out[7] ,
    \sb_1__1__21_chany_top_out[8] ,
    \sb_1__1__21_chany_top_out[9] ,
    \sb_1__1__21_chany_top_out[10] ,
    \sb_1__1__21_chany_top_out[11] ,
    \sb_1__1__21_chany_top_out[12] ,
    \sb_1__1__21_chany_top_out[13] ,
    \sb_1__1__21_chany_top_out[14] ,
    \sb_1__1__21_chany_top_out[15] ,
    \sb_1__1__21_chany_top_out[16] ,
    \sb_1__1__21_chany_top_out[17] ,
    \sb_1__1__21_chany_top_out[18] ,
    \sb_1__1__21_chany_top_out[19] }));
 sb_1__1_ sb_4__2_ (.Test_en_N_out(\Test_enWires[5] ),
    .Test_en_S_in(\Test_enWires[4] ),
    .bottom_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__29_ccff_tail),
    .ccff_tail(sb_1__1__22_ccff_tail),
    .clk_3_N_in(\clk_3_wires[29] ),
    .clk_3_N_out(\clk_3_wires[32] ),
    .left_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[103] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[29] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[32] ),
    .right_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__22_chanx_right_out[0] ,
    \cbx_1__1__22_chanx_right_out[1] ,
    \cbx_1__1__22_chanx_right_out[2] ,
    \cbx_1__1__22_chanx_right_out[3] ,
    \cbx_1__1__22_chanx_right_out[4] ,
    \cbx_1__1__22_chanx_right_out[5] ,
    \cbx_1__1__22_chanx_right_out[6] ,
    \cbx_1__1__22_chanx_right_out[7] ,
    \cbx_1__1__22_chanx_right_out[8] ,
    \cbx_1__1__22_chanx_right_out[9] ,
    \cbx_1__1__22_chanx_right_out[10] ,
    \cbx_1__1__22_chanx_right_out[11] ,
    \cbx_1__1__22_chanx_right_out[12] ,
    \cbx_1__1__22_chanx_right_out[13] ,
    \cbx_1__1__22_chanx_right_out[14] ,
    \cbx_1__1__22_chanx_right_out[15] ,
    \cbx_1__1__22_chanx_right_out[16] ,
    \cbx_1__1__22_chanx_right_out[17] ,
    \cbx_1__1__22_chanx_right_out[18] ,
    \cbx_1__1__22_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__22_chanx_left_out[0] ,
    \sb_1__1__22_chanx_left_out[1] ,
    \sb_1__1__22_chanx_left_out[2] ,
    \sb_1__1__22_chanx_left_out[3] ,
    \sb_1__1__22_chanx_left_out[4] ,
    \sb_1__1__22_chanx_left_out[5] ,
    \sb_1__1__22_chanx_left_out[6] ,
    \sb_1__1__22_chanx_left_out[7] ,
    \sb_1__1__22_chanx_left_out[8] ,
    \sb_1__1__22_chanx_left_out[9] ,
    \sb_1__1__22_chanx_left_out[10] ,
    \sb_1__1__22_chanx_left_out[11] ,
    \sb_1__1__22_chanx_left_out[12] ,
    \sb_1__1__22_chanx_left_out[13] ,
    \sb_1__1__22_chanx_left_out[14] ,
    \sb_1__1__22_chanx_left_out[15] ,
    \sb_1__1__22_chanx_left_out[16] ,
    \sb_1__1__22_chanx_left_out[17] ,
    \sb_1__1__22_chanx_left_out[18] ,
    \sb_1__1__22_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__29_chanx_left_out[0] ,
    \cbx_1__1__29_chanx_left_out[1] ,
    \cbx_1__1__29_chanx_left_out[2] ,
    \cbx_1__1__29_chanx_left_out[3] ,
    \cbx_1__1__29_chanx_left_out[4] ,
    \cbx_1__1__29_chanx_left_out[5] ,
    \cbx_1__1__29_chanx_left_out[6] ,
    \cbx_1__1__29_chanx_left_out[7] ,
    \cbx_1__1__29_chanx_left_out[8] ,
    \cbx_1__1__29_chanx_left_out[9] ,
    \cbx_1__1__29_chanx_left_out[10] ,
    \cbx_1__1__29_chanx_left_out[11] ,
    \cbx_1__1__29_chanx_left_out[12] ,
    \cbx_1__1__29_chanx_left_out[13] ,
    \cbx_1__1__29_chanx_left_out[14] ,
    \cbx_1__1__29_chanx_left_out[15] ,
    \cbx_1__1__29_chanx_left_out[16] ,
    \cbx_1__1__29_chanx_left_out[17] ,
    \cbx_1__1__29_chanx_left_out[18] ,
    \cbx_1__1__29_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__22_chanx_right_out[0] ,
    \sb_1__1__22_chanx_right_out[1] ,
    \sb_1__1__22_chanx_right_out[2] ,
    \sb_1__1__22_chanx_right_out[3] ,
    \sb_1__1__22_chanx_right_out[4] ,
    \sb_1__1__22_chanx_right_out[5] ,
    \sb_1__1__22_chanx_right_out[6] ,
    \sb_1__1__22_chanx_right_out[7] ,
    \sb_1__1__22_chanx_right_out[8] ,
    \sb_1__1__22_chanx_right_out[9] ,
    \sb_1__1__22_chanx_right_out[10] ,
    \sb_1__1__22_chanx_right_out[11] ,
    \sb_1__1__22_chanx_right_out[12] ,
    \sb_1__1__22_chanx_right_out[13] ,
    \sb_1__1__22_chanx_right_out[14] ,
    \sb_1__1__22_chanx_right_out[15] ,
    \sb_1__1__22_chanx_right_out[16] ,
    \sb_1__1__22_chanx_right_out[17] ,
    \sb_1__1__22_chanx_right_out[18] ,
    \sb_1__1__22_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__25_chany_top_out[0] ,
    \cby_1__1__25_chany_top_out[1] ,
    \cby_1__1__25_chany_top_out[2] ,
    \cby_1__1__25_chany_top_out[3] ,
    \cby_1__1__25_chany_top_out[4] ,
    \cby_1__1__25_chany_top_out[5] ,
    \cby_1__1__25_chany_top_out[6] ,
    \cby_1__1__25_chany_top_out[7] ,
    \cby_1__1__25_chany_top_out[8] ,
    \cby_1__1__25_chany_top_out[9] ,
    \cby_1__1__25_chany_top_out[10] ,
    \cby_1__1__25_chany_top_out[11] ,
    \cby_1__1__25_chany_top_out[12] ,
    \cby_1__1__25_chany_top_out[13] ,
    \cby_1__1__25_chany_top_out[14] ,
    \cby_1__1__25_chany_top_out[15] ,
    \cby_1__1__25_chany_top_out[16] ,
    \cby_1__1__25_chany_top_out[17] ,
    \cby_1__1__25_chany_top_out[18] ,
    \cby_1__1__25_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__22_chany_bottom_out[0] ,
    \sb_1__1__22_chany_bottom_out[1] ,
    \sb_1__1__22_chany_bottom_out[2] ,
    \sb_1__1__22_chany_bottom_out[3] ,
    \sb_1__1__22_chany_bottom_out[4] ,
    \sb_1__1__22_chany_bottom_out[5] ,
    \sb_1__1__22_chany_bottom_out[6] ,
    \sb_1__1__22_chany_bottom_out[7] ,
    \sb_1__1__22_chany_bottom_out[8] ,
    \sb_1__1__22_chany_bottom_out[9] ,
    \sb_1__1__22_chany_bottom_out[10] ,
    \sb_1__1__22_chany_bottom_out[11] ,
    \sb_1__1__22_chany_bottom_out[12] ,
    \sb_1__1__22_chany_bottom_out[13] ,
    \sb_1__1__22_chany_bottom_out[14] ,
    \sb_1__1__22_chany_bottom_out[15] ,
    \sb_1__1__22_chany_bottom_out[16] ,
    \sb_1__1__22_chany_bottom_out[17] ,
    \sb_1__1__22_chany_bottom_out[18] ,
    \sb_1__1__22_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__26_chany_bottom_out[0] ,
    \cby_1__1__26_chany_bottom_out[1] ,
    \cby_1__1__26_chany_bottom_out[2] ,
    \cby_1__1__26_chany_bottom_out[3] ,
    \cby_1__1__26_chany_bottom_out[4] ,
    \cby_1__1__26_chany_bottom_out[5] ,
    \cby_1__1__26_chany_bottom_out[6] ,
    \cby_1__1__26_chany_bottom_out[7] ,
    \cby_1__1__26_chany_bottom_out[8] ,
    \cby_1__1__26_chany_bottom_out[9] ,
    \cby_1__1__26_chany_bottom_out[10] ,
    \cby_1__1__26_chany_bottom_out[11] ,
    \cby_1__1__26_chany_bottom_out[12] ,
    \cby_1__1__26_chany_bottom_out[13] ,
    \cby_1__1__26_chany_bottom_out[14] ,
    \cby_1__1__26_chany_bottom_out[15] ,
    \cby_1__1__26_chany_bottom_out[16] ,
    \cby_1__1__26_chany_bottom_out[17] ,
    \cby_1__1__26_chany_bottom_out[18] ,
    \cby_1__1__26_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__22_chany_top_out[0] ,
    \sb_1__1__22_chany_top_out[1] ,
    \sb_1__1__22_chany_top_out[2] ,
    \sb_1__1__22_chany_top_out[3] ,
    \sb_1__1__22_chany_top_out[4] ,
    \sb_1__1__22_chany_top_out[5] ,
    \sb_1__1__22_chany_top_out[6] ,
    \sb_1__1__22_chany_top_out[7] ,
    \sb_1__1__22_chany_top_out[8] ,
    \sb_1__1__22_chany_top_out[9] ,
    \sb_1__1__22_chany_top_out[10] ,
    \sb_1__1__22_chany_top_out[11] ,
    \sb_1__1__22_chany_top_out[12] ,
    \sb_1__1__22_chany_top_out[13] ,
    \sb_1__1__22_chany_top_out[14] ,
    \sb_1__1__22_chany_top_out[15] ,
    \sb_1__1__22_chany_top_out[16] ,
    \sb_1__1__22_chany_top_out[17] ,
    \sb_1__1__22_chany_top_out[18] ,
    \sb_1__1__22_chany_top_out[19] }));
 sb_1__1_ sb_4__3_ (.Test_en_N_out(\Test_enWires[7] ),
    .Test_en_S_in(\Test_enWires[6] ),
    .bottom_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__30_ccff_tail),
    .ccff_tail(sb_1__1__23_ccff_tail),
    .clk_3_N_in(\clk_3_wires[31] ),
    .clk_3_N_out(\clk_3_wires[34] ),
    .left_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[106] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[31] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[34] ),
    .right_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__23_chanx_right_out[0] ,
    \cbx_1__1__23_chanx_right_out[1] ,
    \cbx_1__1__23_chanx_right_out[2] ,
    \cbx_1__1__23_chanx_right_out[3] ,
    \cbx_1__1__23_chanx_right_out[4] ,
    \cbx_1__1__23_chanx_right_out[5] ,
    \cbx_1__1__23_chanx_right_out[6] ,
    \cbx_1__1__23_chanx_right_out[7] ,
    \cbx_1__1__23_chanx_right_out[8] ,
    \cbx_1__1__23_chanx_right_out[9] ,
    \cbx_1__1__23_chanx_right_out[10] ,
    \cbx_1__1__23_chanx_right_out[11] ,
    \cbx_1__1__23_chanx_right_out[12] ,
    \cbx_1__1__23_chanx_right_out[13] ,
    \cbx_1__1__23_chanx_right_out[14] ,
    \cbx_1__1__23_chanx_right_out[15] ,
    \cbx_1__1__23_chanx_right_out[16] ,
    \cbx_1__1__23_chanx_right_out[17] ,
    \cbx_1__1__23_chanx_right_out[18] ,
    \cbx_1__1__23_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__23_chanx_left_out[0] ,
    \sb_1__1__23_chanx_left_out[1] ,
    \sb_1__1__23_chanx_left_out[2] ,
    \sb_1__1__23_chanx_left_out[3] ,
    \sb_1__1__23_chanx_left_out[4] ,
    \sb_1__1__23_chanx_left_out[5] ,
    \sb_1__1__23_chanx_left_out[6] ,
    \sb_1__1__23_chanx_left_out[7] ,
    \sb_1__1__23_chanx_left_out[8] ,
    \sb_1__1__23_chanx_left_out[9] ,
    \sb_1__1__23_chanx_left_out[10] ,
    \sb_1__1__23_chanx_left_out[11] ,
    \sb_1__1__23_chanx_left_out[12] ,
    \sb_1__1__23_chanx_left_out[13] ,
    \sb_1__1__23_chanx_left_out[14] ,
    \sb_1__1__23_chanx_left_out[15] ,
    \sb_1__1__23_chanx_left_out[16] ,
    \sb_1__1__23_chanx_left_out[17] ,
    \sb_1__1__23_chanx_left_out[18] ,
    \sb_1__1__23_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__30_chanx_left_out[0] ,
    \cbx_1__1__30_chanx_left_out[1] ,
    \cbx_1__1__30_chanx_left_out[2] ,
    \cbx_1__1__30_chanx_left_out[3] ,
    \cbx_1__1__30_chanx_left_out[4] ,
    \cbx_1__1__30_chanx_left_out[5] ,
    \cbx_1__1__30_chanx_left_out[6] ,
    \cbx_1__1__30_chanx_left_out[7] ,
    \cbx_1__1__30_chanx_left_out[8] ,
    \cbx_1__1__30_chanx_left_out[9] ,
    \cbx_1__1__30_chanx_left_out[10] ,
    \cbx_1__1__30_chanx_left_out[11] ,
    \cbx_1__1__30_chanx_left_out[12] ,
    \cbx_1__1__30_chanx_left_out[13] ,
    \cbx_1__1__30_chanx_left_out[14] ,
    \cbx_1__1__30_chanx_left_out[15] ,
    \cbx_1__1__30_chanx_left_out[16] ,
    \cbx_1__1__30_chanx_left_out[17] ,
    \cbx_1__1__30_chanx_left_out[18] ,
    \cbx_1__1__30_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__23_chanx_right_out[0] ,
    \sb_1__1__23_chanx_right_out[1] ,
    \sb_1__1__23_chanx_right_out[2] ,
    \sb_1__1__23_chanx_right_out[3] ,
    \sb_1__1__23_chanx_right_out[4] ,
    \sb_1__1__23_chanx_right_out[5] ,
    \sb_1__1__23_chanx_right_out[6] ,
    \sb_1__1__23_chanx_right_out[7] ,
    \sb_1__1__23_chanx_right_out[8] ,
    \sb_1__1__23_chanx_right_out[9] ,
    \sb_1__1__23_chanx_right_out[10] ,
    \sb_1__1__23_chanx_right_out[11] ,
    \sb_1__1__23_chanx_right_out[12] ,
    \sb_1__1__23_chanx_right_out[13] ,
    \sb_1__1__23_chanx_right_out[14] ,
    \sb_1__1__23_chanx_right_out[15] ,
    \sb_1__1__23_chanx_right_out[16] ,
    \sb_1__1__23_chanx_right_out[17] ,
    \sb_1__1__23_chanx_right_out[18] ,
    \sb_1__1__23_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__26_chany_top_out[0] ,
    \cby_1__1__26_chany_top_out[1] ,
    \cby_1__1__26_chany_top_out[2] ,
    \cby_1__1__26_chany_top_out[3] ,
    \cby_1__1__26_chany_top_out[4] ,
    \cby_1__1__26_chany_top_out[5] ,
    \cby_1__1__26_chany_top_out[6] ,
    \cby_1__1__26_chany_top_out[7] ,
    \cby_1__1__26_chany_top_out[8] ,
    \cby_1__1__26_chany_top_out[9] ,
    \cby_1__1__26_chany_top_out[10] ,
    \cby_1__1__26_chany_top_out[11] ,
    \cby_1__1__26_chany_top_out[12] ,
    \cby_1__1__26_chany_top_out[13] ,
    \cby_1__1__26_chany_top_out[14] ,
    \cby_1__1__26_chany_top_out[15] ,
    \cby_1__1__26_chany_top_out[16] ,
    \cby_1__1__26_chany_top_out[17] ,
    \cby_1__1__26_chany_top_out[18] ,
    \cby_1__1__26_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__23_chany_bottom_out[0] ,
    \sb_1__1__23_chany_bottom_out[1] ,
    \sb_1__1__23_chany_bottom_out[2] ,
    \sb_1__1__23_chany_bottom_out[3] ,
    \sb_1__1__23_chany_bottom_out[4] ,
    \sb_1__1__23_chany_bottom_out[5] ,
    \sb_1__1__23_chany_bottom_out[6] ,
    \sb_1__1__23_chany_bottom_out[7] ,
    \sb_1__1__23_chany_bottom_out[8] ,
    \sb_1__1__23_chany_bottom_out[9] ,
    \sb_1__1__23_chany_bottom_out[10] ,
    \sb_1__1__23_chany_bottom_out[11] ,
    \sb_1__1__23_chany_bottom_out[12] ,
    \sb_1__1__23_chany_bottom_out[13] ,
    \sb_1__1__23_chany_bottom_out[14] ,
    \sb_1__1__23_chany_bottom_out[15] ,
    \sb_1__1__23_chany_bottom_out[16] ,
    \sb_1__1__23_chany_bottom_out[17] ,
    \sb_1__1__23_chany_bottom_out[18] ,
    \sb_1__1__23_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__27_chany_bottom_out[0] ,
    \cby_1__1__27_chany_bottom_out[1] ,
    \cby_1__1__27_chany_bottom_out[2] ,
    \cby_1__1__27_chany_bottom_out[3] ,
    \cby_1__1__27_chany_bottom_out[4] ,
    \cby_1__1__27_chany_bottom_out[5] ,
    \cby_1__1__27_chany_bottom_out[6] ,
    \cby_1__1__27_chany_bottom_out[7] ,
    \cby_1__1__27_chany_bottom_out[8] ,
    \cby_1__1__27_chany_bottom_out[9] ,
    \cby_1__1__27_chany_bottom_out[10] ,
    \cby_1__1__27_chany_bottom_out[11] ,
    \cby_1__1__27_chany_bottom_out[12] ,
    \cby_1__1__27_chany_bottom_out[13] ,
    \cby_1__1__27_chany_bottom_out[14] ,
    \cby_1__1__27_chany_bottom_out[15] ,
    \cby_1__1__27_chany_bottom_out[16] ,
    \cby_1__1__27_chany_bottom_out[17] ,
    \cby_1__1__27_chany_bottom_out[18] ,
    \cby_1__1__27_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__23_chany_top_out[0] ,
    \sb_1__1__23_chany_top_out[1] ,
    \sb_1__1__23_chany_top_out[2] ,
    \sb_1__1__23_chany_top_out[3] ,
    \sb_1__1__23_chany_top_out[4] ,
    \sb_1__1__23_chany_top_out[5] ,
    \sb_1__1__23_chany_top_out[6] ,
    \sb_1__1__23_chany_top_out[7] ,
    \sb_1__1__23_chany_top_out[8] ,
    \sb_1__1__23_chany_top_out[9] ,
    \sb_1__1__23_chany_top_out[10] ,
    \sb_1__1__23_chany_top_out[11] ,
    \sb_1__1__23_chany_top_out[12] ,
    \sb_1__1__23_chany_top_out[13] ,
    \sb_1__1__23_chany_top_out[14] ,
    \sb_1__1__23_chany_top_out[15] ,
    \sb_1__1__23_chany_top_out[16] ,
    \sb_1__1__23_chany_top_out[17] ,
    \sb_1__1__23_chany_top_out[18] ,
    \sb_1__1__23_chany_top_out[19] }));
 sb_1__1_ sb_4__4_ (.Test_en_N_out(\Test_enWires[9] ),
    .Test_en_S_in(\Test_enWires[8] ),
    .bottom_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__31_ccff_tail),
    .ccff_tail(sb_1__1__24_ccff_tail),
    .clk_3_E_out(\clk_3_wires[1] ),
    .clk_3_N_in(\clk_3_wires[33] ),
    .clk_3_W_out(\clk_3_wires[3] ),
    .left_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[109] ),
    .prog_clk_3_E_out(\prog_clk_3_wires[1] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[33] ),
    .prog_clk_3_W_out(\prog_clk_3_wires[3] ),
    .right_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__24_chanx_right_out[0] ,
    \cbx_1__1__24_chanx_right_out[1] ,
    \cbx_1__1__24_chanx_right_out[2] ,
    \cbx_1__1__24_chanx_right_out[3] ,
    \cbx_1__1__24_chanx_right_out[4] ,
    \cbx_1__1__24_chanx_right_out[5] ,
    \cbx_1__1__24_chanx_right_out[6] ,
    \cbx_1__1__24_chanx_right_out[7] ,
    \cbx_1__1__24_chanx_right_out[8] ,
    \cbx_1__1__24_chanx_right_out[9] ,
    \cbx_1__1__24_chanx_right_out[10] ,
    \cbx_1__1__24_chanx_right_out[11] ,
    \cbx_1__1__24_chanx_right_out[12] ,
    \cbx_1__1__24_chanx_right_out[13] ,
    \cbx_1__1__24_chanx_right_out[14] ,
    \cbx_1__1__24_chanx_right_out[15] ,
    \cbx_1__1__24_chanx_right_out[16] ,
    \cbx_1__1__24_chanx_right_out[17] ,
    \cbx_1__1__24_chanx_right_out[18] ,
    \cbx_1__1__24_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__24_chanx_left_out[0] ,
    \sb_1__1__24_chanx_left_out[1] ,
    \sb_1__1__24_chanx_left_out[2] ,
    \sb_1__1__24_chanx_left_out[3] ,
    \sb_1__1__24_chanx_left_out[4] ,
    \sb_1__1__24_chanx_left_out[5] ,
    \sb_1__1__24_chanx_left_out[6] ,
    \sb_1__1__24_chanx_left_out[7] ,
    \sb_1__1__24_chanx_left_out[8] ,
    \sb_1__1__24_chanx_left_out[9] ,
    \sb_1__1__24_chanx_left_out[10] ,
    \sb_1__1__24_chanx_left_out[11] ,
    \sb_1__1__24_chanx_left_out[12] ,
    \sb_1__1__24_chanx_left_out[13] ,
    \sb_1__1__24_chanx_left_out[14] ,
    \sb_1__1__24_chanx_left_out[15] ,
    \sb_1__1__24_chanx_left_out[16] ,
    \sb_1__1__24_chanx_left_out[17] ,
    \sb_1__1__24_chanx_left_out[18] ,
    \sb_1__1__24_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__31_chanx_left_out[0] ,
    \cbx_1__1__31_chanx_left_out[1] ,
    \cbx_1__1__31_chanx_left_out[2] ,
    \cbx_1__1__31_chanx_left_out[3] ,
    \cbx_1__1__31_chanx_left_out[4] ,
    \cbx_1__1__31_chanx_left_out[5] ,
    \cbx_1__1__31_chanx_left_out[6] ,
    \cbx_1__1__31_chanx_left_out[7] ,
    \cbx_1__1__31_chanx_left_out[8] ,
    \cbx_1__1__31_chanx_left_out[9] ,
    \cbx_1__1__31_chanx_left_out[10] ,
    \cbx_1__1__31_chanx_left_out[11] ,
    \cbx_1__1__31_chanx_left_out[12] ,
    \cbx_1__1__31_chanx_left_out[13] ,
    \cbx_1__1__31_chanx_left_out[14] ,
    \cbx_1__1__31_chanx_left_out[15] ,
    \cbx_1__1__31_chanx_left_out[16] ,
    \cbx_1__1__31_chanx_left_out[17] ,
    \cbx_1__1__31_chanx_left_out[18] ,
    \cbx_1__1__31_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__24_chanx_right_out[0] ,
    \sb_1__1__24_chanx_right_out[1] ,
    \sb_1__1__24_chanx_right_out[2] ,
    \sb_1__1__24_chanx_right_out[3] ,
    \sb_1__1__24_chanx_right_out[4] ,
    \sb_1__1__24_chanx_right_out[5] ,
    \sb_1__1__24_chanx_right_out[6] ,
    \sb_1__1__24_chanx_right_out[7] ,
    \sb_1__1__24_chanx_right_out[8] ,
    \sb_1__1__24_chanx_right_out[9] ,
    \sb_1__1__24_chanx_right_out[10] ,
    \sb_1__1__24_chanx_right_out[11] ,
    \sb_1__1__24_chanx_right_out[12] ,
    \sb_1__1__24_chanx_right_out[13] ,
    \sb_1__1__24_chanx_right_out[14] ,
    \sb_1__1__24_chanx_right_out[15] ,
    \sb_1__1__24_chanx_right_out[16] ,
    \sb_1__1__24_chanx_right_out[17] ,
    \sb_1__1__24_chanx_right_out[18] ,
    \sb_1__1__24_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__27_chany_top_out[0] ,
    \cby_1__1__27_chany_top_out[1] ,
    \cby_1__1__27_chany_top_out[2] ,
    \cby_1__1__27_chany_top_out[3] ,
    \cby_1__1__27_chany_top_out[4] ,
    \cby_1__1__27_chany_top_out[5] ,
    \cby_1__1__27_chany_top_out[6] ,
    \cby_1__1__27_chany_top_out[7] ,
    \cby_1__1__27_chany_top_out[8] ,
    \cby_1__1__27_chany_top_out[9] ,
    \cby_1__1__27_chany_top_out[10] ,
    \cby_1__1__27_chany_top_out[11] ,
    \cby_1__1__27_chany_top_out[12] ,
    \cby_1__1__27_chany_top_out[13] ,
    \cby_1__1__27_chany_top_out[14] ,
    \cby_1__1__27_chany_top_out[15] ,
    \cby_1__1__27_chany_top_out[16] ,
    \cby_1__1__27_chany_top_out[17] ,
    \cby_1__1__27_chany_top_out[18] ,
    \cby_1__1__27_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__24_chany_bottom_out[0] ,
    \sb_1__1__24_chany_bottom_out[1] ,
    \sb_1__1__24_chany_bottom_out[2] ,
    \sb_1__1__24_chany_bottom_out[3] ,
    \sb_1__1__24_chany_bottom_out[4] ,
    \sb_1__1__24_chany_bottom_out[5] ,
    \sb_1__1__24_chany_bottom_out[6] ,
    \sb_1__1__24_chany_bottom_out[7] ,
    \sb_1__1__24_chany_bottom_out[8] ,
    \sb_1__1__24_chany_bottom_out[9] ,
    \sb_1__1__24_chany_bottom_out[10] ,
    \sb_1__1__24_chany_bottom_out[11] ,
    \sb_1__1__24_chany_bottom_out[12] ,
    \sb_1__1__24_chany_bottom_out[13] ,
    \sb_1__1__24_chany_bottom_out[14] ,
    \sb_1__1__24_chany_bottom_out[15] ,
    \sb_1__1__24_chany_bottom_out[16] ,
    \sb_1__1__24_chany_bottom_out[17] ,
    \sb_1__1__24_chany_bottom_out[18] ,
    \sb_1__1__24_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__28_chany_bottom_out[0] ,
    \cby_1__1__28_chany_bottom_out[1] ,
    \cby_1__1__28_chany_bottom_out[2] ,
    \cby_1__1__28_chany_bottom_out[3] ,
    \cby_1__1__28_chany_bottom_out[4] ,
    \cby_1__1__28_chany_bottom_out[5] ,
    \cby_1__1__28_chany_bottom_out[6] ,
    \cby_1__1__28_chany_bottom_out[7] ,
    \cby_1__1__28_chany_bottom_out[8] ,
    \cby_1__1__28_chany_bottom_out[9] ,
    \cby_1__1__28_chany_bottom_out[10] ,
    \cby_1__1__28_chany_bottom_out[11] ,
    \cby_1__1__28_chany_bottom_out[12] ,
    \cby_1__1__28_chany_bottom_out[13] ,
    \cby_1__1__28_chany_bottom_out[14] ,
    \cby_1__1__28_chany_bottom_out[15] ,
    \cby_1__1__28_chany_bottom_out[16] ,
    \cby_1__1__28_chany_bottom_out[17] ,
    \cby_1__1__28_chany_bottom_out[18] ,
    \cby_1__1__28_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__24_chany_top_out[0] ,
    \sb_1__1__24_chany_top_out[1] ,
    \sb_1__1__24_chany_top_out[2] ,
    \sb_1__1__24_chany_top_out[3] ,
    \sb_1__1__24_chany_top_out[4] ,
    \sb_1__1__24_chany_top_out[5] ,
    \sb_1__1__24_chany_top_out[6] ,
    \sb_1__1__24_chany_top_out[7] ,
    \sb_1__1__24_chany_top_out[8] ,
    \sb_1__1__24_chany_top_out[9] ,
    \sb_1__1__24_chany_top_out[10] ,
    \sb_1__1__24_chany_top_out[11] ,
    \sb_1__1__24_chany_top_out[12] ,
    \sb_1__1__24_chany_top_out[13] ,
    \sb_1__1__24_chany_top_out[14] ,
    \sb_1__1__24_chany_top_out[15] ,
    \sb_1__1__24_chany_top_out[16] ,
    \sb_1__1__24_chany_top_out[17] ,
    \sb_1__1__24_chany_top_out[18] ,
    \sb_1__1__24_chany_top_out[19] }));
 sb_1__1_ sb_4__5_ (.Test_en_N_out(\Test_enWires[11] ),
    .Test_en_S_in(\Test_enWires[10] ),
    .bottom_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__32_ccff_tail),
    .ccff_tail(sb_1__1__25_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[112] ),
    .right_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__25_chanx_right_out[0] ,
    \cbx_1__1__25_chanx_right_out[1] ,
    \cbx_1__1__25_chanx_right_out[2] ,
    \cbx_1__1__25_chanx_right_out[3] ,
    \cbx_1__1__25_chanx_right_out[4] ,
    \cbx_1__1__25_chanx_right_out[5] ,
    \cbx_1__1__25_chanx_right_out[6] ,
    \cbx_1__1__25_chanx_right_out[7] ,
    \cbx_1__1__25_chanx_right_out[8] ,
    \cbx_1__1__25_chanx_right_out[9] ,
    \cbx_1__1__25_chanx_right_out[10] ,
    \cbx_1__1__25_chanx_right_out[11] ,
    \cbx_1__1__25_chanx_right_out[12] ,
    \cbx_1__1__25_chanx_right_out[13] ,
    \cbx_1__1__25_chanx_right_out[14] ,
    \cbx_1__1__25_chanx_right_out[15] ,
    \cbx_1__1__25_chanx_right_out[16] ,
    \cbx_1__1__25_chanx_right_out[17] ,
    \cbx_1__1__25_chanx_right_out[18] ,
    \cbx_1__1__25_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__25_chanx_left_out[0] ,
    \sb_1__1__25_chanx_left_out[1] ,
    \sb_1__1__25_chanx_left_out[2] ,
    \sb_1__1__25_chanx_left_out[3] ,
    \sb_1__1__25_chanx_left_out[4] ,
    \sb_1__1__25_chanx_left_out[5] ,
    \sb_1__1__25_chanx_left_out[6] ,
    \sb_1__1__25_chanx_left_out[7] ,
    \sb_1__1__25_chanx_left_out[8] ,
    \sb_1__1__25_chanx_left_out[9] ,
    \sb_1__1__25_chanx_left_out[10] ,
    \sb_1__1__25_chanx_left_out[11] ,
    \sb_1__1__25_chanx_left_out[12] ,
    \sb_1__1__25_chanx_left_out[13] ,
    \sb_1__1__25_chanx_left_out[14] ,
    \sb_1__1__25_chanx_left_out[15] ,
    \sb_1__1__25_chanx_left_out[16] ,
    \sb_1__1__25_chanx_left_out[17] ,
    \sb_1__1__25_chanx_left_out[18] ,
    \sb_1__1__25_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__32_chanx_left_out[0] ,
    \cbx_1__1__32_chanx_left_out[1] ,
    \cbx_1__1__32_chanx_left_out[2] ,
    \cbx_1__1__32_chanx_left_out[3] ,
    \cbx_1__1__32_chanx_left_out[4] ,
    \cbx_1__1__32_chanx_left_out[5] ,
    \cbx_1__1__32_chanx_left_out[6] ,
    \cbx_1__1__32_chanx_left_out[7] ,
    \cbx_1__1__32_chanx_left_out[8] ,
    \cbx_1__1__32_chanx_left_out[9] ,
    \cbx_1__1__32_chanx_left_out[10] ,
    \cbx_1__1__32_chanx_left_out[11] ,
    \cbx_1__1__32_chanx_left_out[12] ,
    \cbx_1__1__32_chanx_left_out[13] ,
    \cbx_1__1__32_chanx_left_out[14] ,
    \cbx_1__1__32_chanx_left_out[15] ,
    \cbx_1__1__32_chanx_left_out[16] ,
    \cbx_1__1__32_chanx_left_out[17] ,
    \cbx_1__1__32_chanx_left_out[18] ,
    \cbx_1__1__32_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__25_chanx_right_out[0] ,
    \sb_1__1__25_chanx_right_out[1] ,
    \sb_1__1__25_chanx_right_out[2] ,
    \sb_1__1__25_chanx_right_out[3] ,
    \sb_1__1__25_chanx_right_out[4] ,
    \sb_1__1__25_chanx_right_out[5] ,
    \sb_1__1__25_chanx_right_out[6] ,
    \sb_1__1__25_chanx_right_out[7] ,
    \sb_1__1__25_chanx_right_out[8] ,
    \sb_1__1__25_chanx_right_out[9] ,
    \sb_1__1__25_chanx_right_out[10] ,
    \sb_1__1__25_chanx_right_out[11] ,
    \sb_1__1__25_chanx_right_out[12] ,
    \sb_1__1__25_chanx_right_out[13] ,
    \sb_1__1__25_chanx_right_out[14] ,
    \sb_1__1__25_chanx_right_out[15] ,
    \sb_1__1__25_chanx_right_out[16] ,
    \sb_1__1__25_chanx_right_out[17] ,
    \sb_1__1__25_chanx_right_out[18] ,
    \sb_1__1__25_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__28_chany_top_out[0] ,
    \cby_1__1__28_chany_top_out[1] ,
    \cby_1__1__28_chany_top_out[2] ,
    \cby_1__1__28_chany_top_out[3] ,
    \cby_1__1__28_chany_top_out[4] ,
    \cby_1__1__28_chany_top_out[5] ,
    \cby_1__1__28_chany_top_out[6] ,
    \cby_1__1__28_chany_top_out[7] ,
    \cby_1__1__28_chany_top_out[8] ,
    \cby_1__1__28_chany_top_out[9] ,
    \cby_1__1__28_chany_top_out[10] ,
    \cby_1__1__28_chany_top_out[11] ,
    \cby_1__1__28_chany_top_out[12] ,
    \cby_1__1__28_chany_top_out[13] ,
    \cby_1__1__28_chany_top_out[14] ,
    \cby_1__1__28_chany_top_out[15] ,
    \cby_1__1__28_chany_top_out[16] ,
    \cby_1__1__28_chany_top_out[17] ,
    \cby_1__1__28_chany_top_out[18] ,
    \cby_1__1__28_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__25_chany_bottom_out[0] ,
    \sb_1__1__25_chany_bottom_out[1] ,
    \sb_1__1__25_chany_bottom_out[2] ,
    \sb_1__1__25_chany_bottom_out[3] ,
    \sb_1__1__25_chany_bottom_out[4] ,
    \sb_1__1__25_chany_bottom_out[5] ,
    \sb_1__1__25_chany_bottom_out[6] ,
    \sb_1__1__25_chany_bottom_out[7] ,
    \sb_1__1__25_chany_bottom_out[8] ,
    \sb_1__1__25_chany_bottom_out[9] ,
    \sb_1__1__25_chany_bottom_out[10] ,
    \sb_1__1__25_chany_bottom_out[11] ,
    \sb_1__1__25_chany_bottom_out[12] ,
    \sb_1__1__25_chany_bottom_out[13] ,
    \sb_1__1__25_chany_bottom_out[14] ,
    \sb_1__1__25_chany_bottom_out[15] ,
    \sb_1__1__25_chany_bottom_out[16] ,
    \sb_1__1__25_chany_bottom_out[17] ,
    \sb_1__1__25_chany_bottom_out[18] ,
    \sb_1__1__25_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__29_chany_bottom_out[0] ,
    \cby_1__1__29_chany_bottom_out[1] ,
    \cby_1__1__29_chany_bottom_out[2] ,
    \cby_1__1__29_chany_bottom_out[3] ,
    \cby_1__1__29_chany_bottom_out[4] ,
    \cby_1__1__29_chany_bottom_out[5] ,
    \cby_1__1__29_chany_bottom_out[6] ,
    \cby_1__1__29_chany_bottom_out[7] ,
    \cby_1__1__29_chany_bottom_out[8] ,
    \cby_1__1__29_chany_bottom_out[9] ,
    \cby_1__1__29_chany_bottom_out[10] ,
    \cby_1__1__29_chany_bottom_out[11] ,
    \cby_1__1__29_chany_bottom_out[12] ,
    \cby_1__1__29_chany_bottom_out[13] ,
    \cby_1__1__29_chany_bottom_out[14] ,
    \cby_1__1__29_chany_bottom_out[15] ,
    \cby_1__1__29_chany_bottom_out[16] ,
    \cby_1__1__29_chany_bottom_out[17] ,
    \cby_1__1__29_chany_bottom_out[18] ,
    \cby_1__1__29_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__25_chany_top_out[0] ,
    \sb_1__1__25_chany_top_out[1] ,
    \sb_1__1__25_chany_top_out[2] ,
    \sb_1__1__25_chany_top_out[3] ,
    \sb_1__1__25_chany_top_out[4] ,
    \sb_1__1__25_chany_top_out[5] ,
    \sb_1__1__25_chany_top_out[6] ,
    \sb_1__1__25_chany_top_out[7] ,
    \sb_1__1__25_chany_top_out[8] ,
    \sb_1__1__25_chany_top_out[9] ,
    \sb_1__1__25_chany_top_out[10] ,
    \sb_1__1__25_chany_top_out[11] ,
    \sb_1__1__25_chany_top_out[12] ,
    \sb_1__1__25_chany_top_out[13] ,
    \sb_1__1__25_chany_top_out[14] ,
    \sb_1__1__25_chany_top_out[15] ,
    \sb_1__1__25_chany_top_out[16] ,
    \sb_1__1__25_chany_top_out[17] ,
    \sb_1__1__25_chany_top_out[18] ,
    \sb_1__1__25_chany_top_out[19] }));
 sb_1__1_ sb_4__6_ (.Test_en_N_out(\Test_enWires[13] ),
    .Test_en_S_in(\Test_enWires[12] ),
    .bottom_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__33_ccff_tail),
    .ccff_tail(sb_1__1__26_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[115] ),
    .right_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__26_chanx_right_out[0] ,
    \cbx_1__1__26_chanx_right_out[1] ,
    \cbx_1__1__26_chanx_right_out[2] ,
    \cbx_1__1__26_chanx_right_out[3] ,
    \cbx_1__1__26_chanx_right_out[4] ,
    \cbx_1__1__26_chanx_right_out[5] ,
    \cbx_1__1__26_chanx_right_out[6] ,
    \cbx_1__1__26_chanx_right_out[7] ,
    \cbx_1__1__26_chanx_right_out[8] ,
    \cbx_1__1__26_chanx_right_out[9] ,
    \cbx_1__1__26_chanx_right_out[10] ,
    \cbx_1__1__26_chanx_right_out[11] ,
    \cbx_1__1__26_chanx_right_out[12] ,
    \cbx_1__1__26_chanx_right_out[13] ,
    \cbx_1__1__26_chanx_right_out[14] ,
    \cbx_1__1__26_chanx_right_out[15] ,
    \cbx_1__1__26_chanx_right_out[16] ,
    \cbx_1__1__26_chanx_right_out[17] ,
    \cbx_1__1__26_chanx_right_out[18] ,
    \cbx_1__1__26_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__26_chanx_left_out[0] ,
    \sb_1__1__26_chanx_left_out[1] ,
    \sb_1__1__26_chanx_left_out[2] ,
    \sb_1__1__26_chanx_left_out[3] ,
    \sb_1__1__26_chanx_left_out[4] ,
    \sb_1__1__26_chanx_left_out[5] ,
    \sb_1__1__26_chanx_left_out[6] ,
    \sb_1__1__26_chanx_left_out[7] ,
    \sb_1__1__26_chanx_left_out[8] ,
    \sb_1__1__26_chanx_left_out[9] ,
    \sb_1__1__26_chanx_left_out[10] ,
    \sb_1__1__26_chanx_left_out[11] ,
    \sb_1__1__26_chanx_left_out[12] ,
    \sb_1__1__26_chanx_left_out[13] ,
    \sb_1__1__26_chanx_left_out[14] ,
    \sb_1__1__26_chanx_left_out[15] ,
    \sb_1__1__26_chanx_left_out[16] ,
    \sb_1__1__26_chanx_left_out[17] ,
    \sb_1__1__26_chanx_left_out[18] ,
    \sb_1__1__26_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__33_chanx_left_out[0] ,
    \cbx_1__1__33_chanx_left_out[1] ,
    \cbx_1__1__33_chanx_left_out[2] ,
    \cbx_1__1__33_chanx_left_out[3] ,
    \cbx_1__1__33_chanx_left_out[4] ,
    \cbx_1__1__33_chanx_left_out[5] ,
    \cbx_1__1__33_chanx_left_out[6] ,
    \cbx_1__1__33_chanx_left_out[7] ,
    \cbx_1__1__33_chanx_left_out[8] ,
    \cbx_1__1__33_chanx_left_out[9] ,
    \cbx_1__1__33_chanx_left_out[10] ,
    \cbx_1__1__33_chanx_left_out[11] ,
    \cbx_1__1__33_chanx_left_out[12] ,
    \cbx_1__1__33_chanx_left_out[13] ,
    \cbx_1__1__33_chanx_left_out[14] ,
    \cbx_1__1__33_chanx_left_out[15] ,
    \cbx_1__1__33_chanx_left_out[16] ,
    \cbx_1__1__33_chanx_left_out[17] ,
    \cbx_1__1__33_chanx_left_out[18] ,
    \cbx_1__1__33_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__26_chanx_right_out[0] ,
    \sb_1__1__26_chanx_right_out[1] ,
    \sb_1__1__26_chanx_right_out[2] ,
    \sb_1__1__26_chanx_right_out[3] ,
    \sb_1__1__26_chanx_right_out[4] ,
    \sb_1__1__26_chanx_right_out[5] ,
    \sb_1__1__26_chanx_right_out[6] ,
    \sb_1__1__26_chanx_right_out[7] ,
    \sb_1__1__26_chanx_right_out[8] ,
    \sb_1__1__26_chanx_right_out[9] ,
    \sb_1__1__26_chanx_right_out[10] ,
    \sb_1__1__26_chanx_right_out[11] ,
    \sb_1__1__26_chanx_right_out[12] ,
    \sb_1__1__26_chanx_right_out[13] ,
    \sb_1__1__26_chanx_right_out[14] ,
    \sb_1__1__26_chanx_right_out[15] ,
    \sb_1__1__26_chanx_right_out[16] ,
    \sb_1__1__26_chanx_right_out[17] ,
    \sb_1__1__26_chanx_right_out[18] ,
    \sb_1__1__26_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__29_chany_top_out[0] ,
    \cby_1__1__29_chany_top_out[1] ,
    \cby_1__1__29_chany_top_out[2] ,
    \cby_1__1__29_chany_top_out[3] ,
    \cby_1__1__29_chany_top_out[4] ,
    \cby_1__1__29_chany_top_out[5] ,
    \cby_1__1__29_chany_top_out[6] ,
    \cby_1__1__29_chany_top_out[7] ,
    \cby_1__1__29_chany_top_out[8] ,
    \cby_1__1__29_chany_top_out[9] ,
    \cby_1__1__29_chany_top_out[10] ,
    \cby_1__1__29_chany_top_out[11] ,
    \cby_1__1__29_chany_top_out[12] ,
    \cby_1__1__29_chany_top_out[13] ,
    \cby_1__1__29_chany_top_out[14] ,
    \cby_1__1__29_chany_top_out[15] ,
    \cby_1__1__29_chany_top_out[16] ,
    \cby_1__1__29_chany_top_out[17] ,
    \cby_1__1__29_chany_top_out[18] ,
    \cby_1__1__29_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__26_chany_bottom_out[0] ,
    \sb_1__1__26_chany_bottom_out[1] ,
    \sb_1__1__26_chany_bottom_out[2] ,
    \sb_1__1__26_chany_bottom_out[3] ,
    \sb_1__1__26_chany_bottom_out[4] ,
    \sb_1__1__26_chany_bottom_out[5] ,
    \sb_1__1__26_chany_bottom_out[6] ,
    \sb_1__1__26_chany_bottom_out[7] ,
    \sb_1__1__26_chany_bottom_out[8] ,
    \sb_1__1__26_chany_bottom_out[9] ,
    \sb_1__1__26_chany_bottom_out[10] ,
    \sb_1__1__26_chany_bottom_out[11] ,
    \sb_1__1__26_chany_bottom_out[12] ,
    \sb_1__1__26_chany_bottom_out[13] ,
    \sb_1__1__26_chany_bottom_out[14] ,
    \sb_1__1__26_chany_bottom_out[15] ,
    \sb_1__1__26_chany_bottom_out[16] ,
    \sb_1__1__26_chany_bottom_out[17] ,
    \sb_1__1__26_chany_bottom_out[18] ,
    \sb_1__1__26_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__30_chany_bottom_out[0] ,
    \cby_1__1__30_chany_bottom_out[1] ,
    \cby_1__1__30_chany_bottom_out[2] ,
    \cby_1__1__30_chany_bottom_out[3] ,
    \cby_1__1__30_chany_bottom_out[4] ,
    \cby_1__1__30_chany_bottom_out[5] ,
    \cby_1__1__30_chany_bottom_out[6] ,
    \cby_1__1__30_chany_bottom_out[7] ,
    \cby_1__1__30_chany_bottom_out[8] ,
    \cby_1__1__30_chany_bottom_out[9] ,
    \cby_1__1__30_chany_bottom_out[10] ,
    \cby_1__1__30_chany_bottom_out[11] ,
    \cby_1__1__30_chany_bottom_out[12] ,
    \cby_1__1__30_chany_bottom_out[13] ,
    \cby_1__1__30_chany_bottom_out[14] ,
    \cby_1__1__30_chany_bottom_out[15] ,
    \cby_1__1__30_chany_bottom_out[16] ,
    \cby_1__1__30_chany_bottom_out[17] ,
    \cby_1__1__30_chany_bottom_out[18] ,
    \cby_1__1__30_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__26_chany_top_out[0] ,
    \sb_1__1__26_chany_top_out[1] ,
    \sb_1__1__26_chany_top_out[2] ,
    \sb_1__1__26_chany_top_out[3] ,
    \sb_1__1__26_chany_top_out[4] ,
    \sb_1__1__26_chany_top_out[5] ,
    \sb_1__1__26_chany_top_out[6] ,
    \sb_1__1__26_chany_top_out[7] ,
    \sb_1__1__26_chany_top_out[8] ,
    \sb_1__1__26_chany_top_out[9] ,
    \sb_1__1__26_chany_top_out[10] ,
    \sb_1__1__26_chany_top_out[11] ,
    \sb_1__1__26_chany_top_out[12] ,
    \sb_1__1__26_chany_top_out[13] ,
    \sb_1__1__26_chany_top_out[14] ,
    \sb_1__1__26_chany_top_out[15] ,
    \sb_1__1__26_chany_top_out[16] ,
    \sb_1__1__26_chany_top_out[17] ,
    \sb_1__1__26_chany_top_out[18] ,
    \sb_1__1__26_chany_top_out[19] }));
 sb_1__1_ sb_4__7_ (.Test_en_N_out(\Test_enWires[15] ),
    .Test_en_S_in(\Test_enWires[14] ),
    .bottom_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__34_ccff_tail),
    .ccff_tail(sb_1__1__27_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[118] ),
    .right_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__27_chanx_right_out[0] ,
    \cbx_1__1__27_chanx_right_out[1] ,
    \cbx_1__1__27_chanx_right_out[2] ,
    \cbx_1__1__27_chanx_right_out[3] ,
    \cbx_1__1__27_chanx_right_out[4] ,
    \cbx_1__1__27_chanx_right_out[5] ,
    \cbx_1__1__27_chanx_right_out[6] ,
    \cbx_1__1__27_chanx_right_out[7] ,
    \cbx_1__1__27_chanx_right_out[8] ,
    \cbx_1__1__27_chanx_right_out[9] ,
    \cbx_1__1__27_chanx_right_out[10] ,
    \cbx_1__1__27_chanx_right_out[11] ,
    \cbx_1__1__27_chanx_right_out[12] ,
    \cbx_1__1__27_chanx_right_out[13] ,
    \cbx_1__1__27_chanx_right_out[14] ,
    \cbx_1__1__27_chanx_right_out[15] ,
    \cbx_1__1__27_chanx_right_out[16] ,
    \cbx_1__1__27_chanx_right_out[17] ,
    \cbx_1__1__27_chanx_right_out[18] ,
    \cbx_1__1__27_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__27_chanx_left_out[0] ,
    \sb_1__1__27_chanx_left_out[1] ,
    \sb_1__1__27_chanx_left_out[2] ,
    \sb_1__1__27_chanx_left_out[3] ,
    \sb_1__1__27_chanx_left_out[4] ,
    \sb_1__1__27_chanx_left_out[5] ,
    \sb_1__1__27_chanx_left_out[6] ,
    \sb_1__1__27_chanx_left_out[7] ,
    \sb_1__1__27_chanx_left_out[8] ,
    \sb_1__1__27_chanx_left_out[9] ,
    \sb_1__1__27_chanx_left_out[10] ,
    \sb_1__1__27_chanx_left_out[11] ,
    \sb_1__1__27_chanx_left_out[12] ,
    \sb_1__1__27_chanx_left_out[13] ,
    \sb_1__1__27_chanx_left_out[14] ,
    \sb_1__1__27_chanx_left_out[15] ,
    \sb_1__1__27_chanx_left_out[16] ,
    \sb_1__1__27_chanx_left_out[17] ,
    \sb_1__1__27_chanx_left_out[18] ,
    \sb_1__1__27_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__34_chanx_left_out[0] ,
    \cbx_1__1__34_chanx_left_out[1] ,
    \cbx_1__1__34_chanx_left_out[2] ,
    \cbx_1__1__34_chanx_left_out[3] ,
    \cbx_1__1__34_chanx_left_out[4] ,
    \cbx_1__1__34_chanx_left_out[5] ,
    \cbx_1__1__34_chanx_left_out[6] ,
    \cbx_1__1__34_chanx_left_out[7] ,
    \cbx_1__1__34_chanx_left_out[8] ,
    \cbx_1__1__34_chanx_left_out[9] ,
    \cbx_1__1__34_chanx_left_out[10] ,
    \cbx_1__1__34_chanx_left_out[11] ,
    \cbx_1__1__34_chanx_left_out[12] ,
    \cbx_1__1__34_chanx_left_out[13] ,
    \cbx_1__1__34_chanx_left_out[14] ,
    \cbx_1__1__34_chanx_left_out[15] ,
    \cbx_1__1__34_chanx_left_out[16] ,
    \cbx_1__1__34_chanx_left_out[17] ,
    \cbx_1__1__34_chanx_left_out[18] ,
    \cbx_1__1__34_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__27_chanx_right_out[0] ,
    \sb_1__1__27_chanx_right_out[1] ,
    \sb_1__1__27_chanx_right_out[2] ,
    \sb_1__1__27_chanx_right_out[3] ,
    \sb_1__1__27_chanx_right_out[4] ,
    \sb_1__1__27_chanx_right_out[5] ,
    \sb_1__1__27_chanx_right_out[6] ,
    \sb_1__1__27_chanx_right_out[7] ,
    \sb_1__1__27_chanx_right_out[8] ,
    \sb_1__1__27_chanx_right_out[9] ,
    \sb_1__1__27_chanx_right_out[10] ,
    \sb_1__1__27_chanx_right_out[11] ,
    \sb_1__1__27_chanx_right_out[12] ,
    \sb_1__1__27_chanx_right_out[13] ,
    \sb_1__1__27_chanx_right_out[14] ,
    \sb_1__1__27_chanx_right_out[15] ,
    \sb_1__1__27_chanx_right_out[16] ,
    \sb_1__1__27_chanx_right_out[17] ,
    \sb_1__1__27_chanx_right_out[18] ,
    \sb_1__1__27_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__30_chany_top_out[0] ,
    \cby_1__1__30_chany_top_out[1] ,
    \cby_1__1__30_chany_top_out[2] ,
    \cby_1__1__30_chany_top_out[3] ,
    \cby_1__1__30_chany_top_out[4] ,
    \cby_1__1__30_chany_top_out[5] ,
    \cby_1__1__30_chany_top_out[6] ,
    \cby_1__1__30_chany_top_out[7] ,
    \cby_1__1__30_chany_top_out[8] ,
    \cby_1__1__30_chany_top_out[9] ,
    \cby_1__1__30_chany_top_out[10] ,
    \cby_1__1__30_chany_top_out[11] ,
    \cby_1__1__30_chany_top_out[12] ,
    \cby_1__1__30_chany_top_out[13] ,
    \cby_1__1__30_chany_top_out[14] ,
    \cby_1__1__30_chany_top_out[15] ,
    \cby_1__1__30_chany_top_out[16] ,
    \cby_1__1__30_chany_top_out[17] ,
    \cby_1__1__30_chany_top_out[18] ,
    \cby_1__1__30_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__27_chany_bottom_out[0] ,
    \sb_1__1__27_chany_bottom_out[1] ,
    \sb_1__1__27_chany_bottom_out[2] ,
    \sb_1__1__27_chany_bottom_out[3] ,
    \sb_1__1__27_chany_bottom_out[4] ,
    \sb_1__1__27_chany_bottom_out[5] ,
    \sb_1__1__27_chany_bottom_out[6] ,
    \sb_1__1__27_chany_bottom_out[7] ,
    \sb_1__1__27_chany_bottom_out[8] ,
    \sb_1__1__27_chany_bottom_out[9] ,
    \sb_1__1__27_chany_bottom_out[10] ,
    \sb_1__1__27_chany_bottom_out[11] ,
    \sb_1__1__27_chany_bottom_out[12] ,
    \sb_1__1__27_chany_bottom_out[13] ,
    \sb_1__1__27_chany_bottom_out[14] ,
    \sb_1__1__27_chany_bottom_out[15] ,
    \sb_1__1__27_chany_bottom_out[16] ,
    \sb_1__1__27_chany_bottom_out[17] ,
    \sb_1__1__27_chany_bottom_out[18] ,
    \sb_1__1__27_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__31_chany_bottom_out[0] ,
    \cby_1__1__31_chany_bottom_out[1] ,
    \cby_1__1__31_chany_bottom_out[2] ,
    \cby_1__1__31_chany_bottom_out[3] ,
    \cby_1__1__31_chany_bottom_out[4] ,
    \cby_1__1__31_chany_bottom_out[5] ,
    \cby_1__1__31_chany_bottom_out[6] ,
    \cby_1__1__31_chany_bottom_out[7] ,
    \cby_1__1__31_chany_bottom_out[8] ,
    \cby_1__1__31_chany_bottom_out[9] ,
    \cby_1__1__31_chany_bottom_out[10] ,
    \cby_1__1__31_chany_bottom_out[11] ,
    \cby_1__1__31_chany_bottom_out[12] ,
    \cby_1__1__31_chany_bottom_out[13] ,
    \cby_1__1__31_chany_bottom_out[14] ,
    \cby_1__1__31_chany_bottom_out[15] ,
    \cby_1__1__31_chany_bottom_out[16] ,
    \cby_1__1__31_chany_bottom_out[17] ,
    \cby_1__1__31_chany_bottom_out[18] ,
    \cby_1__1__31_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__27_chany_top_out[0] ,
    \sb_1__1__27_chany_top_out[1] ,
    \sb_1__1__27_chany_top_out[2] ,
    \sb_1__1__27_chany_top_out[3] ,
    \sb_1__1__27_chany_top_out[4] ,
    \sb_1__1__27_chany_top_out[5] ,
    \sb_1__1__27_chany_top_out[6] ,
    \sb_1__1__27_chany_top_out[7] ,
    \sb_1__1__27_chany_top_out[8] ,
    \sb_1__1__27_chany_top_out[9] ,
    \sb_1__1__27_chany_top_out[10] ,
    \sb_1__1__27_chany_top_out[11] ,
    \sb_1__1__27_chany_top_out[12] ,
    \sb_1__1__27_chany_top_out[13] ,
    \sb_1__1__27_chany_top_out[14] ,
    \sb_1__1__27_chany_top_out[15] ,
    \sb_1__1__27_chany_top_out[16] ,
    \sb_1__1__27_chany_top_out[17] ,
    \sb_1__1__27_chany_top_out[18] ,
    \sb_1__1__27_chany_top_out[19] }));
 sb_1__2_ sb_4__8_ (.SC_IN_BOT(\scff_Wires[73] ),
    .SC_OUT_BOT(\scff_Wires[74] ),
    .bottom_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_upper),
    .ccff_head(grid_io_top_4_ccff_tail),
    .ccff_tail(sb_1__8__3_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[120] ),
    .right_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__3_chanx_right_out[0] ,
    \cbx_1__8__3_chanx_right_out[1] ,
    \cbx_1__8__3_chanx_right_out[2] ,
    \cbx_1__8__3_chanx_right_out[3] ,
    \cbx_1__8__3_chanx_right_out[4] ,
    \cbx_1__8__3_chanx_right_out[5] ,
    \cbx_1__8__3_chanx_right_out[6] ,
    \cbx_1__8__3_chanx_right_out[7] ,
    \cbx_1__8__3_chanx_right_out[8] ,
    \cbx_1__8__3_chanx_right_out[9] ,
    \cbx_1__8__3_chanx_right_out[10] ,
    \cbx_1__8__3_chanx_right_out[11] ,
    \cbx_1__8__3_chanx_right_out[12] ,
    \cbx_1__8__3_chanx_right_out[13] ,
    \cbx_1__8__3_chanx_right_out[14] ,
    \cbx_1__8__3_chanx_right_out[15] ,
    \cbx_1__8__3_chanx_right_out[16] ,
    \cbx_1__8__3_chanx_right_out[17] ,
    \cbx_1__8__3_chanx_right_out[18] ,
    \cbx_1__8__3_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__8__3_chanx_left_out[0] ,
    \sb_1__8__3_chanx_left_out[1] ,
    \sb_1__8__3_chanx_left_out[2] ,
    \sb_1__8__3_chanx_left_out[3] ,
    \sb_1__8__3_chanx_left_out[4] ,
    \sb_1__8__3_chanx_left_out[5] ,
    \sb_1__8__3_chanx_left_out[6] ,
    \sb_1__8__3_chanx_left_out[7] ,
    \sb_1__8__3_chanx_left_out[8] ,
    \sb_1__8__3_chanx_left_out[9] ,
    \sb_1__8__3_chanx_left_out[10] ,
    \sb_1__8__3_chanx_left_out[11] ,
    \sb_1__8__3_chanx_left_out[12] ,
    \sb_1__8__3_chanx_left_out[13] ,
    \sb_1__8__3_chanx_left_out[14] ,
    \sb_1__8__3_chanx_left_out[15] ,
    \sb_1__8__3_chanx_left_out[16] ,
    \sb_1__8__3_chanx_left_out[17] ,
    \sb_1__8__3_chanx_left_out[18] ,
    \sb_1__8__3_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__8__4_chanx_left_out[0] ,
    \cbx_1__8__4_chanx_left_out[1] ,
    \cbx_1__8__4_chanx_left_out[2] ,
    \cbx_1__8__4_chanx_left_out[3] ,
    \cbx_1__8__4_chanx_left_out[4] ,
    \cbx_1__8__4_chanx_left_out[5] ,
    \cbx_1__8__4_chanx_left_out[6] ,
    \cbx_1__8__4_chanx_left_out[7] ,
    \cbx_1__8__4_chanx_left_out[8] ,
    \cbx_1__8__4_chanx_left_out[9] ,
    \cbx_1__8__4_chanx_left_out[10] ,
    \cbx_1__8__4_chanx_left_out[11] ,
    \cbx_1__8__4_chanx_left_out[12] ,
    \cbx_1__8__4_chanx_left_out[13] ,
    \cbx_1__8__4_chanx_left_out[14] ,
    \cbx_1__8__4_chanx_left_out[15] ,
    \cbx_1__8__4_chanx_left_out[16] ,
    \cbx_1__8__4_chanx_left_out[17] ,
    \cbx_1__8__4_chanx_left_out[18] ,
    \cbx_1__8__4_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__8__3_chanx_right_out[0] ,
    \sb_1__8__3_chanx_right_out[1] ,
    \sb_1__8__3_chanx_right_out[2] ,
    \sb_1__8__3_chanx_right_out[3] ,
    \sb_1__8__3_chanx_right_out[4] ,
    \sb_1__8__3_chanx_right_out[5] ,
    \sb_1__8__3_chanx_right_out[6] ,
    \sb_1__8__3_chanx_right_out[7] ,
    \sb_1__8__3_chanx_right_out[8] ,
    \sb_1__8__3_chanx_right_out[9] ,
    \sb_1__8__3_chanx_right_out[10] ,
    \sb_1__8__3_chanx_right_out[11] ,
    \sb_1__8__3_chanx_right_out[12] ,
    \sb_1__8__3_chanx_right_out[13] ,
    \sb_1__8__3_chanx_right_out[14] ,
    \sb_1__8__3_chanx_right_out[15] ,
    \sb_1__8__3_chanx_right_out[16] ,
    \sb_1__8__3_chanx_right_out[17] ,
    \sb_1__8__3_chanx_right_out[18] ,
    \sb_1__8__3_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__31_chany_top_out[0] ,
    \cby_1__1__31_chany_top_out[1] ,
    \cby_1__1__31_chany_top_out[2] ,
    \cby_1__1__31_chany_top_out[3] ,
    \cby_1__1__31_chany_top_out[4] ,
    \cby_1__1__31_chany_top_out[5] ,
    \cby_1__1__31_chany_top_out[6] ,
    \cby_1__1__31_chany_top_out[7] ,
    \cby_1__1__31_chany_top_out[8] ,
    \cby_1__1__31_chany_top_out[9] ,
    \cby_1__1__31_chany_top_out[10] ,
    \cby_1__1__31_chany_top_out[11] ,
    \cby_1__1__31_chany_top_out[12] ,
    \cby_1__1__31_chany_top_out[13] ,
    \cby_1__1__31_chany_top_out[14] ,
    \cby_1__1__31_chany_top_out[15] ,
    \cby_1__1__31_chany_top_out[16] ,
    \cby_1__1__31_chany_top_out[17] ,
    \cby_1__1__31_chany_top_out[18] ,
    \cby_1__1__31_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__8__3_chany_bottom_out[0] ,
    \sb_1__8__3_chany_bottom_out[1] ,
    \sb_1__8__3_chany_bottom_out[2] ,
    \sb_1__8__3_chany_bottom_out[3] ,
    \sb_1__8__3_chany_bottom_out[4] ,
    \sb_1__8__3_chany_bottom_out[5] ,
    \sb_1__8__3_chany_bottom_out[6] ,
    \sb_1__8__3_chany_bottom_out[7] ,
    \sb_1__8__3_chany_bottom_out[8] ,
    \sb_1__8__3_chany_bottom_out[9] ,
    \sb_1__8__3_chany_bottom_out[10] ,
    \sb_1__8__3_chany_bottom_out[11] ,
    \sb_1__8__3_chany_bottom_out[12] ,
    \sb_1__8__3_chany_bottom_out[13] ,
    \sb_1__8__3_chany_bottom_out[14] ,
    \sb_1__8__3_chany_bottom_out[15] ,
    \sb_1__8__3_chany_bottom_out[16] ,
    \sb_1__8__3_chany_bottom_out[17] ,
    \sb_1__8__3_chany_bottom_out[18] ,
    \sb_1__8__3_chany_bottom_out[19] }));
 sb_1__0_ sb_5__0_ (.SC_IN_TOP(\scff_Wires[92] ),
    .SC_OUT_TOP(\scff_Wires[93] ),
    .ccff_head(grid_io_bottom_2_ccff_tail),
    .ccff_tail(sb_1__0__4_ccff_tail),
    .left_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[123] ),
    .right_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__4_chanx_right_out[0] ,
    \cbx_1__0__4_chanx_right_out[1] ,
    \cbx_1__0__4_chanx_right_out[2] ,
    \cbx_1__0__4_chanx_right_out[3] ,
    \cbx_1__0__4_chanx_right_out[4] ,
    \cbx_1__0__4_chanx_right_out[5] ,
    \cbx_1__0__4_chanx_right_out[6] ,
    \cbx_1__0__4_chanx_right_out[7] ,
    \cbx_1__0__4_chanx_right_out[8] ,
    \cbx_1__0__4_chanx_right_out[9] ,
    \cbx_1__0__4_chanx_right_out[10] ,
    \cbx_1__0__4_chanx_right_out[11] ,
    \cbx_1__0__4_chanx_right_out[12] ,
    \cbx_1__0__4_chanx_right_out[13] ,
    \cbx_1__0__4_chanx_right_out[14] ,
    \cbx_1__0__4_chanx_right_out[15] ,
    \cbx_1__0__4_chanx_right_out[16] ,
    \cbx_1__0__4_chanx_right_out[17] ,
    \cbx_1__0__4_chanx_right_out[18] ,
    \cbx_1__0__4_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__0__4_chanx_left_out[0] ,
    \sb_1__0__4_chanx_left_out[1] ,
    \sb_1__0__4_chanx_left_out[2] ,
    \sb_1__0__4_chanx_left_out[3] ,
    \sb_1__0__4_chanx_left_out[4] ,
    \sb_1__0__4_chanx_left_out[5] ,
    \sb_1__0__4_chanx_left_out[6] ,
    \sb_1__0__4_chanx_left_out[7] ,
    \sb_1__0__4_chanx_left_out[8] ,
    \sb_1__0__4_chanx_left_out[9] ,
    \sb_1__0__4_chanx_left_out[10] ,
    \sb_1__0__4_chanx_left_out[11] ,
    \sb_1__0__4_chanx_left_out[12] ,
    \sb_1__0__4_chanx_left_out[13] ,
    \sb_1__0__4_chanx_left_out[14] ,
    \sb_1__0__4_chanx_left_out[15] ,
    \sb_1__0__4_chanx_left_out[16] ,
    \sb_1__0__4_chanx_left_out[17] ,
    \sb_1__0__4_chanx_left_out[18] ,
    \sb_1__0__4_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__0__5_chanx_left_out[0] ,
    \cbx_1__0__5_chanx_left_out[1] ,
    \cbx_1__0__5_chanx_left_out[2] ,
    \cbx_1__0__5_chanx_left_out[3] ,
    \cbx_1__0__5_chanx_left_out[4] ,
    \cbx_1__0__5_chanx_left_out[5] ,
    \cbx_1__0__5_chanx_left_out[6] ,
    \cbx_1__0__5_chanx_left_out[7] ,
    \cbx_1__0__5_chanx_left_out[8] ,
    \cbx_1__0__5_chanx_left_out[9] ,
    \cbx_1__0__5_chanx_left_out[10] ,
    \cbx_1__0__5_chanx_left_out[11] ,
    \cbx_1__0__5_chanx_left_out[12] ,
    \cbx_1__0__5_chanx_left_out[13] ,
    \cbx_1__0__5_chanx_left_out[14] ,
    \cbx_1__0__5_chanx_left_out[15] ,
    \cbx_1__0__5_chanx_left_out[16] ,
    \cbx_1__0__5_chanx_left_out[17] ,
    \cbx_1__0__5_chanx_left_out[18] ,
    \cbx_1__0__5_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__0__4_chanx_right_out[0] ,
    \sb_1__0__4_chanx_right_out[1] ,
    \sb_1__0__4_chanx_right_out[2] ,
    \sb_1__0__4_chanx_right_out[3] ,
    \sb_1__0__4_chanx_right_out[4] ,
    \sb_1__0__4_chanx_right_out[5] ,
    \sb_1__0__4_chanx_right_out[6] ,
    \sb_1__0__4_chanx_right_out[7] ,
    \sb_1__0__4_chanx_right_out[8] ,
    \sb_1__0__4_chanx_right_out[9] ,
    \sb_1__0__4_chanx_right_out[10] ,
    \sb_1__0__4_chanx_right_out[11] ,
    \sb_1__0__4_chanx_right_out[12] ,
    \sb_1__0__4_chanx_right_out[13] ,
    \sb_1__0__4_chanx_right_out[14] ,
    \sb_1__0__4_chanx_right_out[15] ,
    \sb_1__0__4_chanx_right_out[16] ,
    \sb_1__0__4_chanx_right_out[17] ,
    \sb_1__0__4_chanx_right_out[18] ,
    \sb_1__0__4_chanx_right_out[19] }),
    .chany_top_in({\cby_1__1__32_chany_bottom_out[0] ,
    \cby_1__1__32_chany_bottom_out[1] ,
    \cby_1__1__32_chany_bottom_out[2] ,
    \cby_1__1__32_chany_bottom_out[3] ,
    \cby_1__1__32_chany_bottom_out[4] ,
    \cby_1__1__32_chany_bottom_out[5] ,
    \cby_1__1__32_chany_bottom_out[6] ,
    \cby_1__1__32_chany_bottom_out[7] ,
    \cby_1__1__32_chany_bottom_out[8] ,
    \cby_1__1__32_chany_bottom_out[9] ,
    \cby_1__1__32_chany_bottom_out[10] ,
    \cby_1__1__32_chany_bottom_out[11] ,
    \cby_1__1__32_chany_bottom_out[12] ,
    \cby_1__1__32_chany_bottom_out[13] ,
    \cby_1__1__32_chany_bottom_out[14] ,
    \cby_1__1__32_chany_bottom_out[15] ,
    \cby_1__1__32_chany_bottom_out[16] ,
    \cby_1__1__32_chany_bottom_out[17] ,
    \cby_1__1__32_chany_bottom_out[18] ,
    \cby_1__1__32_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__0__4_chany_top_out[0] ,
    \sb_1__0__4_chany_top_out[1] ,
    \sb_1__0__4_chany_top_out[2] ,
    \sb_1__0__4_chany_top_out[3] ,
    \sb_1__0__4_chany_top_out[4] ,
    \sb_1__0__4_chany_top_out[5] ,
    \sb_1__0__4_chany_top_out[6] ,
    \sb_1__0__4_chany_top_out[7] ,
    \sb_1__0__4_chany_top_out[8] ,
    \sb_1__0__4_chany_top_out[9] ,
    \sb_1__0__4_chany_top_out[10] ,
    \sb_1__0__4_chany_top_out[11] ,
    \sb_1__0__4_chany_top_out[12] ,
    \sb_1__0__4_chany_top_out[13] ,
    \sb_1__0__4_chany_top_out[14] ,
    \sb_1__0__4_chany_top_out[15] ,
    \sb_1__0__4_chany_top_out[16] ,
    \sb_1__0__4_chany_top_out[17] ,
    \sb_1__0__4_chany_top_out[18] ,
    \sb_1__0__4_chany_top_out[19] }));
 sb_1__1_ sb_5__1_ (.bottom_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__35_ccff_tail),
    .ccff_tail(sb_1__1__28_ccff_tail),
    .clk_1_E_out(\clk_1_wires[57] ),
    .clk_1_N_in(\clk_2_wires[34] ),
    .clk_1_W_out(\clk_1_wires[58] ),
    .left_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[126] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[57] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[34] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[58] ),
    .right_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__28_chanx_right_out[0] ,
    \cbx_1__1__28_chanx_right_out[1] ,
    \cbx_1__1__28_chanx_right_out[2] ,
    \cbx_1__1__28_chanx_right_out[3] ,
    \cbx_1__1__28_chanx_right_out[4] ,
    \cbx_1__1__28_chanx_right_out[5] ,
    \cbx_1__1__28_chanx_right_out[6] ,
    \cbx_1__1__28_chanx_right_out[7] ,
    \cbx_1__1__28_chanx_right_out[8] ,
    \cbx_1__1__28_chanx_right_out[9] ,
    \cbx_1__1__28_chanx_right_out[10] ,
    \cbx_1__1__28_chanx_right_out[11] ,
    \cbx_1__1__28_chanx_right_out[12] ,
    \cbx_1__1__28_chanx_right_out[13] ,
    \cbx_1__1__28_chanx_right_out[14] ,
    \cbx_1__1__28_chanx_right_out[15] ,
    \cbx_1__1__28_chanx_right_out[16] ,
    \cbx_1__1__28_chanx_right_out[17] ,
    \cbx_1__1__28_chanx_right_out[18] ,
    \cbx_1__1__28_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__28_chanx_left_out[0] ,
    \sb_1__1__28_chanx_left_out[1] ,
    \sb_1__1__28_chanx_left_out[2] ,
    \sb_1__1__28_chanx_left_out[3] ,
    \sb_1__1__28_chanx_left_out[4] ,
    \sb_1__1__28_chanx_left_out[5] ,
    \sb_1__1__28_chanx_left_out[6] ,
    \sb_1__1__28_chanx_left_out[7] ,
    \sb_1__1__28_chanx_left_out[8] ,
    \sb_1__1__28_chanx_left_out[9] ,
    \sb_1__1__28_chanx_left_out[10] ,
    \sb_1__1__28_chanx_left_out[11] ,
    \sb_1__1__28_chanx_left_out[12] ,
    \sb_1__1__28_chanx_left_out[13] ,
    \sb_1__1__28_chanx_left_out[14] ,
    \sb_1__1__28_chanx_left_out[15] ,
    \sb_1__1__28_chanx_left_out[16] ,
    \sb_1__1__28_chanx_left_out[17] ,
    \sb_1__1__28_chanx_left_out[18] ,
    \sb_1__1__28_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__35_chanx_left_out[0] ,
    \cbx_1__1__35_chanx_left_out[1] ,
    \cbx_1__1__35_chanx_left_out[2] ,
    \cbx_1__1__35_chanx_left_out[3] ,
    \cbx_1__1__35_chanx_left_out[4] ,
    \cbx_1__1__35_chanx_left_out[5] ,
    \cbx_1__1__35_chanx_left_out[6] ,
    \cbx_1__1__35_chanx_left_out[7] ,
    \cbx_1__1__35_chanx_left_out[8] ,
    \cbx_1__1__35_chanx_left_out[9] ,
    \cbx_1__1__35_chanx_left_out[10] ,
    \cbx_1__1__35_chanx_left_out[11] ,
    \cbx_1__1__35_chanx_left_out[12] ,
    \cbx_1__1__35_chanx_left_out[13] ,
    \cbx_1__1__35_chanx_left_out[14] ,
    \cbx_1__1__35_chanx_left_out[15] ,
    \cbx_1__1__35_chanx_left_out[16] ,
    \cbx_1__1__35_chanx_left_out[17] ,
    \cbx_1__1__35_chanx_left_out[18] ,
    \cbx_1__1__35_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__28_chanx_right_out[0] ,
    \sb_1__1__28_chanx_right_out[1] ,
    \sb_1__1__28_chanx_right_out[2] ,
    \sb_1__1__28_chanx_right_out[3] ,
    \sb_1__1__28_chanx_right_out[4] ,
    \sb_1__1__28_chanx_right_out[5] ,
    \sb_1__1__28_chanx_right_out[6] ,
    \sb_1__1__28_chanx_right_out[7] ,
    \sb_1__1__28_chanx_right_out[8] ,
    \sb_1__1__28_chanx_right_out[9] ,
    \sb_1__1__28_chanx_right_out[10] ,
    \sb_1__1__28_chanx_right_out[11] ,
    \sb_1__1__28_chanx_right_out[12] ,
    \sb_1__1__28_chanx_right_out[13] ,
    \sb_1__1__28_chanx_right_out[14] ,
    \sb_1__1__28_chanx_right_out[15] ,
    \sb_1__1__28_chanx_right_out[16] ,
    \sb_1__1__28_chanx_right_out[17] ,
    \sb_1__1__28_chanx_right_out[18] ,
    \sb_1__1__28_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__32_chany_top_out[0] ,
    \cby_1__1__32_chany_top_out[1] ,
    \cby_1__1__32_chany_top_out[2] ,
    \cby_1__1__32_chany_top_out[3] ,
    \cby_1__1__32_chany_top_out[4] ,
    \cby_1__1__32_chany_top_out[5] ,
    \cby_1__1__32_chany_top_out[6] ,
    \cby_1__1__32_chany_top_out[7] ,
    \cby_1__1__32_chany_top_out[8] ,
    \cby_1__1__32_chany_top_out[9] ,
    \cby_1__1__32_chany_top_out[10] ,
    \cby_1__1__32_chany_top_out[11] ,
    \cby_1__1__32_chany_top_out[12] ,
    \cby_1__1__32_chany_top_out[13] ,
    \cby_1__1__32_chany_top_out[14] ,
    \cby_1__1__32_chany_top_out[15] ,
    \cby_1__1__32_chany_top_out[16] ,
    \cby_1__1__32_chany_top_out[17] ,
    \cby_1__1__32_chany_top_out[18] ,
    \cby_1__1__32_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__28_chany_bottom_out[0] ,
    \sb_1__1__28_chany_bottom_out[1] ,
    \sb_1__1__28_chany_bottom_out[2] ,
    \sb_1__1__28_chany_bottom_out[3] ,
    \sb_1__1__28_chany_bottom_out[4] ,
    \sb_1__1__28_chany_bottom_out[5] ,
    \sb_1__1__28_chany_bottom_out[6] ,
    \sb_1__1__28_chany_bottom_out[7] ,
    \sb_1__1__28_chany_bottom_out[8] ,
    \sb_1__1__28_chany_bottom_out[9] ,
    \sb_1__1__28_chany_bottom_out[10] ,
    \sb_1__1__28_chany_bottom_out[11] ,
    \sb_1__1__28_chany_bottom_out[12] ,
    \sb_1__1__28_chany_bottom_out[13] ,
    \sb_1__1__28_chany_bottom_out[14] ,
    \sb_1__1__28_chany_bottom_out[15] ,
    \sb_1__1__28_chany_bottom_out[16] ,
    \sb_1__1__28_chany_bottom_out[17] ,
    \sb_1__1__28_chany_bottom_out[18] ,
    \sb_1__1__28_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__33_chany_bottom_out[0] ,
    \cby_1__1__33_chany_bottom_out[1] ,
    \cby_1__1__33_chany_bottom_out[2] ,
    \cby_1__1__33_chany_bottom_out[3] ,
    \cby_1__1__33_chany_bottom_out[4] ,
    \cby_1__1__33_chany_bottom_out[5] ,
    \cby_1__1__33_chany_bottom_out[6] ,
    \cby_1__1__33_chany_bottom_out[7] ,
    \cby_1__1__33_chany_bottom_out[8] ,
    \cby_1__1__33_chany_bottom_out[9] ,
    \cby_1__1__33_chany_bottom_out[10] ,
    \cby_1__1__33_chany_bottom_out[11] ,
    \cby_1__1__33_chany_bottom_out[12] ,
    \cby_1__1__33_chany_bottom_out[13] ,
    \cby_1__1__33_chany_bottom_out[14] ,
    \cby_1__1__33_chany_bottom_out[15] ,
    \cby_1__1__33_chany_bottom_out[16] ,
    \cby_1__1__33_chany_bottom_out[17] ,
    \cby_1__1__33_chany_bottom_out[18] ,
    \cby_1__1__33_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__28_chany_top_out[0] ,
    \sb_1__1__28_chany_top_out[1] ,
    \sb_1__1__28_chany_top_out[2] ,
    \sb_1__1__28_chany_top_out[3] ,
    \sb_1__1__28_chany_top_out[4] ,
    \sb_1__1__28_chany_top_out[5] ,
    \sb_1__1__28_chany_top_out[6] ,
    \sb_1__1__28_chany_top_out[7] ,
    \sb_1__1__28_chany_top_out[8] ,
    \sb_1__1__28_chany_top_out[9] ,
    \sb_1__1__28_chany_top_out[10] ,
    \sb_1__1__28_chany_top_out[11] ,
    \sb_1__1__28_chany_top_out[12] ,
    \sb_1__1__28_chany_top_out[13] ,
    \sb_1__1__28_chany_top_out[14] ,
    \sb_1__1__28_chany_top_out[15] ,
    \sb_1__1__28_chany_top_out[16] ,
    \sb_1__1__28_chany_top_out[17] ,
    \sb_1__1__28_chany_top_out[18] ,
    \sb_1__1__28_chany_top_out[19] }));
 sb_1__1_ sb_5__2_ (.bottom_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__36_ccff_tail),
    .ccff_tail(sb_1__1__29_ccff_tail),
    .clk_2_N_in(\clk_2_wires[30] ),
    .clk_2_N_out(\clk_2_wires[31] ),
    .clk_2_S_out(\clk_2_wires[33] ),
    .left_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[129] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[30] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[31] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[33] ),
    .right_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__29_chanx_right_out[0] ,
    \cbx_1__1__29_chanx_right_out[1] ,
    \cbx_1__1__29_chanx_right_out[2] ,
    \cbx_1__1__29_chanx_right_out[3] ,
    \cbx_1__1__29_chanx_right_out[4] ,
    \cbx_1__1__29_chanx_right_out[5] ,
    \cbx_1__1__29_chanx_right_out[6] ,
    \cbx_1__1__29_chanx_right_out[7] ,
    \cbx_1__1__29_chanx_right_out[8] ,
    \cbx_1__1__29_chanx_right_out[9] ,
    \cbx_1__1__29_chanx_right_out[10] ,
    \cbx_1__1__29_chanx_right_out[11] ,
    \cbx_1__1__29_chanx_right_out[12] ,
    \cbx_1__1__29_chanx_right_out[13] ,
    \cbx_1__1__29_chanx_right_out[14] ,
    \cbx_1__1__29_chanx_right_out[15] ,
    \cbx_1__1__29_chanx_right_out[16] ,
    \cbx_1__1__29_chanx_right_out[17] ,
    \cbx_1__1__29_chanx_right_out[18] ,
    \cbx_1__1__29_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__29_chanx_left_out[0] ,
    \sb_1__1__29_chanx_left_out[1] ,
    \sb_1__1__29_chanx_left_out[2] ,
    \sb_1__1__29_chanx_left_out[3] ,
    \sb_1__1__29_chanx_left_out[4] ,
    \sb_1__1__29_chanx_left_out[5] ,
    \sb_1__1__29_chanx_left_out[6] ,
    \sb_1__1__29_chanx_left_out[7] ,
    \sb_1__1__29_chanx_left_out[8] ,
    \sb_1__1__29_chanx_left_out[9] ,
    \sb_1__1__29_chanx_left_out[10] ,
    \sb_1__1__29_chanx_left_out[11] ,
    \sb_1__1__29_chanx_left_out[12] ,
    \sb_1__1__29_chanx_left_out[13] ,
    \sb_1__1__29_chanx_left_out[14] ,
    \sb_1__1__29_chanx_left_out[15] ,
    \sb_1__1__29_chanx_left_out[16] ,
    \sb_1__1__29_chanx_left_out[17] ,
    \sb_1__1__29_chanx_left_out[18] ,
    \sb_1__1__29_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__36_chanx_left_out[0] ,
    \cbx_1__1__36_chanx_left_out[1] ,
    \cbx_1__1__36_chanx_left_out[2] ,
    \cbx_1__1__36_chanx_left_out[3] ,
    \cbx_1__1__36_chanx_left_out[4] ,
    \cbx_1__1__36_chanx_left_out[5] ,
    \cbx_1__1__36_chanx_left_out[6] ,
    \cbx_1__1__36_chanx_left_out[7] ,
    \cbx_1__1__36_chanx_left_out[8] ,
    \cbx_1__1__36_chanx_left_out[9] ,
    \cbx_1__1__36_chanx_left_out[10] ,
    \cbx_1__1__36_chanx_left_out[11] ,
    \cbx_1__1__36_chanx_left_out[12] ,
    \cbx_1__1__36_chanx_left_out[13] ,
    \cbx_1__1__36_chanx_left_out[14] ,
    \cbx_1__1__36_chanx_left_out[15] ,
    \cbx_1__1__36_chanx_left_out[16] ,
    \cbx_1__1__36_chanx_left_out[17] ,
    \cbx_1__1__36_chanx_left_out[18] ,
    \cbx_1__1__36_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__29_chanx_right_out[0] ,
    \sb_1__1__29_chanx_right_out[1] ,
    \sb_1__1__29_chanx_right_out[2] ,
    \sb_1__1__29_chanx_right_out[3] ,
    \sb_1__1__29_chanx_right_out[4] ,
    \sb_1__1__29_chanx_right_out[5] ,
    \sb_1__1__29_chanx_right_out[6] ,
    \sb_1__1__29_chanx_right_out[7] ,
    \sb_1__1__29_chanx_right_out[8] ,
    \sb_1__1__29_chanx_right_out[9] ,
    \sb_1__1__29_chanx_right_out[10] ,
    \sb_1__1__29_chanx_right_out[11] ,
    \sb_1__1__29_chanx_right_out[12] ,
    \sb_1__1__29_chanx_right_out[13] ,
    \sb_1__1__29_chanx_right_out[14] ,
    \sb_1__1__29_chanx_right_out[15] ,
    \sb_1__1__29_chanx_right_out[16] ,
    \sb_1__1__29_chanx_right_out[17] ,
    \sb_1__1__29_chanx_right_out[18] ,
    \sb_1__1__29_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__33_chany_top_out[0] ,
    \cby_1__1__33_chany_top_out[1] ,
    \cby_1__1__33_chany_top_out[2] ,
    \cby_1__1__33_chany_top_out[3] ,
    \cby_1__1__33_chany_top_out[4] ,
    \cby_1__1__33_chany_top_out[5] ,
    \cby_1__1__33_chany_top_out[6] ,
    \cby_1__1__33_chany_top_out[7] ,
    \cby_1__1__33_chany_top_out[8] ,
    \cby_1__1__33_chany_top_out[9] ,
    \cby_1__1__33_chany_top_out[10] ,
    \cby_1__1__33_chany_top_out[11] ,
    \cby_1__1__33_chany_top_out[12] ,
    \cby_1__1__33_chany_top_out[13] ,
    \cby_1__1__33_chany_top_out[14] ,
    \cby_1__1__33_chany_top_out[15] ,
    \cby_1__1__33_chany_top_out[16] ,
    \cby_1__1__33_chany_top_out[17] ,
    \cby_1__1__33_chany_top_out[18] ,
    \cby_1__1__33_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__29_chany_bottom_out[0] ,
    \sb_1__1__29_chany_bottom_out[1] ,
    \sb_1__1__29_chany_bottom_out[2] ,
    \sb_1__1__29_chany_bottom_out[3] ,
    \sb_1__1__29_chany_bottom_out[4] ,
    \sb_1__1__29_chany_bottom_out[5] ,
    \sb_1__1__29_chany_bottom_out[6] ,
    \sb_1__1__29_chany_bottom_out[7] ,
    \sb_1__1__29_chany_bottom_out[8] ,
    \sb_1__1__29_chany_bottom_out[9] ,
    \sb_1__1__29_chany_bottom_out[10] ,
    \sb_1__1__29_chany_bottom_out[11] ,
    \sb_1__1__29_chany_bottom_out[12] ,
    \sb_1__1__29_chany_bottom_out[13] ,
    \sb_1__1__29_chany_bottom_out[14] ,
    \sb_1__1__29_chany_bottom_out[15] ,
    \sb_1__1__29_chany_bottom_out[16] ,
    \sb_1__1__29_chany_bottom_out[17] ,
    \sb_1__1__29_chany_bottom_out[18] ,
    \sb_1__1__29_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__34_chany_bottom_out[0] ,
    \cby_1__1__34_chany_bottom_out[1] ,
    \cby_1__1__34_chany_bottom_out[2] ,
    \cby_1__1__34_chany_bottom_out[3] ,
    \cby_1__1__34_chany_bottom_out[4] ,
    \cby_1__1__34_chany_bottom_out[5] ,
    \cby_1__1__34_chany_bottom_out[6] ,
    \cby_1__1__34_chany_bottom_out[7] ,
    \cby_1__1__34_chany_bottom_out[8] ,
    \cby_1__1__34_chany_bottom_out[9] ,
    \cby_1__1__34_chany_bottom_out[10] ,
    \cby_1__1__34_chany_bottom_out[11] ,
    \cby_1__1__34_chany_bottom_out[12] ,
    \cby_1__1__34_chany_bottom_out[13] ,
    \cby_1__1__34_chany_bottom_out[14] ,
    \cby_1__1__34_chany_bottom_out[15] ,
    \cby_1__1__34_chany_bottom_out[16] ,
    \cby_1__1__34_chany_bottom_out[17] ,
    \cby_1__1__34_chany_bottom_out[18] ,
    \cby_1__1__34_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__29_chany_top_out[0] ,
    \sb_1__1__29_chany_top_out[1] ,
    \sb_1__1__29_chany_top_out[2] ,
    \sb_1__1__29_chany_top_out[3] ,
    \sb_1__1__29_chany_top_out[4] ,
    \sb_1__1__29_chany_top_out[5] ,
    \sb_1__1__29_chany_top_out[6] ,
    \sb_1__1__29_chany_top_out[7] ,
    \sb_1__1__29_chany_top_out[8] ,
    \sb_1__1__29_chany_top_out[9] ,
    \sb_1__1__29_chany_top_out[10] ,
    \sb_1__1__29_chany_top_out[11] ,
    \sb_1__1__29_chany_top_out[12] ,
    \sb_1__1__29_chany_top_out[13] ,
    \sb_1__1__29_chany_top_out[14] ,
    \sb_1__1__29_chany_top_out[15] ,
    \sb_1__1__29_chany_top_out[16] ,
    \sb_1__1__29_chany_top_out[17] ,
    \sb_1__1__29_chany_top_out[18] ,
    \sb_1__1__29_chany_top_out[19] }));
 sb_1__1_ sb_5__3_ (.bottom_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__37_ccff_tail),
    .ccff_tail(sb_1__1__30_ccff_tail),
    .clk_1_E_out(\clk_1_wires[64] ),
    .clk_1_N_in(\clk_2_wires[32] ),
    .clk_1_W_out(\clk_1_wires[65] ),
    .left_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[132] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[64] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[32] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[65] ),
    .right_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__30_chanx_right_out[0] ,
    \cbx_1__1__30_chanx_right_out[1] ,
    \cbx_1__1__30_chanx_right_out[2] ,
    \cbx_1__1__30_chanx_right_out[3] ,
    \cbx_1__1__30_chanx_right_out[4] ,
    \cbx_1__1__30_chanx_right_out[5] ,
    \cbx_1__1__30_chanx_right_out[6] ,
    \cbx_1__1__30_chanx_right_out[7] ,
    \cbx_1__1__30_chanx_right_out[8] ,
    \cbx_1__1__30_chanx_right_out[9] ,
    \cbx_1__1__30_chanx_right_out[10] ,
    \cbx_1__1__30_chanx_right_out[11] ,
    \cbx_1__1__30_chanx_right_out[12] ,
    \cbx_1__1__30_chanx_right_out[13] ,
    \cbx_1__1__30_chanx_right_out[14] ,
    \cbx_1__1__30_chanx_right_out[15] ,
    \cbx_1__1__30_chanx_right_out[16] ,
    \cbx_1__1__30_chanx_right_out[17] ,
    \cbx_1__1__30_chanx_right_out[18] ,
    \cbx_1__1__30_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__30_chanx_left_out[0] ,
    \sb_1__1__30_chanx_left_out[1] ,
    \sb_1__1__30_chanx_left_out[2] ,
    \sb_1__1__30_chanx_left_out[3] ,
    \sb_1__1__30_chanx_left_out[4] ,
    \sb_1__1__30_chanx_left_out[5] ,
    \sb_1__1__30_chanx_left_out[6] ,
    \sb_1__1__30_chanx_left_out[7] ,
    \sb_1__1__30_chanx_left_out[8] ,
    \sb_1__1__30_chanx_left_out[9] ,
    \sb_1__1__30_chanx_left_out[10] ,
    \sb_1__1__30_chanx_left_out[11] ,
    \sb_1__1__30_chanx_left_out[12] ,
    \sb_1__1__30_chanx_left_out[13] ,
    \sb_1__1__30_chanx_left_out[14] ,
    \sb_1__1__30_chanx_left_out[15] ,
    \sb_1__1__30_chanx_left_out[16] ,
    \sb_1__1__30_chanx_left_out[17] ,
    \sb_1__1__30_chanx_left_out[18] ,
    \sb_1__1__30_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__37_chanx_left_out[0] ,
    \cbx_1__1__37_chanx_left_out[1] ,
    \cbx_1__1__37_chanx_left_out[2] ,
    \cbx_1__1__37_chanx_left_out[3] ,
    \cbx_1__1__37_chanx_left_out[4] ,
    \cbx_1__1__37_chanx_left_out[5] ,
    \cbx_1__1__37_chanx_left_out[6] ,
    \cbx_1__1__37_chanx_left_out[7] ,
    \cbx_1__1__37_chanx_left_out[8] ,
    \cbx_1__1__37_chanx_left_out[9] ,
    \cbx_1__1__37_chanx_left_out[10] ,
    \cbx_1__1__37_chanx_left_out[11] ,
    \cbx_1__1__37_chanx_left_out[12] ,
    \cbx_1__1__37_chanx_left_out[13] ,
    \cbx_1__1__37_chanx_left_out[14] ,
    \cbx_1__1__37_chanx_left_out[15] ,
    \cbx_1__1__37_chanx_left_out[16] ,
    \cbx_1__1__37_chanx_left_out[17] ,
    \cbx_1__1__37_chanx_left_out[18] ,
    \cbx_1__1__37_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__30_chanx_right_out[0] ,
    \sb_1__1__30_chanx_right_out[1] ,
    \sb_1__1__30_chanx_right_out[2] ,
    \sb_1__1__30_chanx_right_out[3] ,
    \sb_1__1__30_chanx_right_out[4] ,
    \sb_1__1__30_chanx_right_out[5] ,
    \sb_1__1__30_chanx_right_out[6] ,
    \sb_1__1__30_chanx_right_out[7] ,
    \sb_1__1__30_chanx_right_out[8] ,
    \sb_1__1__30_chanx_right_out[9] ,
    \sb_1__1__30_chanx_right_out[10] ,
    \sb_1__1__30_chanx_right_out[11] ,
    \sb_1__1__30_chanx_right_out[12] ,
    \sb_1__1__30_chanx_right_out[13] ,
    \sb_1__1__30_chanx_right_out[14] ,
    \sb_1__1__30_chanx_right_out[15] ,
    \sb_1__1__30_chanx_right_out[16] ,
    \sb_1__1__30_chanx_right_out[17] ,
    \sb_1__1__30_chanx_right_out[18] ,
    \sb_1__1__30_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__34_chany_top_out[0] ,
    \cby_1__1__34_chany_top_out[1] ,
    \cby_1__1__34_chany_top_out[2] ,
    \cby_1__1__34_chany_top_out[3] ,
    \cby_1__1__34_chany_top_out[4] ,
    \cby_1__1__34_chany_top_out[5] ,
    \cby_1__1__34_chany_top_out[6] ,
    \cby_1__1__34_chany_top_out[7] ,
    \cby_1__1__34_chany_top_out[8] ,
    \cby_1__1__34_chany_top_out[9] ,
    \cby_1__1__34_chany_top_out[10] ,
    \cby_1__1__34_chany_top_out[11] ,
    \cby_1__1__34_chany_top_out[12] ,
    \cby_1__1__34_chany_top_out[13] ,
    \cby_1__1__34_chany_top_out[14] ,
    \cby_1__1__34_chany_top_out[15] ,
    \cby_1__1__34_chany_top_out[16] ,
    \cby_1__1__34_chany_top_out[17] ,
    \cby_1__1__34_chany_top_out[18] ,
    \cby_1__1__34_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__30_chany_bottom_out[0] ,
    \sb_1__1__30_chany_bottom_out[1] ,
    \sb_1__1__30_chany_bottom_out[2] ,
    \sb_1__1__30_chany_bottom_out[3] ,
    \sb_1__1__30_chany_bottom_out[4] ,
    \sb_1__1__30_chany_bottom_out[5] ,
    \sb_1__1__30_chany_bottom_out[6] ,
    \sb_1__1__30_chany_bottom_out[7] ,
    \sb_1__1__30_chany_bottom_out[8] ,
    \sb_1__1__30_chany_bottom_out[9] ,
    \sb_1__1__30_chany_bottom_out[10] ,
    \sb_1__1__30_chany_bottom_out[11] ,
    \sb_1__1__30_chany_bottom_out[12] ,
    \sb_1__1__30_chany_bottom_out[13] ,
    \sb_1__1__30_chany_bottom_out[14] ,
    \sb_1__1__30_chany_bottom_out[15] ,
    \sb_1__1__30_chany_bottom_out[16] ,
    \sb_1__1__30_chany_bottom_out[17] ,
    \sb_1__1__30_chany_bottom_out[18] ,
    \sb_1__1__30_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__35_chany_bottom_out[0] ,
    \cby_1__1__35_chany_bottom_out[1] ,
    \cby_1__1__35_chany_bottom_out[2] ,
    \cby_1__1__35_chany_bottom_out[3] ,
    \cby_1__1__35_chany_bottom_out[4] ,
    \cby_1__1__35_chany_bottom_out[5] ,
    \cby_1__1__35_chany_bottom_out[6] ,
    \cby_1__1__35_chany_bottom_out[7] ,
    \cby_1__1__35_chany_bottom_out[8] ,
    \cby_1__1__35_chany_bottom_out[9] ,
    \cby_1__1__35_chany_bottom_out[10] ,
    \cby_1__1__35_chany_bottom_out[11] ,
    \cby_1__1__35_chany_bottom_out[12] ,
    \cby_1__1__35_chany_bottom_out[13] ,
    \cby_1__1__35_chany_bottom_out[14] ,
    \cby_1__1__35_chany_bottom_out[15] ,
    \cby_1__1__35_chany_bottom_out[16] ,
    \cby_1__1__35_chany_bottom_out[17] ,
    \cby_1__1__35_chany_bottom_out[18] ,
    \cby_1__1__35_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__30_chany_top_out[0] ,
    \sb_1__1__30_chany_top_out[1] ,
    \sb_1__1__30_chany_top_out[2] ,
    \sb_1__1__30_chany_top_out[3] ,
    \sb_1__1__30_chany_top_out[4] ,
    \sb_1__1__30_chany_top_out[5] ,
    \sb_1__1__30_chany_top_out[6] ,
    \sb_1__1__30_chany_top_out[7] ,
    \sb_1__1__30_chany_top_out[8] ,
    \sb_1__1__30_chany_top_out[9] ,
    \sb_1__1__30_chany_top_out[10] ,
    \sb_1__1__30_chany_top_out[11] ,
    \sb_1__1__30_chany_top_out[12] ,
    \sb_1__1__30_chany_top_out[13] ,
    \sb_1__1__30_chany_top_out[14] ,
    \sb_1__1__30_chany_top_out[15] ,
    \sb_1__1__30_chany_top_out[16] ,
    \sb_1__1__30_chany_top_out[17] ,
    \sb_1__1__30_chany_top_out[18] ,
    \sb_1__1__30_chany_top_out[19] }));
 sb_1__1_ sb_5__4_ (.bottom_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__38_ccff_tail),
    .ccff_tail(sb_1__1__31_ccff_tail),
    .clk_3_E_out(\clk_3_wires[6] ),
    .clk_3_N_in(\clk_3_wires[2] ),
    .left_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[135] ),
    .prog_clk_3_E_out(\prog_clk_3_wires[6] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[2] ),
    .right_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__31_chanx_right_out[0] ,
    \cbx_1__1__31_chanx_right_out[1] ,
    \cbx_1__1__31_chanx_right_out[2] ,
    \cbx_1__1__31_chanx_right_out[3] ,
    \cbx_1__1__31_chanx_right_out[4] ,
    \cbx_1__1__31_chanx_right_out[5] ,
    \cbx_1__1__31_chanx_right_out[6] ,
    \cbx_1__1__31_chanx_right_out[7] ,
    \cbx_1__1__31_chanx_right_out[8] ,
    \cbx_1__1__31_chanx_right_out[9] ,
    \cbx_1__1__31_chanx_right_out[10] ,
    \cbx_1__1__31_chanx_right_out[11] ,
    \cbx_1__1__31_chanx_right_out[12] ,
    \cbx_1__1__31_chanx_right_out[13] ,
    \cbx_1__1__31_chanx_right_out[14] ,
    \cbx_1__1__31_chanx_right_out[15] ,
    \cbx_1__1__31_chanx_right_out[16] ,
    \cbx_1__1__31_chanx_right_out[17] ,
    \cbx_1__1__31_chanx_right_out[18] ,
    \cbx_1__1__31_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__31_chanx_left_out[0] ,
    \sb_1__1__31_chanx_left_out[1] ,
    \sb_1__1__31_chanx_left_out[2] ,
    \sb_1__1__31_chanx_left_out[3] ,
    \sb_1__1__31_chanx_left_out[4] ,
    \sb_1__1__31_chanx_left_out[5] ,
    \sb_1__1__31_chanx_left_out[6] ,
    \sb_1__1__31_chanx_left_out[7] ,
    \sb_1__1__31_chanx_left_out[8] ,
    \sb_1__1__31_chanx_left_out[9] ,
    \sb_1__1__31_chanx_left_out[10] ,
    \sb_1__1__31_chanx_left_out[11] ,
    \sb_1__1__31_chanx_left_out[12] ,
    \sb_1__1__31_chanx_left_out[13] ,
    \sb_1__1__31_chanx_left_out[14] ,
    \sb_1__1__31_chanx_left_out[15] ,
    \sb_1__1__31_chanx_left_out[16] ,
    \sb_1__1__31_chanx_left_out[17] ,
    \sb_1__1__31_chanx_left_out[18] ,
    \sb_1__1__31_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__38_chanx_left_out[0] ,
    \cbx_1__1__38_chanx_left_out[1] ,
    \cbx_1__1__38_chanx_left_out[2] ,
    \cbx_1__1__38_chanx_left_out[3] ,
    \cbx_1__1__38_chanx_left_out[4] ,
    \cbx_1__1__38_chanx_left_out[5] ,
    \cbx_1__1__38_chanx_left_out[6] ,
    \cbx_1__1__38_chanx_left_out[7] ,
    \cbx_1__1__38_chanx_left_out[8] ,
    \cbx_1__1__38_chanx_left_out[9] ,
    \cbx_1__1__38_chanx_left_out[10] ,
    \cbx_1__1__38_chanx_left_out[11] ,
    \cbx_1__1__38_chanx_left_out[12] ,
    \cbx_1__1__38_chanx_left_out[13] ,
    \cbx_1__1__38_chanx_left_out[14] ,
    \cbx_1__1__38_chanx_left_out[15] ,
    \cbx_1__1__38_chanx_left_out[16] ,
    \cbx_1__1__38_chanx_left_out[17] ,
    \cbx_1__1__38_chanx_left_out[18] ,
    \cbx_1__1__38_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__31_chanx_right_out[0] ,
    \sb_1__1__31_chanx_right_out[1] ,
    \sb_1__1__31_chanx_right_out[2] ,
    \sb_1__1__31_chanx_right_out[3] ,
    \sb_1__1__31_chanx_right_out[4] ,
    \sb_1__1__31_chanx_right_out[5] ,
    \sb_1__1__31_chanx_right_out[6] ,
    \sb_1__1__31_chanx_right_out[7] ,
    \sb_1__1__31_chanx_right_out[8] ,
    \sb_1__1__31_chanx_right_out[9] ,
    \sb_1__1__31_chanx_right_out[10] ,
    \sb_1__1__31_chanx_right_out[11] ,
    \sb_1__1__31_chanx_right_out[12] ,
    \sb_1__1__31_chanx_right_out[13] ,
    \sb_1__1__31_chanx_right_out[14] ,
    \sb_1__1__31_chanx_right_out[15] ,
    \sb_1__1__31_chanx_right_out[16] ,
    \sb_1__1__31_chanx_right_out[17] ,
    \sb_1__1__31_chanx_right_out[18] ,
    \sb_1__1__31_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__35_chany_top_out[0] ,
    \cby_1__1__35_chany_top_out[1] ,
    \cby_1__1__35_chany_top_out[2] ,
    \cby_1__1__35_chany_top_out[3] ,
    \cby_1__1__35_chany_top_out[4] ,
    \cby_1__1__35_chany_top_out[5] ,
    \cby_1__1__35_chany_top_out[6] ,
    \cby_1__1__35_chany_top_out[7] ,
    \cby_1__1__35_chany_top_out[8] ,
    \cby_1__1__35_chany_top_out[9] ,
    \cby_1__1__35_chany_top_out[10] ,
    \cby_1__1__35_chany_top_out[11] ,
    \cby_1__1__35_chany_top_out[12] ,
    \cby_1__1__35_chany_top_out[13] ,
    \cby_1__1__35_chany_top_out[14] ,
    \cby_1__1__35_chany_top_out[15] ,
    \cby_1__1__35_chany_top_out[16] ,
    \cby_1__1__35_chany_top_out[17] ,
    \cby_1__1__35_chany_top_out[18] ,
    \cby_1__1__35_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__31_chany_bottom_out[0] ,
    \sb_1__1__31_chany_bottom_out[1] ,
    \sb_1__1__31_chany_bottom_out[2] ,
    \sb_1__1__31_chany_bottom_out[3] ,
    \sb_1__1__31_chany_bottom_out[4] ,
    \sb_1__1__31_chany_bottom_out[5] ,
    \sb_1__1__31_chany_bottom_out[6] ,
    \sb_1__1__31_chany_bottom_out[7] ,
    \sb_1__1__31_chany_bottom_out[8] ,
    \sb_1__1__31_chany_bottom_out[9] ,
    \sb_1__1__31_chany_bottom_out[10] ,
    \sb_1__1__31_chany_bottom_out[11] ,
    \sb_1__1__31_chany_bottom_out[12] ,
    \sb_1__1__31_chany_bottom_out[13] ,
    \sb_1__1__31_chany_bottom_out[14] ,
    \sb_1__1__31_chany_bottom_out[15] ,
    \sb_1__1__31_chany_bottom_out[16] ,
    \sb_1__1__31_chany_bottom_out[17] ,
    \sb_1__1__31_chany_bottom_out[18] ,
    \sb_1__1__31_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__36_chany_bottom_out[0] ,
    \cby_1__1__36_chany_bottom_out[1] ,
    \cby_1__1__36_chany_bottom_out[2] ,
    \cby_1__1__36_chany_bottom_out[3] ,
    \cby_1__1__36_chany_bottom_out[4] ,
    \cby_1__1__36_chany_bottom_out[5] ,
    \cby_1__1__36_chany_bottom_out[6] ,
    \cby_1__1__36_chany_bottom_out[7] ,
    \cby_1__1__36_chany_bottom_out[8] ,
    \cby_1__1__36_chany_bottom_out[9] ,
    \cby_1__1__36_chany_bottom_out[10] ,
    \cby_1__1__36_chany_bottom_out[11] ,
    \cby_1__1__36_chany_bottom_out[12] ,
    \cby_1__1__36_chany_bottom_out[13] ,
    \cby_1__1__36_chany_bottom_out[14] ,
    \cby_1__1__36_chany_bottom_out[15] ,
    \cby_1__1__36_chany_bottom_out[16] ,
    \cby_1__1__36_chany_bottom_out[17] ,
    \cby_1__1__36_chany_bottom_out[18] ,
    \cby_1__1__36_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__31_chany_top_out[0] ,
    \sb_1__1__31_chany_top_out[1] ,
    \sb_1__1__31_chany_top_out[2] ,
    \sb_1__1__31_chany_top_out[3] ,
    \sb_1__1__31_chany_top_out[4] ,
    \sb_1__1__31_chany_top_out[5] ,
    \sb_1__1__31_chany_top_out[6] ,
    \sb_1__1__31_chany_top_out[7] ,
    \sb_1__1__31_chany_top_out[8] ,
    \sb_1__1__31_chany_top_out[9] ,
    \sb_1__1__31_chany_top_out[10] ,
    \sb_1__1__31_chany_top_out[11] ,
    \sb_1__1__31_chany_top_out[12] ,
    \sb_1__1__31_chany_top_out[13] ,
    \sb_1__1__31_chany_top_out[14] ,
    \sb_1__1__31_chany_top_out[15] ,
    \sb_1__1__31_chany_top_out[16] ,
    \sb_1__1__31_chany_top_out[17] ,
    \sb_1__1__31_chany_top_out[18] ,
    \sb_1__1__31_chany_top_out[19] }));
 sb_1__1_ sb_5__5_ (.bottom_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__39_ccff_tail),
    .ccff_tail(sb_1__1__32_ccff_tail),
    .clk_1_E_out(\clk_1_wires[71] ),
    .clk_1_N_in(\clk_2_wires[47] ),
    .clk_1_W_out(\clk_1_wires[72] ),
    .left_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[138] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[71] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[47] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[72] ),
    .right_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__32_chanx_right_out[0] ,
    \cbx_1__1__32_chanx_right_out[1] ,
    \cbx_1__1__32_chanx_right_out[2] ,
    \cbx_1__1__32_chanx_right_out[3] ,
    \cbx_1__1__32_chanx_right_out[4] ,
    \cbx_1__1__32_chanx_right_out[5] ,
    \cbx_1__1__32_chanx_right_out[6] ,
    \cbx_1__1__32_chanx_right_out[7] ,
    \cbx_1__1__32_chanx_right_out[8] ,
    \cbx_1__1__32_chanx_right_out[9] ,
    \cbx_1__1__32_chanx_right_out[10] ,
    \cbx_1__1__32_chanx_right_out[11] ,
    \cbx_1__1__32_chanx_right_out[12] ,
    \cbx_1__1__32_chanx_right_out[13] ,
    \cbx_1__1__32_chanx_right_out[14] ,
    \cbx_1__1__32_chanx_right_out[15] ,
    \cbx_1__1__32_chanx_right_out[16] ,
    \cbx_1__1__32_chanx_right_out[17] ,
    \cbx_1__1__32_chanx_right_out[18] ,
    \cbx_1__1__32_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__32_chanx_left_out[0] ,
    \sb_1__1__32_chanx_left_out[1] ,
    \sb_1__1__32_chanx_left_out[2] ,
    \sb_1__1__32_chanx_left_out[3] ,
    \sb_1__1__32_chanx_left_out[4] ,
    \sb_1__1__32_chanx_left_out[5] ,
    \sb_1__1__32_chanx_left_out[6] ,
    \sb_1__1__32_chanx_left_out[7] ,
    \sb_1__1__32_chanx_left_out[8] ,
    \sb_1__1__32_chanx_left_out[9] ,
    \sb_1__1__32_chanx_left_out[10] ,
    \sb_1__1__32_chanx_left_out[11] ,
    \sb_1__1__32_chanx_left_out[12] ,
    \sb_1__1__32_chanx_left_out[13] ,
    \sb_1__1__32_chanx_left_out[14] ,
    \sb_1__1__32_chanx_left_out[15] ,
    \sb_1__1__32_chanx_left_out[16] ,
    \sb_1__1__32_chanx_left_out[17] ,
    \sb_1__1__32_chanx_left_out[18] ,
    \sb_1__1__32_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__39_chanx_left_out[0] ,
    \cbx_1__1__39_chanx_left_out[1] ,
    \cbx_1__1__39_chanx_left_out[2] ,
    \cbx_1__1__39_chanx_left_out[3] ,
    \cbx_1__1__39_chanx_left_out[4] ,
    \cbx_1__1__39_chanx_left_out[5] ,
    \cbx_1__1__39_chanx_left_out[6] ,
    \cbx_1__1__39_chanx_left_out[7] ,
    \cbx_1__1__39_chanx_left_out[8] ,
    \cbx_1__1__39_chanx_left_out[9] ,
    \cbx_1__1__39_chanx_left_out[10] ,
    \cbx_1__1__39_chanx_left_out[11] ,
    \cbx_1__1__39_chanx_left_out[12] ,
    \cbx_1__1__39_chanx_left_out[13] ,
    \cbx_1__1__39_chanx_left_out[14] ,
    \cbx_1__1__39_chanx_left_out[15] ,
    \cbx_1__1__39_chanx_left_out[16] ,
    \cbx_1__1__39_chanx_left_out[17] ,
    \cbx_1__1__39_chanx_left_out[18] ,
    \cbx_1__1__39_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__32_chanx_right_out[0] ,
    \sb_1__1__32_chanx_right_out[1] ,
    \sb_1__1__32_chanx_right_out[2] ,
    \sb_1__1__32_chanx_right_out[3] ,
    \sb_1__1__32_chanx_right_out[4] ,
    \sb_1__1__32_chanx_right_out[5] ,
    \sb_1__1__32_chanx_right_out[6] ,
    \sb_1__1__32_chanx_right_out[7] ,
    \sb_1__1__32_chanx_right_out[8] ,
    \sb_1__1__32_chanx_right_out[9] ,
    \sb_1__1__32_chanx_right_out[10] ,
    \sb_1__1__32_chanx_right_out[11] ,
    \sb_1__1__32_chanx_right_out[12] ,
    \sb_1__1__32_chanx_right_out[13] ,
    \sb_1__1__32_chanx_right_out[14] ,
    \sb_1__1__32_chanx_right_out[15] ,
    \sb_1__1__32_chanx_right_out[16] ,
    \sb_1__1__32_chanx_right_out[17] ,
    \sb_1__1__32_chanx_right_out[18] ,
    \sb_1__1__32_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__36_chany_top_out[0] ,
    \cby_1__1__36_chany_top_out[1] ,
    \cby_1__1__36_chany_top_out[2] ,
    \cby_1__1__36_chany_top_out[3] ,
    \cby_1__1__36_chany_top_out[4] ,
    \cby_1__1__36_chany_top_out[5] ,
    \cby_1__1__36_chany_top_out[6] ,
    \cby_1__1__36_chany_top_out[7] ,
    \cby_1__1__36_chany_top_out[8] ,
    \cby_1__1__36_chany_top_out[9] ,
    \cby_1__1__36_chany_top_out[10] ,
    \cby_1__1__36_chany_top_out[11] ,
    \cby_1__1__36_chany_top_out[12] ,
    \cby_1__1__36_chany_top_out[13] ,
    \cby_1__1__36_chany_top_out[14] ,
    \cby_1__1__36_chany_top_out[15] ,
    \cby_1__1__36_chany_top_out[16] ,
    \cby_1__1__36_chany_top_out[17] ,
    \cby_1__1__36_chany_top_out[18] ,
    \cby_1__1__36_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__32_chany_bottom_out[0] ,
    \sb_1__1__32_chany_bottom_out[1] ,
    \sb_1__1__32_chany_bottom_out[2] ,
    \sb_1__1__32_chany_bottom_out[3] ,
    \sb_1__1__32_chany_bottom_out[4] ,
    \sb_1__1__32_chany_bottom_out[5] ,
    \sb_1__1__32_chany_bottom_out[6] ,
    \sb_1__1__32_chany_bottom_out[7] ,
    \sb_1__1__32_chany_bottom_out[8] ,
    \sb_1__1__32_chany_bottom_out[9] ,
    \sb_1__1__32_chany_bottom_out[10] ,
    \sb_1__1__32_chany_bottom_out[11] ,
    \sb_1__1__32_chany_bottom_out[12] ,
    \sb_1__1__32_chany_bottom_out[13] ,
    \sb_1__1__32_chany_bottom_out[14] ,
    \sb_1__1__32_chany_bottom_out[15] ,
    \sb_1__1__32_chany_bottom_out[16] ,
    \sb_1__1__32_chany_bottom_out[17] ,
    \sb_1__1__32_chany_bottom_out[18] ,
    \sb_1__1__32_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__37_chany_bottom_out[0] ,
    \cby_1__1__37_chany_bottom_out[1] ,
    \cby_1__1__37_chany_bottom_out[2] ,
    \cby_1__1__37_chany_bottom_out[3] ,
    \cby_1__1__37_chany_bottom_out[4] ,
    \cby_1__1__37_chany_bottom_out[5] ,
    \cby_1__1__37_chany_bottom_out[6] ,
    \cby_1__1__37_chany_bottom_out[7] ,
    \cby_1__1__37_chany_bottom_out[8] ,
    \cby_1__1__37_chany_bottom_out[9] ,
    \cby_1__1__37_chany_bottom_out[10] ,
    \cby_1__1__37_chany_bottom_out[11] ,
    \cby_1__1__37_chany_bottom_out[12] ,
    \cby_1__1__37_chany_bottom_out[13] ,
    \cby_1__1__37_chany_bottom_out[14] ,
    \cby_1__1__37_chany_bottom_out[15] ,
    \cby_1__1__37_chany_bottom_out[16] ,
    \cby_1__1__37_chany_bottom_out[17] ,
    \cby_1__1__37_chany_bottom_out[18] ,
    \cby_1__1__37_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__32_chany_top_out[0] ,
    \sb_1__1__32_chany_top_out[1] ,
    \sb_1__1__32_chany_top_out[2] ,
    \sb_1__1__32_chany_top_out[3] ,
    \sb_1__1__32_chany_top_out[4] ,
    \sb_1__1__32_chany_top_out[5] ,
    \sb_1__1__32_chany_top_out[6] ,
    \sb_1__1__32_chany_top_out[7] ,
    \sb_1__1__32_chany_top_out[8] ,
    \sb_1__1__32_chany_top_out[9] ,
    \sb_1__1__32_chany_top_out[10] ,
    \sb_1__1__32_chany_top_out[11] ,
    \sb_1__1__32_chany_top_out[12] ,
    \sb_1__1__32_chany_top_out[13] ,
    \sb_1__1__32_chany_top_out[14] ,
    \sb_1__1__32_chany_top_out[15] ,
    \sb_1__1__32_chany_top_out[16] ,
    \sb_1__1__32_chany_top_out[17] ,
    \sb_1__1__32_chany_top_out[18] ,
    \sb_1__1__32_chany_top_out[19] }));
 sb_1__1_ sb_5__6_ (.bottom_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__40_ccff_tail),
    .ccff_tail(sb_1__1__33_ccff_tail),
    .clk_2_N_in(\clk_2_wires[43] ),
    .clk_2_N_out(\clk_2_wires[44] ),
    .clk_2_S_out(\clk_2_wires[46] ),
    .left_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[141] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[43] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[44] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[46] ),
    .right_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__33_chanx_right_out[0] ,
    \cbx_1__1__33_chanx_right_out[1] ,
    \cbx_1__1__33_chanx_right_out[2] ,
    \cbx_1__1__33_chanx_right_out[3] ,
    \cbx_1__1__33_chanx_right_out[4] ,
    \cbx_1__1__33_chanx_right_out[5] ,
    \cbx_1__1__33_chanx_right_out[6] ,
    \cbx_1__1__33_chanx_right_out[7] ,
    \cbx_1__1__33_chanx_right_out[8] ,
    \cbx_1__1__33_chanx_right_out[9] ,
    \cbx_1__1__33_chanx_right_out[10] ,
    \cbx_1__1__33_chanx_right_out[11] ,
    \cbx_1__1__33_chanx_right_out[12] ,
    \cbx_1__1__33_chanx_right_out[13] ,
    \cbx_1__1__33_chanx_right_out[14] ,
    \cbx_1__1__33_chanx_right_out[15] ,
    \cbx_1__1__33_chanx_right_out[16] ,
    \cbx_1__1__33_chanx_right_out[17] ,
    \cbx_1__1__33_chanx_right_out[18] ,
    \cbx_1__1__33_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__33_chanx_left_out[0] ,
    \sb_1__1__33_chanx_left_out[1] ,
    \sb_1__1__33_chanx_left_out[2] ,
    \sb_1__1__33_chanx_left_out[3] ,
    \sb_1__1__33_chanx_left_out[4] ,
    \sb_1__1__33_chanx_left_out[5] ,
    \sb_1__1__33_chanx_left_out[6] ,
    \sb_1__1__33_chanx_left_out[7] ,
    \sb_1__1__33_chanx_left_out[8] ,
    \sb_1__1__33_chanx_left_out[9] ,
    \sb_1__1__33_chanx_left_out[10] ,
    \sb_1__1__33_chanx_left_out[11] ,
    \sb_1__1__33_chanx_left_out[12] ,
    \sb_1__1__33_chanx_left_out[13] ,
    \sb_1__1__33_chanx_left_out[14] ,
    \sb_1__1__33_chanx_left_out[15] ,
    \sb_1__1__33_chanx_left_out[16] ,
    \sb_1__1__33_chanx_left_out[17] ,
    \sb_1__1__33_chanx_left_out[18] ,
    \sb_1__1__33_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__40_chanx_left_out[0] ,
    \cbx_1__1__40_chanx_left_out[1] ,
    \cbx_1__1__40_chanx_left_out[2] ,
    \cbx_1__1__40_chanx_left_out[3] ,
    \cbx_1__1__40_chanx_left_out[4] ,
    \cbx_1__1__40_chanx_left_out[5] ,
    \cbx_1__1__40_chanx_left_out[6] ,
    \cbx_1__1__40_chanx_left_out[7] ,
    \cbx_1__1__40_chanx_left_out[8] ,
    \cbx_1__1__40_chanx_left_out[9] ,
    \cbx_1__1__40_chanx_left_out[10] ,
    \cbx_1__1__40_chanx_left_out[11] ,
    \cbx_1__1__40_chanx_left_out[12] ,
    \cbx_1__1__40_chanx_left_out[13] ,
    \cbx_1__1__40_chanx_left_out[14] ,
    \cbx_1__1__40_chanx_left_out[15] ,
    \cbx_1__1__40_chanx_left_out[16] ,
    \cbx_1__1__40_chanx_left_out[17] ,
    \cbx_1__1__40_chanx_left_out[18] ,
    \cbx_1__1__40_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__33_chanx_right_out[0] ,
    \sb_1__1__33_chanx_right_out[1] ,
    \sb_1__1__33_chanx_right_out[2] ,
    \sb_1__1__33_chanx_right_out[3] ,
    \sb_1__1__33_chanx_right_out[4] ,
    \sb_1__1__33_chanx_right_out[5] ,
    \sb_1__1__33_chanx_right_out[6] ,
    \sb_1__1__33_chanx_right_out[7] ,
    \sb_1__1__33_chanx_right_out[8] ,
    \sb_1__1__33_chanx_right_out[9] ,
    \sb_1__1__33_chanx_right_out[10] ,
    \sb_1__1__33_chanx_right_out[11] ,
    \sb_1__1__33_chanx_right_out[12] ,
    \sb_1__1__33_chanx_right_out[13] ,
    \sb_1__1__33_chanx_right_out[14] ,
    \sb_1__1__33_chanx_right_out[15] ,
    \sb_1__1__33_chanx_right_out[16] ,
    \sb_1__1__33_chanx_right_out[17] ,
    \sb_1__1__33_chanx_right_out[18] ,
    \sb_1__1__33_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__37_chany_top_out[0] ,
    \cby_1__1__37_chany_top_out[1] ,
    \cby_1__1__37_chany_top_out[2] ,
    \cby_1__1__37_chany_top_out[3] ,
    \cby_1__1__37_chany_top_out[4] ,
    \cby_1__1__37_chany_top_out[5] ,
    \cby_1__1__37_chany_top_out[6] ,
    \cby_1__1__37_chany_top_out[7] ,
    \cby_1__1__37_chany_top_out[8] ,
    \cby_1__1__37_chany_top_out[9] ,
    \cby_1__1__37_chany_top_out[10] ,
    \cby_1__1__37_chany_top_out[11] ,
    \cby_1__1__37_chany_top_out[12] ,
    \cby_1__1__37_chany_top_out[13] ,
    \cby_1__1__37_chany_top_out[14] ,
    \cby_1__1__37_chany_top_out[15] ,
    \cby_1__1__37_chany_top_out[16] ,
    \cby_1__1__37_chany_top_out[17] ,
    \cby_1__1__37_chany_top_out[18] ,
    \cby_1__1__37_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__33_chany_bottom_out[0] ,
    \sb_1__1__33_chany_bottom_out[1] ,
    \sb_1__1__33_chany_bottom_out[2] ,
    \sb_1__1__33_chany_bottom_out[3] ,
    \sb_1__1__33_chany_bottom_out[4] ,
    \sb_1__1__33_chany_bottom_out[5] ,
    \sb_1__1__33_chany_bottom_out[6] ,
    \sb_1__1__33_chany_bottom_out[7] ,
    \sb_1__1__33_chany_bottom_out[8] ,
    \sb_1__1__33_chany_bottom_out[9] ,
    \sb_1__1__33_chany_bottom_out[10] ,
    \sb_1__1__33_chany_bottom_out[11] ,
    \sb_1__1__33_chany_bottom_out[12] ,
    \sb_1__1__33_chany_bottom_out[13] ,
    \sb_1__1__33_chany_bottom_out[14] ,
    \sb_1__1__33_chany_bottom_out[15] ,
    \sb_1__1__33_chany_bottom_out[16] ,
    \sb_1__1__33_chany_bottom_out[17] ,
    \sb_1__1__33_chany_bottom_out[18] ,
    \sb_1__1__33_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__38_chany_bottom_out[0] ,
    \cby_1__1__38_chany_bottom_out[1] ,
    \cby_1__1__38_chany_bottom_out[2] ,
    \cby_1__1__38_chany_bottom_out[3] ,
    \cby_1__1__38_chany_bottom_out[4] ,
    \cby_1__1__38_chany_bottom_out[5] ,
    \cby_1__1__38_chany_bottom_out[6] ,
    \cby_1__1__38_chany_bottom_out[7] ,
    \cby_1__1__38_chany_bottom_out[8] ,
    \cby_1__1__38_chany_bottom_out[9] ,
    \cby_1__1__38_chany_bottom_out[10] ,
    \cby_1__1__38_chany_bottom_out[11] ,
    \cby_1__1__38_chany_bottom_out[12] ,
    \cby_1__1__38_chany_bottom_out[13] ,
    \cby_1__1__38_chany_bottom_out[14] ,
    \cby_1__1__38_chany_bottom_out[15] ,
    \cby_1__1__38_chany_bottom_out[16] ,
    \cby_1__1__38_chany_bottom_out[17] ,
    \cby_1__1__38_chany_bottom_out[18] ,
    \cby_1__1__38_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__33_chany_top_out[0] ,
    \sb_1__1__33_chany_top_out[1] ,
    \sb_1__1__33_chany_top_out[2] ,
    \sb_1__1__33_chany_top_out[3] ,
    \sb_1__1__33_chany_top_out[4] ,
    \sb_1__1__33_chany_top_out[5] ,
    \sb_1__1__33_chany_top_out[6] ,
    \sb_1__1__33_chany_top_out[7] ,
    \sb_1__1__33_chany_top_out[8] ,
    \sb_1__1__33_chany_top_out[9] ,
    \sb_1__1__33_chany_top_out[10] ,
    \sb_1__1__33_chany_top_out[11] ,
    \sb_1__1__33_chany_top_out[12] ,
    \sb_1__1__33_chany_top_out[13] ,
    \sb_1__1__33_chany_top_out[14] ,
    \sb_1__1__33_chany_top_out[15] ,
    \sb_1__1__33_chany_top_out[16] ,
    \sb_1__1__33_chany_top_out[17] ,
    \sb_1__1__33_chany_top_out[18] ,
    \sb_1__1__33_chany_top_out[19] }));
 sb_1__1_ sb_5__7_ (.bottom_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__41_ccff_tail),
    .ccff_tail(sb_1__1__34_ccff_tail),
    .clk_1_E_out(\clk_1_wires[78] ),
    .clk_1_N_in(\clk_2_wires[45] ),
    .clk_1_W_out(\clk_1_wires[79] ),
    .left_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[144] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[78] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[45] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[79] ),
    .right_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__34_chanx_right_out[0] ,
    \cbx_1__1__34_chanx_right_out[1] ,
    \cbx_1__1__34_chanx_right_out[2] ,
    \cbx_1__1__34_chanx_right_out[3] ,
    \cbx_1__1__34_chanx_right_out[4] ,
    \cbx_1__1__34_chanx_right_out[5] ,
    \cbx_1__1__34_chanx_right_out[6] ,
    \cbx_1__1__34_chanx_right_out[7] ,
    \cbx_1__1__34_chanx_right_out[8] ,
    \cbx_1__1__34_chanx_right_out[9] ,
    \cbx_1__1__34_chanx_right_out[10] ,
    \cbx_1__1__34_chanx_right_out[11] ,
    \cbx_1__1__34_chanx_right_out[12] ,
    \cbx_1__1__34_chanx_right_out[13] ,
    \cbx_1__1__34_chanx_right_out[14] ,
    \cbx_1__1__34_chanx_right_out[15] ,
    \cbx_1__1__34_chanx_right_out[16] ,
    \cbx_1__1__34_chanx_right_out[17] ,
    \cbx_1__1__34_chanx_right_out[18] ,
    \cbx_1__1__34_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__34_chanx_left_out[0] ,
    \sb_1__1__34_chanx_left_out[1] ,
    \sb_1__1__34_chanx_left_out[2] ,
    \sb_1__1__34_chanx_left_out[3] ,
    \sb_1__1__34_chanx_left_out[4] ,
    \sb_1__1__34_chanx_left_out[5] ,
    \sb_1__1__34_chanx_left_out[6] ,
    \sb_1__1__34_chanx_left_out[7] ,
    \sb_1__1__34_chanx_left_out[8] ,
    \sb_1__1__34_chanx_left_out[9] ,
    \sb_1__1__34_chanx_left_out[10] ,
    \sb_1__1__34_chanx_left_out[11] ,
    \sb_1__1__34_chanx_left_out[12] ,
    \sb_1__1__34_chanx_left_out[13] ,
    \sb_1__1__34_chanx_left_out[14] ,
    \sb_1__1__34_chanx_left_out[15] ,
    \sb_1__1__34_chanx_left_out[16] ,
    \sb_1__1__34_chanx_left_out[17] ,
    \sb_1__1__34_chanx_left_out[18] ,
    \sb_1__1__34_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__41_chanx_left_out[0] ,
    \cbx_1__1__41_chanx_left_out[1] ,
    \cbx_1__1__41_chanx_left_out[2] ,
    \cbx_1__1__41_chanx_left_out[3] ,
    \cbx_1__1__41_chanx_left_out[4] ,
    \cbx_1__1__41_chanx_left_out[5] ,
    \cbx_1__1__41_chanx_left_out[6] ,
    \cbx_1__1__41_chanx_left_out[7] ,
    \cbx_1__1__41_chanx_left_out[8] ,
    \cbx_1__1__41_chanx_left_out[9] ,
    \cbx_1__1__41_chanx_left_out[10] ,
    \cbx_1__1__41_chanx_left_out[11] ,
    \cbx_1__1__41_chanx_left_out[12] ,
    \cbx_1__1__41_chanx_left_out[13] ,
    \cbx_1__1__41_chanx_left_out[14] ,
    \cbx_1__1__41_chanx_left_out[15] ,
    \cbx_1__1__41_chanx_left_out[16] ,
    \cbx_1__1__41_chanx_left_out[17] ,
    \cbx_1__1__41_chanx_left_out[18] ,
    \cbx_1__1__41_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__34_chanx_right_out[0] ,
    \sb_1__1__34_chanx_right_out[1] ,
    \sb_1__1__34_chanx_right_out[2] ,
    \sb_1__1__34_chanx_right_out[3] ,
    \sb_1__1__34_chanx_right_out[4] ,
    \sb_1__1__34_chanx_right_out[5] ,
    \sb_1__1__34_chanx_right_out[6] ,
    \sb_1__1__34_chanx_right_out[7] ,
    \sb_1__1__34_chanx_right_out[8] ,
    \sb_1__1__34_chanx_right_out[9] ,
    \sb_1__1__34_chanx_right_out[10] ,
    \sb_1__1__34_chanx_right_out[11] ,
    \sb_1__1__34_chanx_right_out[12] ,
    \sb_1__1__34_chanx_right_out[13] ,
    \sb_1__1__34_chanx_right_out[14] ,
    \sb_1__1__34_chanx_right_out[15] ,
    \sb_1__1__34_chanx_right_out[16] ,
    \sb_1__1__34_chanx_right_out[17] ,
    \sb_1__1__34_chanx_right_out[18] ,
    \sb_1__1__34_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__38_chany_top_out[0] ,
    \cby_1__1__38_chany_top_out[1] ,
    \cby_1__1__38_chany_top_out[2] ,
    \cby_1__1__38_chany_top_out[3] ,
    \cby_1__1__38_chany_top_out[4] ,
    \cby_1__1__38_chany_top_out[5] ,
    \cby_1__1__38_chany_top_out[6] ,
    \cby_1__1__38_chany_top_out[7] ,
    \cby_1__1__38_chany_top_out[8] ,
    \cby_1__1__38_chany_top_out[9] ,
    \cby_1__1__38_chany_top_out[10] ,
    \cby_1__1__38_chany_top_out[11] ,
    \cby_1__1__38_chany_top_out[12] ,
    \cby_1__1__38_chany_top_out[13] ,
    \cby_1__1__38_chany_top_out[14] ,
    \cby_1__1__38_chany_top_out[15] ,
    \cby_1__1__38_chany_top_out[16] ,
    \cby_1__1__38_chany_top_out[17] ,
    \cby_1__1__38_chany_top_out[18] ,
    \cby_1__1__38_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__34_chany_bottom_out[0] ,
    \sb_1__1__34_chany_bottom_out[1] ,
    \sb_1__1__34_chany_bottom_out[2] ,
    \sb_1__1__34_chany_bottom_out[3] ,
    \sb_1__1__34_chany_bottom_out[4] ,
    \sb_1__1__34_chany_bottom_out[5] ,
    \sb_1__1__34_chany_bottom_out[6] ,
    \sb_1__1__34_chany_bottom_out[7] ,
    \sb_1__1__34_chany_bottom_out[8] ,
    \sb_1__1__34_chany_bottom_out[9] ,
    \sb_1__1__34_chany_bottom_out[10] ,
    \sb_1__1__34_chany_bottom_out[11] ,
    \sb_1__1__34_chany_bottom_out[12] ,
    \sb_1__1__34_chany_bottom_out[13] ,
    \sb_1__1__34_chany_bottom_out[14] ,
    \sb_1__1__34_chany_bottom_out[15] ,
    \sb_1__1__34_chany_bottom_out[16] ,
    \sb_1__1__34_chany_bottom_out[17] ,
    \sb_1__1__34_chany_bottom_out[18] ,
    \sb_1__1__34_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__39_chany_bottom_out[0] ,
    \cby_1__1__39_chany_bottom_out[1] ,
    \cby_1__1__39_chany_bottom_out[2] ,
    \cby_1__1__39_chany_bottom_out[3] ,
    \cby_1__1__39_chany_bottom_out[4] ,
    \cby_1__1__39_chany_bottom_out[5] ,
    \cby_1__1__39_chany_bottom_out[6] ,
    \cby_1__1__39_chany_bottom_out[7] ,
    \cby_1__1__39_chany_bottom_out[8] ,
    \cby_1__1__39_chany_bottom_out[9] ,
    \cby_1__1__39_chany_bottom_out[10] ,
    \cby_1__1__39_chany_bottom_out[11] ,
    \cby_1__1__39_chany_bottom_out[12] ,
    \cby_1__1__39_chany_bottom_out[13] ,
    \cby_1__1__39_chany_bottom_out[14] ,
    \cby_1__1__39_chany_bottom_out[15] ,
    \cby_1__1__39_chany_bottom_out[16] ,
    \cby_1__1__39_chany_bottom_out[17] ,
    \cby_1__1__39_chany_bottom_out[18] ,
    \cby_1__1__39_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__34_chany_top_out[0] ,
    \sb_1__1__34_chany_top_out[1] ,
    \sb_1__1__34_chany_top_out[2] ,
    \sb_1__1__34_chany_top_out[3] ,
    \sb_1__1__34_chany_top_out[4] ,
    \sb_1__1__34_chany_top_out[5] ,
    \sb_1__1__34_chany_top_out[6] ,
    \sb_1__1__34_chany_top_out[7] ,
    \sb_1__1__34_chany_top_out[8] ,
    \sb_1__1__34_chany_top_out[9] ,
    \sb_1__1__34_chany_top_out[10] ,
    \sb_1__1__34_chany_top_out[11] ,
    \sb_1__1__34_chany_top_out[12] ,
    \sb_1__1__34_chany_top_out[13] ,
    \sb_1__1__34_chany_top_out[14] ,
    \sb_1__1__34_chany_top_out[15] ,
    \sb_1__1__34_chany_top_out[16] ,
    \sb_1__1__34_chany_top_out[17] ,
    \sb_1__1__34_chany_top_out[18] ,
    \sb_1__1__34_chany_top_out[19] }));
 sb_1__2_ sb_5__8_ (.bottom_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_upper),
    .ccff_head(grid_io_top_5_ccff_tail),
    .ccff_tail(sb_1__8__4_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[146] ),
    .right_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__4_chanx_right_out[0] ,
    \cbx_1__8__4_chanx_right_out[1] ,
    \cbx_1__8__4_chanx_right_out[2] ,
    \cbx_1__8__4_chanx_right_out[3] ,
    \cbx_1__8__4_chanx_right_out[4] ,
    \cbx_1__8__4_chanx_right_out[5] ,
    \cbx_1__8__4_chanx_right_out[6] ,
    \cbx_1__8__4_chanx_right_out[7] ,
    \cbx_1__8__4_chanx_right_out[8] ,
    \cbx_1__8__4_chanx_right_out[9] ,
    \cbx_1__8__4_chanx_right_out[10] ,
    \cbx_1__8__4_chanx_right_out[11] ,
    \cbx_1__8__4_chanx_right_out[12] ,
    \cbx_1__8__4_chanx_right_out[13] ,
    \cbx_1__8__4_chanx_right_out[14] ,
    \cbx_1__8__4_chanx_right_out[15] ,
    \cbx_1__8__4_chanx_right_out[16] ,
    \cbx_1__8__4_chanx_right_out[17] ,
    \cbx_1__8__4_chanx_right_out[18] ,
    \cbx_1__8__4_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__8__4_chanx_left_out[0] ,
    \sb_1__8__4_chanx_left_out[1] ,
    \sb_1__8__4_chanx_left_out[2] ,
    \sb_1__8__4_chanx_left_out[3] ,
    \sb_1__8__4_chanx_left_out[4] ,
    \sb_1__8__4_chanx_left_out[5] ,
    \sb_1__8__4_chanx_left_out[6] ,
    \sb_1__8__4_chanx_left_out[7] ,
    \sb_1__8__4_chanx_left_out[8] ,
    \sb_1__8__4_chanx_left_out[9] ,
    \sb_1__8__4_chanx_left_out[10] ,
    \sb_1__8__4_chanx_left_out[11] ,
    \sb_1__8__4_chanx_left_out[12] ,
    \sb_1__8__4_chanx_left_out[13] ,
    \sb_1__8__4_chanx_left_out[14] ,
    \sb_1__8__4_chanx_left_out[15] ,
    \sb_1__8__4_chanx_left_out[16] ,
    \sb_1__8__4_chanx_left_out[17] ,
    \sb_1__8__4_chanx_left_out[18] ,
    \sb_1__8__4_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__8__5_chanx_left_out[0] ,
    \cbx_1__8__5_chanx_left_out[1] ,
    \cbx_1__8__5_chanx_left_out[2] ,
    \cbx_1__8__5_chanx_left_out[3] ,
    \cbx_1__8__5_chanx_left_out[4] ,
    \cbx_1__8__5_chanx_left_out[5] ,
    \cbx_1__8__5_chanx_left_out[6] ,
    \cbx_1__8__5_chanx_left_out[7] ,
    \cbx_1__8__5_chanx_left_out[8] ,
    \cbx_1__8__5_chanx_left_out[9] ,
    \cbx_1__8__5_chanx_left_out[10] ,
    \cbx_1__8__5_chanx_left_out[11] ,
    \cbx_1__8__5_chanx_left_out[12] ,
    \cbx_1__8__5_chanx_left_out[13] ,
    \cbx_1__8__5_chanx_left_out[14] ,
    \cbx_1__8__5_chanx_left_out[15] ,
    \cbx_1__8__5_chanx_left_out[16] ,
    \cbx_1__8__5_chanx_left_out[17] ,
    \cbx_1__8__5_chanx_left_out[18] ,
    \cbx_1__8__5_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__8__4_chanx_right_out[0] ,
    \sb_1__8__4_chanx_right_out[1] ,
    \sb_1__8__4_chanx_right_out[2] ,
    \sb_1__8__4_chanx_right_out[3] ,
    \sb_1__8__4_chanx_right_out[4] ,
    \sb_1__8__4_chanx_right_out[5] ,
    \sb_1__8__4_chanx_right_out[6] ,
    \sb_1__8__4_chanx_right_out[7] ,
    \sb_1__8__4_chanx_right_out[8] ,
    \sb_1__8__4_chanx_right_out[9] ,
    \sb_1__8__4_chanx_right_out[10] ,
    \sb_1__8__4_chanx_right_out[11] ,
    \sb_1__8__4_chanx_right_out[12] ,
    \sb_1__8__4_chanx_right_out[13] ,
    \sb_1__8__4_chanx_right_out[14] ,
    \sb_1__8__4_chanx_right_out[15] ,
    \sb_1__8__4_chanx_right_out[16] ,
    \sb_1__8__4_chanx_right_out[17] ,
    \sb_1__8__4_chanx_right_out[18] ,
    \sb_1__8__4_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__39_chany_top_out[0] ,
    \cby_1__1__39_chany_top_out[1] ,
    \cby_1__1__39_chany_top_out[2] ,
    \cby_1__1__39_chany_top_out[3] ,
    \cby_1__1__39_chany_top_out[4] ,
    \cby_1__1__39_chany_top_out[5] ,
    \cby_1__1__39_chany_top_out[6] ,
    \cby_1__1__39_chany_top_out[7] ,
    \cby_1__1__39_chany_top_out[8] ,
    \cby_1__1__39_chany_top_out[9] ,
    \cby_1__1__39_chany_top_out[10] ,
    \cby_1__1__39_chany_top_out[11] ,
    \cby_1__1__39_chany_top_out[12] ,
    \cby_1__1__39_chany_top_out[13] ,
    \cby_1__1__39_chany_top_out[14] ,
    \cby_1__1__39_chany_top_out[15] ,
    \cby_1__1__39_chany_top_out[16] ,
    \cby_1__1__39_chany_top_out[17] ,
    \cby_1__1__39_chany_top_out[18] ,
    \cby_1__1__39_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__8__4_chany_bottom_out[0] ,
    \sb_1__8__4_chany_bottom_out[1] ,
    \sb_1__8__4_chany_bottom_out[2] ,
    \sb_1__8__4_chany_bottom_out[3] ,
    \sb_1__8__4_chany_bottom_out[4] ,
    \sb_1__8__4_chany_bottom_out[5] ,
    \sb_1__8__4_chany_bottom_out[6] ,
    \sb_1__8__4_chany_bottom_out[7] ,
    \sb_1__8__4_chany_bottom_out[8] ,
    \sb_1__8__4_chany_bottom_out[9] ,
    \sb_1__8__4_chany_bottom_out[10] ,
    \sb_1__8__4_chany_bottom_out[11] ,
    \sb_1__8__4_chany_bottom_out[12] ,
    \sb_1__8__4_chany_bottom_out[13] ,
    \sb_1__8__4_chany_bottom_out[14] ,
    \sb_1__8__4_chany_bottom_out[15] ,
    \sb_1__8__4_chany_bottom_out[16] ,
    \sb_1__8__4_chany_bottom_out[17] ,
    \sb_1__8__4_chany_bottom_out[18] ,
    \sb_1__8__4_chany_bottom_out[19] }));
 sb_1__0_ sb_6__0_ (.ccff_head(grid_io_bottom_1_ccff_tail),
    .ccff_tail(sb_1__0__5_ccff_tail),
    .left_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[149] ),
    .right_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__5_chanx_right_out[0] ,
    \cbx_1__0__5_chanx_right_out[1] ,
    \cbx_1__0__5_chanx_right_out[2] ,
    \cbx_1__0__5_chanx_right_out[3] ,
    \cbx_1__0__5_chanx_right_out[4] ,
    \cbx_1__0__5_chanx_right_out[5] ,
    \cbx_1__0__5_chanx_right_out[6] ,
    \cbx_1__0__5_chanx_right_out[7] ,
    \cbx_1__0__5_chanx_right_out[8] ,
    \cbx_1__0__5_chanx_right_out[9] ,
    \cbx_1__0__5_chanx_right_out[10] ,
    \cbx_1__0__5_chanx_right_out[11] ,
    \cbx_1__0__5_chanx_right_out[12] ,
    \cbx_1__0__5_chanx_right_out[13] ,
    \cbx_1__0__5_chanx_right_out[14] ,
    \cbx_1__0__5_chanx_right_out[15] ,
    \cbx_1__0__5_chanx_right_out[16] ,
    \cbx_1__0__5_chanx_right_out[17] ,
    \cbx_1__0__5_chanx_right_out[18] ,
    \cbx_1__0__5_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__0__5_chanx_left_out[0] ,
    \sb_1__0__5_chanx_left_out[1] ,
    \sb_1__0__5_chanx_left_out[2] ,
    \sb_1__0__5_chanx_left_out[3] ,
    \sb_1__0__5_chanx_left_out[4] ,
    \sb_1__0__5_chanx_left_out[5] ,
    \sb_1__0__5_chanx_left_out[6] ,
    \sb_1__0__5_chanx_left_out[7] ,
    \sb_1__0__5_chanx_left_out[8] ,
    \sb_1__0__5_chanx_left_out[9] ,
    \sb_1__0__5_chanx_left_out[10] ,
    \sb_1__0__5_chanx_left_out[11] ,
    \sb_1__0__5_chanx_left_out[12] ,
    \sb_1__0__5_chanx_left_out[13] ,
    \sb_1__0__5_chanx_left_out[14] ,
    \sb_1__0__5_chanx_left_out[15] ,
    \sb_1__0__5_chanx_left_out[16] ,
    \sb_1__0__5_chanx_left_out[17] ,
    \sb_1__0__5_chanx_left_out[18] ,
    \sb_1__0__5_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__0__6_chanx_left_out[0] ,
    \cbx_1__0__6_chanx_left_out[1] ,
    \cbx_1__0__6_chanx_left_out[2] ,
    \cbx_1__0__6_chanx_left_out[3] ,
    \cbx_1__0__6_chanx_left_out[4] ,
    \cbx_1__0__6_chanx_left_out[5] ,
    \cbx_1__0__6_chanx_left_out[6] ,
    \cbx_1__0__6_chanx_left_out[7] ,
    \cbx_1__0__6_chanx_left_out[8] ,
    \cbx_1__0__6_chanx_left_out[9] ,
    \cbx_1__0__6_chanx_left_out[10] ,
    \cbx_1__0__6_chanx_left_out[11] ,
    \cbx_1__0__6_chanx_left_out[12] ,
    \cbx_1__0__6_chanx_left_out[13] ,
    \cbx_1__0__6_chanx_left_out[14] ,
    \cbx_1__0__6_chanx_left_out[15] ,
    \cbx_1__0__6_chanx_left_out[16] ,
    \cbx_1__0__6_chanx_left_out[17] ,
    \cbx_1__0__6_chanx_left_out[18] ,
    \cbx_1__0__6_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__0__5_chanx_right_out[0] ,
    \sb_1__0__5_chanx_right_out[1] ,
    \sb_1__0__5_chanx_right_out[2] ,
    \sb_1__0__5_chanx_right_out[3] ,
    \sb_1__0__5_chanx_right_out[4] ,
    \sb_1__0__5_chanx_right_out[5] ,
    \sb_1__0__5_chanx_right_out[6] ,
    \sb_1__0__5_chanx_right_out[7] ,
    \sb_1__0__5_chanx_right_out[8] ,
    \sb_1__0__5_chanx_right_out[9] ,
    \sb_1__0__5_chanx_right_out[10] ,
    \sb_1__0__5_chanx_right_out[11] ,
    \sb_1__0__5_chanx_right_out[12] ,
    \sb_1__0__5_chanx_right_out[13] ,
    \sb_1__0__5_chanx_right_out[14] ,
    \sb_1__0__5_chanx_right_out[15] ,
    \sb_1__0__5_chanx_right_out[16] ,
    \sb_1__0__5_chanx_right_out[17] ,
    \sb_1__0__5_chanx_right_out[18] ,
    \sb_1__0__5_chanx_right_out[19] }),
    .chany_top_in({\cby_1__1__40_chany_bottom_out[0] ,
    \cby_1__1__40_chany_bottom_out[1] ,
    \cby_1__1__40_chany_bottom_out[2] ,
    \cby_1__1__40_chany_bottom_out[3] ,
    \cby_1__1__40_chany_bottom_out[4] ,
    \cby_1__1__40_chany_bottom_out[5] ,
    \cby_1__1__40_chany_bottom_out[6] ,
    \cby_1__1__40_chany_bottom_out[7] ,
    \cby_1__1__40_chany_bottom_out[8] ,
    \cby_1__1__40_chany_bottom_out[9] ,
    \cby_1__1__40_chany_bottom_out[10] ,
    \cby_1__1__40_chany_bottom_out[11] ,
    \cby_1__1__40_chany_bottom_out[12] ,
    \cby_1__1__40_chany_bottom_out[13] ,
    \cby_1__1__40_chany_bottom_out[14] ,
    \cby_1__1__40_chany_bottom_out[15] ,
    \cby_1__1__40_chany_bottom_out[16] ,
    \cby_1__1__40_chany_bottom_out[17] ,
    \cby_1__1__40_chany_bottom_out[18] ,
    \cby_1__1__40_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__0__5_chany_top_out[0] ,
    \sb_1__0__5_chany_top_out[1] ,
    \sb_1__0__5_chany_top_out[2] ,
    \sb_1__0__5_chany_top_out[3] ,
    \sb_1__0__5_chany_top_out[4] ,
    \sb_1__0__5_chany_top_out[5] ,
    \sb_1__0__5_chany_top_out[6] ,
    \sb_1__0__5_chany_top_out[7] ,
    \sb_1__0__5_chany_top_out[8] ,
    \sb_1__0__5_chany_top_out[9] ,
    \sb_1__0__5_chany_top_out[10] ,
    \sb_1__0__5_chany_top_out[11] ,
    \sb_1__0__5_chany_top_out[12] ,
    \sb_1__0__5_chany_top_out[13] ,
    \sb_1__0__5_chany_top_out[14] ,
    \sb_1__0__5_chany_top_out[15] ,
    \sb_1__0__5_chany_top_out[16] ,
    \sb_1__0__5_chany_top_out[17] ,
    \sb_1__0__5_chany_top_out[18] ,
    \sb_1__0__5_chany_top_out[19] }));
 sb_1__1_ sb_6__1_ (.bottom_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__42_ccff_tail),
    .ccff_tail(sb_1__1__35_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[152] ),
    .right_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__35_chanx_right_out[0] ,
    \cbx_1__1__35_chanx_right_out[1] ,
    \cbx_1__1__35_chanx_right_out[2] ,
    \cbx_1__1__35_chanx_right_out[3] ,
    \cbx_1__1__35_chanx_right_out[4] ,
    \cbx_1__1__35_chanx_right_out[5] ,
    \cbx_1__1__35_chanx_right_out[6] ,
    \cbx_1__1__35_chanx_right_out[7] ,
    \cbx_1__1__35_chanx_right_out[8] ,
    \cbx_1__1__35_chanx_right_out[9] ,
    \cbx_1__1__35_chanx_right_out[10] ,
    \cbx_1__1__35_chanx_right_out[11] ,
    \cbx_1__1__35_chanx_right_out[12] ,
    \cbx_1__1__35_chanx_right_out[13] ,
    \cbx_1__1__35_chanx_right_out[14] ,
    \cbx_1__1__35_chanx_right_out[15] ,
    \cbx_1__1__35_chanx_right_out[16] ,
    \cbx_1__1__35_chanx_right_out[17] ,
    \cbx_1__1__35_chanx_right_out[18] ,
    \cbx_1__1__35_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__35_chanx_left_out[0] ,
    \sb_1__1__35_chanx_left_out[1] ,
    \sb_1__1__35_chanx_left_out[2] ,
    \sb_1__1__35_chanx_left_out[3] ,
    \sb_1__1__35_chanx_left_out[4] ,
    \sb_1__1__35_chanx_left_out[5] ,
    \sb_1__1__35_chanx_left_out[6] ,
    \sb_1__1__35_chanx_left_out[7] ,
    \sb_1__1__35_chanx_left_out[8] ,
    \sb_1__1__35_chanx_left_out[9] ,
    \sb_1__1__35_chanx_left_out[10] ,
    \sb_1__1__35_chanx_left_out[11] ,
    \sb_1__1__35_chanx_left_out[12] ,
    \sb_1__1__35_chanx_left_out[13] ,
    \sb_1__1__35_chanx_left_out[14] ,
    \sb_1__1__35_chanx_left_out[15] ,
    \sb_1__1__35_chanx_left_out[16] ,
    \sb_1__1__35_chanx_left_out[17] ,
    \sb_1__1__35_chanx_left_out[18] ,
    \sb_1__1__35_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__42_chanx_left_out[0] ,
    \cbx_1__1__42_chanx_left_out[1] ,
    \cbx_1__1__42_chanx_left_out[2] ,
    \cbx_1__1__42_chanx_left_out[3] ,
    \cbx_1__1__42_chanx_left_out[4] ,
    \cbx_1__1__42_chanx_left_out[5] ,
    \cbx_1__1__42_chanx_left_out[6] ,
    \cbx_1__1__42_chanx_left_out[7] ,
    \cbx_1__1__42_chanx_left_out[8] ,
    \cbx_1__1__42_chanx_left_out[9] ,
    \cbx_1__1__42_chanx_left_out[10] ,
    \cbx_1__1__42_chanx_left_out[11] ,
    \cbx_1__1__42_chanx_left_out[12] ,
    \cbx_1__1__42_chanx_left_out[13] ,
    \cbx_1__1__42_chanx_left_out[14] ,
    \cbx_1__1__42_chanx_left_out[15] ,
    \cbx_1__1__42_chanx_left_out[16] ,
    \cbx_1__1__42_chanx_left_out[17] ,
    \cbx_1__1__42_chanx_left_out[18] ,
    \cbx_1__1__42_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__35_chanx_right_out[0] ,
    \sb_1__1__35_chanx_right_out[1] ,
    \sb_1__1__35_chanx_right_out[2] ,
    \sb_1__1__35_chanx_right_out[3] ,
    \sb_1__1__35_chanx_right_out[4] ,
    \sb_1__1__35_chanx_right_out[5] ,
    \sb_1__1__35_chanx_right_out[6] ,
    \sb_1__1__35_chanx_right_out[7] ,
    \sb_1__1__35_chanx_right_out[8] ,
    \sb_1__1__35_chanx_right_out[9] ,
    \sb_1__1__35_chanx_right_out[10] ,
    \sb_1__1__35_chanx_right_out[11] ,
    \sb_1__1__35_chanx_right_out[12] ,
    \sb_1__1__35_chanx_right_out[13] ,
    \sb_1__1__35_chanx_right_out[14] ,
    \sb_1__1__35_chanx_right_out[15] ,
    \sb_1__1__35_chanx_right_out[16] ,
    \sb_1__1__35_chanx_right_out[17] ,
    \sb_1__1__35_chanx_right_out[18] ,
    \sb_1__1__35_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__40_chany_top_out[0] ,
    \cby_1__1__40_chany_top_out[1] ,
    \cby_1__1__40_chany_top_out[2] ,
    \cby_1__1__40_chany_top_out[3] ,
    \cby_1__1__40_chany_top_out[4] ,
    \cby_1__1__40_chany_top_out[5] ,
    \cby_1__1__40_chany_top_out[6] ,
    \cby_1__1__40_chany_top_out[7] ,
    \cby_1__1__40_chany_top_out[8] ,
    \cby_1__1__40_chany_top_out[9] ,
    \cby_1__1__40_chany_top_out[10] ,
    \cby_1__1__40_chany_top_out[11] ,
    \cby_1__1__40_chany_top_out[12] ,
    \cby_1__1__40_chany_top_out[13] ,
    \cby_1__1__40_chany_top_out[14] ,
    \cby_1__1__40_chany_top_out[15] ,
    \cby_1__1__40_chany_top_out[16] ,
    \cby_1__1__40_chany_top_out[17] ,
    \cby_1__1__40_chany_top_out[18] ,
    \cby_1__1__40_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__35_chany_bottom_out[0] ,
    \sb_1__1__35_chany_bottom_out[1] ,
    \sb_1__1__35_chany_bottom_out[2] ,
    \sb_1__1__35_chany_bottom_out[3] ,
    \sb_1__1__35_chany_bottom_out[4] ,
    \sb_1__1__35_chany_bottom_out[5] ,
    \sb_1__1__35_chany_bottom_out[6] ,
    \sb_1__1__35_chany_bottom_out[7] ,
    \sb_1__1__35_chany_bottom_out[8] ,
    \sb_1__1__35_chany_bottom_out[9] ,
    \sb_1__1__35_chany_bottom_out[10] ,
    \sb_1__1__35_chany_bottom_out[11] ,
    \sb_1__1__35_chany_bottom_out[12] ,
    \sb_1__1__35_chany_bottom_out[13] ,
    \sb_1__1__35_chany_bottom_out[14] ,
    \sb_1__1__35_chany_bottom_out[15] ,
    \sb_1__1__35_chany_bottom_out[16] ,
    \sb_1__1__35_chany_bottom_out[17] ,
    \sb_1__1__35_chany_bottom_out[18] ,
    \sb_1__1__35_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__41_chany_bottom_out[0] ,
    \cby_1__1__41_chany_bottom_out[1] ,
    \cby_1__1__41_chany_bottom_out[2] ,
    \cby_1__1__41_chany_bottom_out[3] ,
    \cby_1__1__41_chany_bottom_out[4] ,
    \cby_1__1__41_chany_bottom_out[5] ,
    \cby_1__1__41_chany_bottom_out[6] ,
    \cby_1__1__41_chany_bottom_out[7] ,
    \cby_1__1__41_chany_bottom_out[8] ,
    \cby_1__1__41_chany_bottom_out[9] ,
    \cby_1__1__41_chany_bottom_out[10] ,
    \cby_1__1__41_chany_bottom_out[11] ,
    \cby_1__1__41_chany_bottom_out[12] ,
    \cby_1__1__41_chany_bottom_out[13] ,
    \cby_1__1__41_chany_bottom_out[14] ,
    \cby_1__1__41_chany_bottom_out[15] ,
    \cby_1__1__41_chany_bottom_out[16] ,
    \cby_1__1__41_chany_bottom_out[17] ,
    \cby_1__1__41_chany_bottom_out[18] ,
    \cby_1__1__41_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__35_chany_top_out[0] ,
    \sb_1__1__35_chany_top_out[1] ,
    \sb_1__1__35_chany_top_out[2] ,
    \sb_1__1__35_chany_top_out[3] ,
    \sb_1__1__35_chany_top_out[4] ,
    \sb_1__1__35_chany_top_out[5] ,
    \sb_1__1__35_chany_top_out[6] ,
    \sb_1__1__35_chany_top_out[7] ,
    \sb_1__1__35_chany_top_out[8] ,
    \sb_1__1__35_chany_top_out[9] ,
    \sb_1__1__35_chany_top_out[10] ,
    \sb_1__1__35_chany_top_out[11] ,
    \sb_1__1__35_chany_top_out[12] ,
    \sb_1__1__35_chany_top_out[13] ,
    \sb_1__1__35_chany_top_out[14] ,
    \sb_1__1__35_chany_top_out[15] ,
    \sb_1__1__35_chany_top_out[16] ,
    \sb_1__1__35_chany_top_out[17] ,
    \sb_1__1__35_chany_top_out[18] ,
    \sb_1__1__35_chany_top_out[19] }));
 sb_1__1_ sb_6__2_ (.bottom_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__43_ccff_tail),
    .ccff_tail(sb_1__1__36_ccff_tail),
    .clk_2_E_out(\clk_2_wires[27] ),
    .clk_2_N_in(\clk_3_wires[25] ),
    .clk_2_W_out(\clk_2_wires[29] ),
    .left_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[155] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[27] ),
    .prog_clk_2_N_in(\prog_clk_3_wires[25] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[29] ),
    .right_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__36_chanx_right_out[0] ,
    \cbx_1__1__36_chanx_right_out[1] ,
    \cbx_1__1__36_chanx_right_out[2] ,
    \cbx_1__1__36_chanx_right_out[3] ,
    \cbx_1__1__36_chanx_right_out[4] ,
    \cbx_1__1__36_chanx_right_out[5] ,
    \cbx_1__1__36_chanx_right_out[6] ,
    \cbx_1__1__36_chanx_right_out[7] ,
    \cbx_1__1__36_chanx_right_out[8] ,
    \cbx_1__1__36_chanx_right_out[9] ,
    \cbx_1__1__36_chanx_right_out[10] ,
    \cbx_1__1__36_chanx_right_out[11] ,
    \cbx_1__1__36_chanx_right_out[12] ,
    \cbx_1__1__36_chanx_right_out[13] ,
    \cbx_1__1__36_chanx_right_out[14] ,
    \cbx_1__1__36_chanx_right_out[15] ,
    \cbx_1__1__36_chanx_right_out[16] ,
    \cbx_1__1__36_chanx_right_out[17] ,
    \cbx_1__1__36_chanx_right_out[18] ,
    \cbx_1__1__36_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__36_chanx_left_out[0] ,
    \sb_1__1__36_chanx_left_out[1] ,
    \sb_1__1__36_chanx_left_out[2] ,
    \sb_1__1__36_chanx_left_out[3] ,
    \sb_1__1__36_chanx_left_out[4] ,
    \sb_1__1__36_chanx_left_out[5] ,
    \sb_1__1__36_chanx_left_out[6] ,
    \sb_1__1__36_chanx_left_out[7] ,
    \sb_1__1__36_chanx_left_out[8] ,
    \sb_1__1__36_chanx_left_out[9] ,
    \sb_1__1__36_chanx_left_out[10] ,
    \sb_1__1__36_chanx_left_out[11] ,
    \sb_1__1__36_chanx_left_out[12] ,
    \sb_1__1__36_chanx_left_out[13] ,
    \sb_1__1__36_chanx_left_out[14] ,
    \sb_1__1__36_chanx_left_out[15] ,
    \sb_1__1__36_chanx_left_out[16] ,
    \sb_1__1__36_chanx_left_out[17] ,
    \sb_1__1__36_chanx_left_out[18] ,
    \sb_1__1__36_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__43_chanx_left_out[0] ,
    \cbx_1__1__43_chanx_left_out[1] ,
    \cbx_1__1__43_chanx_left_out[2] ,
    \cbx_1__1__43_chanx_left_out[3] ,
    \cbx_1__1__43_chanx_left_out[4] ,
    \cbx_1__1__43_chanx_left_out[5] ,
    \cbx_1__1__43_chanx_left_out[6] ,
    \cbx_1__1__43_chanx_left_out[7] ,
    \cbx_1__1__43_chanx_left_out[8] ,
    \cbx_1__1__43_chanx_left_out[9] ,
    \cbx_1__1__43_chanx_left_out[10] ,
    \cbx_1__1__43_chanx_left_out[11] ,
    \cbx_1__1__43_chanx_left_out[12] ,
    \cbx_1__1__43_chanx_left_out[13] ,
    \cbx_1__1__43_chanx_left_out[14] ,
    \cbx_1__1__43_chanx_left_out[15] ,
    \cbx_1__1__43_chanx_left_out[16] ,
    \cbx_1__1__43_chanx_left_out[17] ,
    \cbx_1__1__43_chanx_left_out[18] ,
    \cbx_1__1__43_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__36_chanx_right_out[0] ,
    \sb_1__1__36_chanx_right_out[1] ,
    \sb_1__1__36_chanx_right_out[2] ,
    \sb_1__1__36_chanx_right_out[3] ,
    \sb_1__1__36_chanx_right_out[4] ,
    \sb_1__1__36_chanx_right_out[5] ,
    \sb_1__1__36_chanx_right_out[6] ,
    \sb_1__1__36_chanx_right_out[7] ,
    \sb_1__1__36_chanx_right_out[8] ,
    \sb_1__1__36_chanx_right_out[9] ,
    \sb_1__1__36_chanx_right_out[10] ,
    \sb_1__1__36_chanx_right_out[11] ,
    \sb_1__1__36_chanx_right_out[12] ,
    \sb_1__1__36_chanx_right_out[13] ,
    \sb_1__1__36_chanx_right_out[14] ,
    \sb_1__1__36_chanx_right_out[15] ,
    \sb_1__1__36_chanx_right_out[16] ,
    \sb_1__1__36_chanx_right_out[17] ,
    \sb_1__1__36_chanx_right_out[18] ,
    \sb_1__1__36_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__41_chany_top_out[0] ,
    \cby_1__1__41_chany_top_out[1] ,
    \cby_1__1__41_chany_top_out[2] ,
    \cby_1__1__41_chany_top_out[3] ,
    \cby_1__1__41_chany_top_out[4] ,
    \cby_1__1__41_chany_top_out[5] ,
    \cby_1__1__41_chany_top_out[6] ,
    \cby_1__1__41_chany_top_out[7] ,
    \cby_1__1__41_chany_top_out[8] ,
    \cby_1__1__41_chany_top_out[9] ,
    \cby_1__1__41_chany_top_out[10] ,
    \cby_1__1__41_chany_top_out[11] ,
    \cby_1__1__41_chany_top_out[12] ,
    \cby_1__1__41_chany_top_out[13] ,
    \cby_1__1__41_chany_top_out[14] ,
    \cby_1__1__41_chany_top_out[15] ,
    \cby_1__1__41_chany_top_out[16] ,
    \cby_1__1__41_chany_top_out[17] ,
    \cby_1__1__41_chany_top_out[18] ,
    \cby_1__1__41_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__36_chany_bottom_out[0] ,
    \sb_1__1__36_chany_bottom_out[1] ,
    \sb_1__1__36_chany_bottom_out[2] ,
    \sb_1__1__36_chany_bottom_out[3] ,
    \sb_1__1__36_chany_bottom_out[4] ,
    \sb_1__1__36_chany_bottom_out[5] ,
    \sb_1__1__36_chany_bottom_out[6] ,
    \sb_1__1__36_chany_bottom_out[7] ,
    \sb_1__1__36_chany_bottom_out[8] ,
    \sb_1__1__36_chany_bottom_out[9] ,
    \sb_1__1__36_chany_bottom_out[10] ,
    \sb_1__1__36_chany_bottom_out[11] ,
    \sb_1__1__36_chany_bottom_out[12] ,
    \sb_1__1__36_chany_bottom_out[13] ,
    \sb_1__1__36_chany_bottom_out[14] ,
    \sb_1__1__36_chany_bottom_out[15] ,
    \sb_1__1__36_chany_bottom_out[16] ,
    \sb_1__1__36_chany_bottom_out[17] ,
    \sb_1__1__36_chany_bottom_out[18] ,
    \sb_1__1__36_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__42_chany_bottom_out[0] ,
    \cby_1__1__42_chany_bottom_out[1] ,
    \cby_1__1__42_chany_bottom_out[2] ,
    \cby_1__1__42_chany_bottom_out[3] ,
    \cby_1__1__42_chany_bottom_out[4] ,
    \cby_1__1__42_chany_bottom_out[5] ,
    \cby_1__1__42_chany_bottom_out[6] ,
    \cby_1__1__42_chany_bottom_out[7] ,
    \cby_1__1__42_chany_bottom_out[8] ,
    \cby_1__1__42_chany_bottom_out[9] ,
    \cby_1__1__42_chany_bottom_out[10] ,
    \cby_1__1__42_chany_bottom_out[11] ,
    \cby_1__1__42_chany_bottom_out[12] ,
    \cby_1__1__42_chany_bottom_out[13] ,
    \cby_1__1__42_chany_bottom_out[14] ,
    \cby_1__1__42_chany_bottom_out[15] ,
    \cby_1__1__42_chany_bottom_out[16] ,
    \cby_1__1__42_chany_bottom_out[17] ,
    \cby_1__1__42_chany_bottom_out[18] ,
    \cby_1__1__42_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__36_chany_top_out[0] ,
    \sb_1__1__36_chany_top_out[1] ,
    \sb_1__1__36_chany_top_out[2] ,
    \sb_1__1__36_chany_top_out[3] ,
    \sb_1__1__36_chany_top_out[4] ,
    \sb_1__1__36_chany_top_out[5] ,
    \sb_1__1__36_chany_top_out[6] ,
    \sb_1__1__36_chany_top_out[7] ,
    \sb_1__1__36_chany_top_out[8] ,
    \sb_1__1__36_chany_top_out[9] ,
    \sb_1__1__36_chany_top_out[10] ,
    \sb_1__1__36_chany_top_out[11] ,
    \sb_1__1__36_chany_top_out[12] ,
    \sb_1__1__36_chany_top_out[13] ,
    \sb_1__1__36_chany_top_out[14] ,
    \sb_1__1__36_chany_top_out[15] ,
    \sb_1__1__36_chany_top_out[16] ,
    \sb_1__1__36_chany_top_out[17] ,
    \sb_1__1__36_chany_top_out[18] ,
    \sb_1__1__36_chany_top_out[19] }));
 sb_1__1_ sb_6__3_ (.bottom_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__44_ccff_tail),
    .ccff_tail(sb_1__1__37_ccff_tail),
    .clk_3_N_in(\clk_3_wires[21] ),
    .clk_3_S_out(\clk_3_wires[24] ),
    .left_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[158] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[21] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[24] ),
    .right_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__37_chanx_right_out[0] ,
    \cbx_1__1__37_chanx_right_out[1] ,
    \cbx_1__1__37_chanx_right_out[2] ,
    \cbx_1__1__37_chanx_right_out[3] ,
    \cbx_1__1__37_chanx_right_out[4] ,
    \cbx_1__1__37_chanx_right_out[5] ,
    \cbx_1__1__37_chanx_right_out[6] ,
    \cbx_1__1__37_chanx_right_out[7] ,
    \cbx_1__1__37_chanx_right_out[8] ,
    \cbx_1__1__37_chanx_right_out[9] ,
    \cbx_1__1__37_chanx_right_out[10] ,
    \cbx_1__1__37_chanx_right_out[11] ,
    \cbx_1__1__37_chanx_right_out[12] ,
    \cbx_1__1__37_chanx_right_out[13] ,
    \cbx_1__1__37_chanx_right_out[14] ,
    \cbx_1__1__37_chanx_right_out[15] ,
    \cbx_1__1__37_chanx_right_out[16] ,
    \cbx_1__1__37_chanx_right_out[17] ,
    \cbx_1__1__37_chanx_right_out[18] ,
    \cbx_1__1__37_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__37_chanx_left_out[0] ,
    \sb_1__1__37_chanx_left_out[1] ,
    \sb_1__1__37_chanx_left_out[2] ,
    \sb_1__1__37_chanx_left_out[3] ,
    \sb_1__1__37_chanx_left_out[4] ,
    \sb_1__1__37_chanx_left_out[5] ,
    \sb_1__1__37_chanx_left_out[6] ,
    \sb_1__1__37_chanx_left_out[7] ,
    \sb_1__1__37_chanx_left_out[8] ,
    \sb_1__1__37_chanx_left_out[9] ,
    \sb_1__1__37_chanx_left_out[10] ,
    \sb_1__1__37_chanx_left_out[11] ,
    \sb_1__1__37_chanx_left_out[12] ,
    \sb_1__1__37_chanx_left_out[13] ,
    \sb_1__1__37_chanx_left_out[14] ,
    \sb_1__1__37_chanx_left_out[15] ,
    \sb_1__1__37_chanx_left_out[16] ,
    \sb_1__1__37_chanx_left_out[17] ,
    \sb_1__1__37_chanx_left_out[18] ,
    \sb_1__1__37_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__44_chanx_left_out[0] ,
    \cbx_1__1__44_chanx_left_out[1] ,
    \cbx_1__1__44_chanx_left_out[2] ,
    \cbx_1__1__44_chanx_left_out[3] ,
    \cbx_1__1__44_chanx_left_out[4] ,
    \cbx_1__1__44_chanx_left_out[5] ,
    \cbx_1__1__44_chanx_left_out[6] ,
    \cbx_1__1__44_chanx_left_out[7] ,
    \cbx_1__1__44_chanx_left_out[8] ,
    \cbx_1__1__44_chanx_left_out[9] ,
    \cbx_1__1__44_chanx_left_out[10] ,
    \cbx_1__1__44_chanx_left_out[11] ,
    \cbx_1__1__44_chanx_left_out[12] ,
    \cbx_1__1__44_chanx_left_out[13] ,
    \cbx_1__1__44_chanx_left_out[14] ,
    \cbx_1__1__44_chanx_left_out[15] ,
    \cbx_1__1__44_chanx_left_out[16] ,
    \cbx_1__1__44_chanx_left_out[17] ,
    \cbx_1__1__44_chanx_left_out[18] ,
    \cbx_1__1__44_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__37_chanx_right_out[0] ,
    \sb_1__1__37_chanx_right_out[1] ,
    \sb_1__1__37_chanx_right_out[2] ,
    \sb_1__1__37_chanx_right_out[3] ,
    \sb_1__1__37_chanx_right_out[4] ,
    \sb_1__1__37_chanx_right_out[5] ,
    \sb_1__1__37_chanx_right_out[6] ,
    \sb_1__1__37_chanx_right_out[7] ,
    \sb_1__1__37_chanx_right_out[8] ,
    \sb_1__1__37_chanx_right_out[9] ,
    \sb_1__1__37_chanx_right_out[10] ,
    \sb_1__1__37_chanx_right_out[11] ,
    \sb_1__1__37_chanx_right_out[12] ,
    \sb_1__1__37_chanx_right_out[13] ,
    \sb_1__1__37_chanx_right_out[14] ,
    \sb_1__1__37_chanx_right_out[15] ,
    \sb_1__1__37_chanx_right_out[16] ,
    \sb_1__1__37_chanx_right_out[17] ,
    \sb_1__1__37_chanx_right_out[18] ,
    \sb_1__1__37_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__42_chany_top_out[0] ,
    \cby_1__1__42_chany_top_out[1] ,
    \cby_1__1__42_chany_top_out[2] ,
    \cby_1__1__42_chany_top_out[3] ,
    \cby_1__1__42_chany_top_out[4] ,
    \cby_1__1__42_chany_top_out[5] ,
    \cby_1__1__42_chany_top_out[6] ,
    \cby_1__1__42_chany_top_out[7] ,
    \cby_1__1__42_chany_top_out[8] ,
    \cby_1__1__42_chany_top_out[9] ,
    \cby_1__1__42_chany_top_out[10] ,
    \cby_1__1__42_chany_top_out[11] ,
    \cby_1__1__42_chany_top_out[12] ,
    \cby_1__1__42_chany_top_out[13] ,
    \cby_1__1__42_chany_top_out[14] ,
    \cby_1__1__42_chany_top_out[15] ,
    \cby_1__1__42_chany_top_out[16] ,
    \cby_1__1__42_chany_top_out[17] ,
    \cby_1__1__42_chany_top_out[18] ,
    \cby_1__1__42_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__37_chany_bottom_out[0] ,
    \sb_1__1__37_chany_bottom_out[1] ,
    \sb_1__1__37_chany_bottom_out[2] ,
    \sb_1__1__37_chany_bottom_out[3] ,
    \sb_1__1__37_chany_bottom_out[4] ,
    \sb_1__1__37_chany_bottom_out[5] ,
    \sb_1__1__37_chany_bottom_out[6] ,
    \sb_1__1__37_chany_bottom_out[7] ,
    \sb_1__1__37_chany_bottom_out[8] ,
    \sb_1__1__37_chany_bottom_out[9] ,
    \sb_1__1__37_chany_bottom_out[10] ,
    \sb_1__1__37_chany_bottom_out[11] ,
    \sb_1__1__37_chany_bottom_out[12] ,
    \sb_1__1__37_chany_bottom_out[13] ,
    \sb_1__1__37_chany_bottom_out[14] ,
    \sb_1__1__37_chany_bottom_out[15] ,
    \sb_1__1__37_chany_bottom_out[16] ,
    \sb_1__1__37_chany_bottom_out[17] ,
    \sb_1__1__37_chany_bottom_out[18] ,
    \sb_1__1__37_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__43_chany_bottom_out[0] ,
    \cby_1__1__43_chany_bottom_out[1] ,
    \cby_1__1__43_chany_bottom_out[2] ,
    \cby_1__1__43_chany_bottom_out[3] ,
    \cby_1__1__43_chany_bottom_out[4] ,
    \cby_1__1__43_chany_bottom_out[5] ,
    \cby_1__1__43_chany_bottom_out[6] ,
    \cby_1__1__43_chany_bottom_out[7] ,
    \cby_1__1__43_chany_bottom_out[8] ,
    \cby_1__1__43_chany_bottom_out[9] ,
    \cby_1__1__43_chany_bottom_out[10] ,
    \cby_1__1__43_chany_bottom_out[11] ,
    \cby_1__1__43_chany_bottom_out[12] ,
    \cby_1__1__43_chany_bottom_out[13] ,
    \cby_1__1__43_chany_bottom_out[14] ,
    \cby_1__1__43_chany_bottom_out[15] ,
    \cby_1__1__43_chany_bottom_out[16] ,
    \cby_1__1__43_chany_bottom_out[17] ,
    \cby_1__1__43_chany_bottom_out[18] ,
    \cby_1__1__43_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__37_chany_top_out[0] ,
    \sb_1__1__37_chany_top_out[1] ,
    \sb_1__1__37_chany_top_out[2] ,
    \sb_1__1__37_chany_top_out[3] ,
    \sb_1__1__37_chany_top_out[4] ,
    \sb_1__1__37_chany_top_out[5] ,
    \sb_1__1__37_chany_top_out[6] ,
    \sb_1__1__37_chany_top_out[7] ,
    \sb_1__1__37_chany_top_out[8] ,
    \sb_1__1__37_chany_top_out[9] ,
    \sb_1__1__37_chany_top_out[10] ,
    \sb_1__1__37_chany_top_out[11] ,
    \sb_1__1__37_chany_top_out[12] ,
    \sb_1__1__37_chany_top_out[13] ,
    \sb_1__1__37_chany_top_out[14] ,
    \sb_1__1__37_chany_top_out[15] ,
    \sb_1__1__37_chany_top_out[16] ,
    \sb_1__1__37_chany_top_out[17] ,
    \sb_1__1__37_chany_top_out[18] ,
    \sb_1__1__37_chany_top_out[19] }));
 sb_1__1_ sb_6__4_ (.bottom_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__45_ccff_tail),
    .ccff_tail(sb_1__1__38_ccff_tail),
    .clk_3_N_in(\clk_3_wires[7] ),
    .clk_3_N_out(\clk_3_wires[18] ),
    .clk_3_S_out(\clk_3_wires[20] ),
    .left_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[161] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[7] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[18] ),
    .prog_clk_3_S_out(\prog_clk_3_wires[20] ),
    .right_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__38_chanx_right_out[0] ,
    \cbx_1__1__38_chanx_right_out[1] ,
    \cbx_1__1__38_chanx_right_out[2] ,
    \cbx_1__1__38_chanx_right_out[3] ,
    \cbx_1__1__38_chanx_right_out[4] ,
    \cbx_1__1__38_chanx_right_out[5] ,
    \cbx_1__1__38_chanx_right_out[6] ,
    \cbx_1__1__38_chanx_right_out[7] ,
    \cbx_1__1__38_chanx_right_out[8] ,
    \cbx_1__1__38_chanx_right_out[9] ,
    \cbx_1__1__38_chanx_right_out[10] ,
    \cbx_1__1__38_chanx_right_out[11] ,
    \cbx_1__1__38_chanx_right_out[12] ,
    \cbx_1__1__38_chanx_right_out[13] ,
    \cbx_1__1__38_chanx_right_out[14] ,
    \cbx_1__1__38_chanx_right_out[15] ,
    \cbx_1__1__38_chanx_right_out[16] ,
    \cbx_1__1__38_chanx_right_out[17] ,
    \cbx_1__1__38_chanx_right_out[18] ,
    \cbx_1__1__38_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__38_chanx_left_out[0] ,
    \sb_1__1__38_chanx_left_out[1] ,
    \sb_1__1__38_chanx_left_out[2] ,
    \sb_1__1__38_chanx_left_out[3] ,
    \sb_1__1__38_chanx_left_out[4] ,
    \sb_1__1__38_chanx_left_out[5] ,
    \sb_1__1__38_chanx_left_out[6] ,
    \sb_1__1__38_chanx_left_out[7] ,
    \sb_1__1__38_chanx_left_out[8] ,
    \sb_1__1__38_chanx_left_out[9] ,
    \sb_1__1__38_chanx_left_out[10] ,
    \sb_1__1__38_chanx_left_out[11] ,
    \sb_1__1__38_chanx_left_out[12] ,
    \sb_1__1__38_chanx_left_out[13] ,
    \sb_1__1__38_chanx_left_out[14] ,
    \sb_1__1__38_chanx_left_out[15] ,
    \sb_1__1__38_chanx_left_out[16] ,
    \sb_1__1__38_chanx_left_out[17] ,
    \sb_1__1__38_chanx_left_out[18] ,
    \sb_1__1__38_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__45_chanx_left_out[0] ,
    \cbx_1__1__45_chanx_left_out[1] ,
    \cbx_1__1__45_chanx_left_out[2] ,
    \cbx_1__1__45_chanx_left_out[3] ,
    \cbx_1__1__45_chanx_left_out[4] ,
    \cbx_1__1__45_chanx_left_out[5] ,
    \cbx_1__1__45_chanx_left_out[6] ,
    \cbx_1__1__45_chanx_left_out[7] ,
    \cbx_1__1__45_chanx_left_out[8] ,
    \cbx_1__1__45_chanx_left_out[9] ,
    \cbx_1__1__45_chanx_left_out[10] ,
    \cbx_1__1__45_chanx_left_out[11] ,
    \cbx_1__1__45_chanx_left_out[12] ,
    \cbx_1__1__45_chanx_left_out[13] ,
    \cbx_1__1__45_chanx_left_out[14] ,
    \cbx_1__1__45_chanx_left_out[15] ,
    \cbx_1__1__45_chanx_left_out[16] ,
    \cbx_1__1__45_chanx_left_out[17] ,
    \cbx_1__1__45_chanx_left_out[18] ,
    \cbx_1__1__45_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__38_chanx_right_out[0] ,
    \sb_1__1__38_chanx_right_out[1] ,
    \sb_1__1__38_chanx_right_out[2] ,
    \sb_1__1__38_chanx_right_out[3] ,
    \sb_1__1__38_chanx_right_out[4] ,
    \sb_1__1__38_chanx_right_out[5] ,
    \sb_1__1__38_chanx_right_out[6] ,
    \sb_1__1__38_chanx_right_out[7] ,
    \sb_1__1__38_chanx_right_out[8] ,
    \sb_1__1__38_chanx_right_out[9] ,
    \sb_1__1__38_chanx_right_out[10] ,
    \sb_1__1__38_chanx_right_out[11] ,
    \sb_1__1__38_chanx_right_out[12] ,
    \sb_1__1__38_chanx_right_out[13] ,
    \sb_1__1__38_chanx_right_out[14] ,
    \sb_1__1__38_chanx_right_out[15] ,
    \sb_1__1__38_chanx_right_out[16] ,
    \sb_1__1__38_chanx_right_out[17] ,
    \sb_1__1__38_chanx_right_out[18] ,
    \sb_1__1__38_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__43_chany_top_out[0] ,
    \cby_1__1__43_chany_top_out[1] ,
    \cby_1__1__43_chany_top_out[2] ,
    \cby_1__1__43_chany_top_out[3] ,
    \cby_1__1__43_chany_top_out[4] ,
    \cby_1__1__43_chany_top_out[5] ,
    \cby_1__1__43_chany_top_out[6] ,
    \cby_1__1__43_chany_top_out[7] ,
    \cby_1__1__43_chany_top_out[8] ,
    \cby_1__1__43_chany_top_out[9] ,
    \cby_1__1__43_chany_top_out[10] ,
    \cby_1__1__43_chany_top_out[11] ,
    \cby_1__1__43_chany_top_out[12] ,
    \cby_1__1__43_chany_top_out[13] ,
    \cby_1__1__43_chany_top_out[14] ,
    \cby_1__1__43_chany_top_out[15] ,
    \cby_1__1__43_chany_top_out[16] ,
    \cby_1__1__43_chany_top_out[17] ,
    \cby_1__1__43_chany_top_out[18] ,
    \cby_1__1__43_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__38_chany_bottom_out[0] ,
    \sb_1__1__38_chany_bottom_out[1] ,
    \sb_1__1__38_chany_bottom_out[2] ,
    \sb_1__1__38_chany_bottom_out[3] ,
    \sb_1__1__38_chany_bottom_out[4] ,
    \sb_1__1__38_chany_bottom_out[5] ,
    \sb_1__1__38_chany_bottom_out[6] ,
    \sb_1__1__38_chany_bottom_out[7] ,
    \sb_1__1__38_chany_bottom_out[8] ,
    \sb_1__1__38_chany_bottom_out[9] ,
    \sb_1__1__38_chany_bottom_out[10] ,
    \sb_1__1__38_chany_bottom_out[11] ,
    \sb_1__1__38_chany_bottom_out[12] ,
    \sb_1__1__38_chany_bottom_out[13] ,
    \sb_1__1__38_chany_bottom_out[14] ,
    \sb_1__1__38_chany_bottom_out[15] ,
    \sb_1__1__38_chany_bottom_out[16] ,
    \sb_1__1__38_chany_bottom_out[17] ,
    \sb_1__1__38_chany_bottom_out[18] ,
    \sb_1__1__38_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__44_chany_bottom_out[0] ,
    \cby_1__1__44_chany_bottom_out[1] ,
    \cby_1__1__44_chany_bottom_out[2] ,
    \cby_1__1__44_chany_bottom_out[3] ,
    \cby_1__1__44_chany_bottom_out[4] ,
    \cby_1__1__44_chany_bottom_out[5] ,
    \cby_1__1__44_chany_bottom_out[6] ,
    \cby_1__1__44_chany_bottom_out[7] ,
    \cby_1__1__44_chany_bottom_out[8] ,
    \cby_1__1__44_chany_bottom_out[9] ,
    \cby_1__1__44_chany_bottom_out[10] ,
    \cby_1__1__44_chany_bottom_out[11] ,
    \cby_1__1__44_chany_bottom_out[12] ,
    \cby_1__1__44_chany_bottom_out[13] ,
    \cby_1__1__44_chany_bottom_out[14] ,
    \cby_1__1__44_chany_bottom_out[15] ,
    \cby_1__1__44_chany_bottom_out[16] ,
    \cby_1__1__44_chany_bottom_out[17] ,
    \cby_1__1__44_chany_bottom_out[18] ,
    \cby_1__1__44_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__38_chany_top_out[0] ,
    \sb_1__1__38_chany_top_out[1] ,
    \sb_1__1__38_chany_top_out[2] ,
    \sb_1__1__38_chany_top_out[3] ,
    \sb_1__1__38_chany_top_out[4] ,
    \sb_1__1__38_chany_top_out[5] ,
    \sb_1__1__38_chany_top_out[6] ,
    \sb_1__1__38_chany_top_out[7] ,
    \sb_1__1__38_chany_top_out[8] ,
    \sb_1__1__38_chany_top_out[9] ,
    \sb_1__1__38_chany_top_out[10] ,
    \sb_1__1__38_chany_top_out[11] ,
    \sb_1__1__38_chany_top_out[12] ,
    \sb_1__1__38_chany_top_out[13] ,
    \sb_1__1__38_chany_top_out[14] ,
    \sb_1__1__38_chany_top_out[15] ,
    \sb_1__1__38_chany_top_out[16] ,
    \sb_1__1__38_chany_top_out[17] ,
    \sb_1__1__38_chany_top_out[18] ,
    \sb_1__1__38_chany_top_out[19] }));
 sb_1__1_ sb_6__5_ (.bottom_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__46_ccff_tail),
    .ccff_tail(sb_1__1__39_ccff_tail),
    .clk_3_N_in(\clk_3_wires[19] ),
    .clk_3_N_out(\clk_3_wires[22] ),
    .left_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[164] ),
    .prog_clk_3_N_in(\prog_clk_3_wires[19] ),
    .prog_clk_3_N_out(\prog_clk_3_wires[22] ),
    .right_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__39_chanx_right_out[0] ,
    \cbx_1__1__39_chanx_right_out[1] ,
    \cbx_1__1__39_chanx_right_out[2] ,
    \cbx_1__1__39_chanx_right_out[3] ,
    \cbx_1__1__39_chanx_right_out[4] ,
    \cbx_1__1__39_chanx_right_out[5] ,
    \cbx_1__1__39_chanx_right_out[6] ,
    \cbx_1__1__39_chanx_right_out[7] ,
    \cbx_1__1__39_chanx_right_out[8] ,
    \cbx_1__1__39_chanx_right_out[9] ,
    \cbx_1__1__39_chanx_right_out[10] ,
    \cbx_1__1__39_chanx_right_out[11] ,
    \cbx_1__1__39_chanx_right_out[12] ,
    \cbx_1__1__39_chanx_right_out[13] ,
    \cbx_1__1__39_chanx_right_out[14] ,
    \cbx_1__1__39_chanx_right_out[15] ,
    \cbx_1__1__39_chanx_right_out[16] ,
    \cbx_1__1__39_chanx_right_out[17] ,
    \cbx_1__1__39_chanx_right_out[18] ,
    \cbx_1__1__39_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__39_chanx_left_out[0] ,
    \sb_1__1__39_chanx_left_out[1] ,
    \sb_1__1__39_chanx_left_out[2] ,
    \sb_1__1__39_chanx_left_out[3] ,
    \sb_1__1__39_chanx_left_out[4] ,
    \sb_1__1__39_chanx_left_out[5] ,
    \sb_1__1__39_chanx_left_out[6] ,
    \sb_1__1__39_chanx_left_out[7] ,
    \sb_1__1__39_chanx_left_out[8] ,
    \sb_1__1__39_chanx_left_out[9] ,
    \sb_1__1__39_chanx_left_out[10] ,
    \sb_1__1__39_chanx_left_out[11] ,
    \sb_1__1__39_chanx_left_out[12] ,
    \sb_1__1__39_chanx_left_out[13] ,
    \sb_1__1__39_chanx_left_out[14] ,
    \sb_1__1__39_chanx_left_out[15] ,
    \sb_1__1__39_chanx_left_out[16] ,
    \sb_1__1__39_chanx_left_out[17] ,
    \sb_1__1__39_chanx_left_out[18] ,
    \sb_1__1__39_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__46_chanx_left_out[0] ,
    \cbx_1__1__46_chanx_left_out[1] ,
    \cbx_1__1__46_chanx_left_out[2] ,
    \cbx_1__1__46_chanx_left_out[3] ,
    \cbx_1__1__46_chanx_left_out[4] ,
    \cbx_1__1__46_chanx_left_out[5] ,
    \cbx_1__1__46_chanx_left_out[6] ,
    \cbx_1__1__46_chanx_left_out[7] ,
    \cbx_1__1__46_chanx_left_out[8] ,
    \cbx_1__1__46_chanx_left_out[9] ,
    \cbx_1__1__46_chanx_left_out[10] ,
    \cbx_1__1__46_chanx_left_out[11] ,
    \cbx_1__1__46_chanx_left_out[12] ,
    \cbx_1__1__46_chanx_left_out[13] ,
    \cbx_1__1__46_chanx_left_out[14] ,
    \cbx_1__1__46_chanx_left_out[15] ,
    \cbx_1__1__46_chanx_left_out[16] ,
    \cbx_1__1__46_chanx_left_out[17] ,
    \cbx_1__1__46_chanx_left_out[18] ,
    \cbx_1__1__46_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__39_chanx_right_out[0] ,
    \sb_1__1__39_chanx_right_out[1] ,
    \sb_1__1__39_chanx_right_out[2] ,
    \sb_1__1__39_chanx_right_out[3] ,
    \sb_1__1__39_chanx_right_out[4] ,
    \sb_1__1__39_chanx_right_out[5] ,
    \sb_1__1__39_chanx_right_out[6] ,
    \sb_1__1__39_chanx_right_out[7] ,
    \sb_1__1__39_chanx_right_out[8] ,
    \sb_1__1__39_chanx_right_out[9] ,
    \sb_1__1__39_chanx_right_out[10] ,
    \sb_1__1__39_chanx_right_out[11] ,
    \sb_1__1__39_chanx_right_out[12] ,
    \sb_1__1__39_chanx_right_out[13] ,
    \sb_1__1__39_chanx_right_out[14] ,
    \sb_1__1__39_chanx_right_out[15] ,
    \sb_1__1__39_chanx_right_out[16] ,
    \sb_1__1__39_chanx_right_out[17] ,
    \sb_1__1__39_chanx_right_out[18] ,
    \sb_1__1__39_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__44_chany_top_out[0] ,
    \cby_1__1__44_chany_top_out[1] ,
    \cby_1__1__44_chany_top_out[2] ,
    \cby_1__1__44_chany_top_out[3] ,
    \cby_1__1__44_chany_top_out[4] ,
    \cby_1__1__44_chany_top_out[5] ,
    \cby_1__1__44_chany_top_out[6] ,
    \cby_1__1__44_chany_top_out[7] ,
    \cby_1__1__44_chany_top_out[8] ,
    \cby_1__1__44_chany_top_out[9] ,
    \cby_1__1__44_chany_top_out[10] ,
    \cby_1__1__44_chany_top_out[11] ,
    \cby_1__1__44_chany_top_out[12] ,
    \cby_1__1__44_chany_top_out[13] ,
    \cby_1__1__44_chany_top_out[14] ,
    \cby_1__1__44_chany_top_out[15] ,
    \cby_1__1__44_chany_top_out[16] ,
    \cby_1__1__44_chany_top_out[17] ,
    \cby_1__1__44_chany_top_out[18] ,
    \cby_1__1__44_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__39_chany_bottom_out[0] ,
    \sb_1__1__39_chany_bottom_out[1] ,
    \sb_1__1__39_chany_bottom_out[2] ,
    \sb_1__1__39_chany_bottom_out[3] ,
    \sb_1__1__39_chany_bottom_out[4] ,
    \sb_1__1__39_chany_bottom_out[5] ,
    \sb_1__1__39_chany_bottom_out[6] ,
    \sb_1__1__39_chany_bottom_out[7] ,
    \sb_1__1__39_chany_bottom_out[8] ,
    \sb_1__1__39_chany_bottom_out[9] ,
    \sb_1__1__39_chany_bottom_out[10] ,
    \sb_1__1__39_chany_bottom_out[11] ,
    \sb_1__1__39_chany_bottom_out[12] ,
    \sb_1__1__39_chany_bottom_out[13] ,
    \sb_1__1__39_chany_bottom_out[14] ,
    \sb_1__1__39_chany_bottom_out[15] ,
    \sb_1__1__39_chany_bottom_out[16] ,
    \sb_1__1__39_chany_bottom_out[17] ,
    \sb_1__1__39_chany_bottom_out[18] ,
    \sb_1__1__39_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__45_chany_bottom_out[0] ,
    \cby_1__1__45_chany_bottom_out[1] ,
    \cby_1__1__45_chany_bottom_out[2] ,
    \cby_1__1__45_chany_bottom_out[3] ,
    \cby_1__1__45_chany_bottom_out[4] ,
    \cby_1__1__45_chany_bottom_out[5] ,
    \cby_1__1__45_chany_bottom_out[6] ,
    \cby_1__1__45_chany_bottom_out[7] ,
    \cby_1__1__45_chany_bottom_out[8] ,
    \cby_1__1__45_chany_bottom_out[9] ,
    \cby_1__1__45_chany_bottom_out[10] ,
    \cby_1__1__45_chany_bottom_out[11] ,
    \cby_1__1__45_chany_bottom_out[12] ,
    \cby_1__1__45_chany_bottom_out[13] ,
    \cby_1__1__45_chany_bottom_out[14] ,
    \cby_1__1__45_chany_bottom_out[15] ,
    \cby_1__1__45_chany_bottom_out[16] ,
    \cby_1__1__45_chany_bottom_out[17] ,
    \cby_1__1__45_chany_bottom_out[18] ,
    \cby_1__1__45_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__39_chany_top_out[0] ,
    \sb_1__1__39_chany_top_out[1] ,
    \sb_1__1__39_chany_top_out[2] ,
    \sb_1__1__39_chany_top_out[3] ,
    \sb_1__1__39_chany_top_out[4] ,
    \sb_1__1__39_chany_top_out[5] ,
    \sb_1__1__39_chany_top_out[6] ,
    \sb_1__1__39_chany_top_out[7] ,
    \sb_1__1__39_chany_top_out[8] ,
    \sb_1__1__39_chany_top_out[9] ,
    \sb_1__1__39_chany_top_out[10] ,
    \sb_1__1__39_chany_top_out[11] ,
    \sb_1__1__39_chany_top_out[12] ,
    \sb_1__1__39_chany_top_out[13] ,
    \sb_1__1__39_chany_top_out[14] ,
    \sb_1__1__39_chany_top_out[15] ,
    \sb_1__1__39_chany_top_out[16] ,
    \sb_1__1__39_chany_top_out[17] ,
    \sb_1__1__39_chany_top_out[18] ,
    \sb_1__1__39_chany_top_out[19] }));
 sb_1__1_ sb_6__6_ (.bottom_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__47_ccff_tail),
    .ccff_tail(sb_1__1__40_ccff_tail),
    .clk_2_E_out(\clk_2_wires[40] ),
    .clk_2_N_in(\clk_3_wires[23] ),
    .clk_2_W_out(\clk_2_wires[42] ),
    .left_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[167] ),
    .prog_clk_2_E_out(\prog_clk_2_wires[40] ),
    .prog_clk_2_N_in(\prog_clk_3_wires[23] ),
    .prog_clk_2_W_out(\prog_clk_2_wires[42] ),
    .right_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__40_chanx_right_out[0] ,
    \cbx_1__1__40_chanx_right_out[1] ,
    \cbx_1__1__40_chanx_right_out[2] ,
    \cbx_1__1__40_chanx_right_out[3] ,
    \cbx_1__1__40_chanx_right_out[4] ,
    \cbx_1__1__40_chanx_right_out[5] ,
    \cbx_1__1__40_chanx_right_out[6] ,
    \cbx_1__1__40_chanx_right_out[7] ,
    \cbx_1__1__40_chanx_right_out[8] ,
    \cbx_1__1__40_chanx_right_out[9] ,
    \cbx_1__1__40_chanx_right_out[10] ,
    \cbx_1__1__40_chanx_right_out[11] ,
    \cbx_1__1__40_chanx_right_out[12] ,
    \cbx_1__1__40_chanx_right_out[13] ,
    \cbx_1__1__40_chanx_right_out[14] ,
    \cbx_1__1__40_chanx_right_out[15] ,
    \cbx_1__1__40_chanx_right_out[16] ,
    \cbx_1__1__40_chanx_right_out[17] ,
    \cbx_1__1__40_chanx_right_out[18] ,
    \cbx_1__1__40_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__40_chanx_left_out[0] ,
    \sb_1__1__40_chanx_left_out[1] ,
    \sb_1__1__40_chanx_left_out[2] ,
    \sb_1__1__40_chanx_left_out[3] ,
    \sb_1__1__40_chanx_left_out[4] ,
    \sb_1__1__40_chanx_left_out[5] ,
    \sb_1__1__40_chanx_left_out[6] ,
    \sb_1__1__40_chanx_left_out[7] ,
    \sb_1__1__40_chanx_left_out[8] ,
    \sb_1__1__40_chanx_left_out[9] ,
    \sb_1__1__40_chanx_left_out[10] ,
    \sb_1__1__40_chanx_left_out[11] ,
    \sb_1__1__40_chanx_left_out[12] ,
    \sb_1__1__40_chanx_left_out[13] ,
    \sb_1__1__40_chanx_left_out[14] ,
    \sb_1__1__40_chanx_left_out[15] ,
    \sb_1__1__40_chanx_left_out[16] ,
    \sb_1__1__40_chanx_left_out[17] ,
    \sb_1__1__40_chanx_left_out[18] ,
    \sb_1__1__40_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__47_chanx_left_out[0] ,
    \cbx_1__1__47_chanx_left_out[1] ,
    \cbx_1__1__47_chanx_left_out[2] ,
    \cbx_1__1__47_chanx_left_out[3] ,
    \cbx_1__1__47_chanx_left_out[4] ,
    \cbx_1__1__47_chanx_left_out[5] ,
    \cbx_1__1__47_chanx_left_out[6] ,
    \cbx_1__1__47_chanx_left_out[7] ,
    \cbx_1__1__47_chanx_left_out[8] ,
    \cbx_1__1__47_chanx_left_out[9] ,
    \cbx_1__1__47_chanx_left_out[10] ,
    \cbx_1__1__47_chanx_left_out[11] ,
    \cbx_1__1__47_chanx_left_out[12] ,
    \cbx_1__1__47_chanx_left_out[13] ,
    \cbx_1__1__47_chanx_left_out[14] ,
    \cbx_1__1__47_chanx_left_out[15] ,
    \cbx_1__1__47_chanx_left_out[16] ,
    \cbx_1__1__47_chanx_left_out[17] ,
    \cbx_1__1__47_chanx_left_out[18] ,
    \cbx_1__1__47_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__40_chanx_right_out[0] ,
    \sb_1__1__40_chanx_right_out[1] ,
    \sb_1__1__40_chanx_right_out[2] ,
    \sb_1__1__40_chanx_right_out[3] ,
    \sb_1__1__40_chanx_right_out[4] ,
    \sb_1__1__40_chanx_right_out[5] ,
    \sb_1__1__40_chanx_right_out[6] ,
    \sb_1__1__40_chanx_right_out[7] ,
    \sb_1__1__40_chanx_right_out[8] ,
    \sb_1__1__40_chanx_right_out[9] ,
    \sb_1__1__40_chanx_right_out[10] ,
    \sb_1__1__40_chanx_right_out[11] ,
    \sb_1__1__40_chanx_right_out[12] ,
    \sb_1__1__40_chanx_right_out[13] ,
    \sb_1__1__40_chanx_right_out[14] ,
    \sb_1__1__40_chanx_right_out[15] ,
    \sb_1__1__40_chanx_right_out[16] ,
    \sb_1__1__40_chanx_right_out[17] ,
    \sb_1__1__40_chanx_right_out[18] ,
    \sb_1__1__40_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__45_chany_top_out[0] ,
    \cby_1__1__45_chany_top_out[1] ,
    \cby_1__1__45_chany_top_out[2] ,
    \cby_1__1__45_chany_top_out[3] ,
    \cby_1__1__45_chany_top_out[4] ,
    \cby_1__1__45_chany_top_out[5] ,
    \cby_1__1__45_chany_top_out[6] ,
    \cby_1__1__45_chany_top_out[7] ,
    \cby_1__1__45_chany_top_out[8] ,
    \cby_1__1__45_chany_top_out[9] ,
    \cby_1__1__45_chany_top_out[10] ,
    \cby_1__1__45_chany_top_out[11] ,
    \cby_1__1__45_chany_top_out[12] ,
    \cby_1__1__45_chany_top_out[13] ,
    \cby_1__1__45_chany_top_out[14] ,
    \cby_1__1__45_chany_top_out[15] ,
    \cby_1__1__45_chany_top_out[16] ,
    \cby_1__1__45_chany_top_out[17] ,
    \cby_1__1__45_chany_top_out[18] ,
    \cby_1__1__45_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__40_chany_bottom_out[0] ,
    \sb_1__1__40_chany_bottom_out[1] ,
    \sb_1__1__40_chany_bottom_out[2] ,
    \sb_1__1__40_chany_bottom_out[3] ,
    \sb_1__1__40_chany_bottom_out[4] ,
    \sb_1__1__40_chany_bottom_out[5] ,
    \sb_1__1__40_chany_bottom_out[6] ,
    \sb_1__1__40_chany_bottom_out[7] ,
    \sb_1__1__40_chany_bottom_out[8] ,
    \sb_1__1__40_chany_bottom_out[9] ,
    \sb_1__1__40_chany_bottom_out[10] ,
    \sb_1__1__40_chany_bottom_out[11] ,
    \sb_1__1__40_chany_bottom_out[12] ,
    \sb_1__1__40_chany_bottom_out[13] ,
    \sb_1__1__40_chany_bottom_out[14] ,
    \sb_1__1__40_chany_bottom_out[15] ,
    \sb_1__1__40_chany_bottom_out[16] ,
    \sb_1__1__40_chany_bottom_out[17] ,
    \sb_1__1__40_chany_bottom_out[18] ,
    \sb_1__1__40_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__46_chany_bottom_out[0] ,
    \cby_1__1__46_chany_bottom_out[1] ,
    \cby_1__1__46_chany_bottom_out[2] ,
    \cby_1__1__46_chany_bottom_out[3] ,
    \cby_1__1__46_chany_bottom_out[4] ,
    \cby_1__1__46_chany_bottom_out[5] ,
    \cby_1__1__46_chany_bottom_out[6] ,
    \cby_1__1__46_chany_bottom_out[7] ,
    \cby_1__1__46_chany_bottom_out[8] ,
    \cby_1__1__46_chany_bottom_out[9] ,
    \cby_1__1__46_chany_bottom_out[10] ,
    \cby_1__1__46_chany_bottom_out[11] ,
    \cby_1__1__46_chany_bottom_out[12] ,
    \cby_1__1__46_chany_bottom_out[13] ,
    \cby_1__1__46_chany_bottom_out[14] ,
    \cby_1__1__46_chany_bottom_out[15] ,
    \cby_1__1__46_chany_bottom_out[16] ,
    \cby_1__1__46_chany_bottom_out[17] ,
    \cby_1__1__46_chany_bottom_out[18] ,
    \cby_1__1__46_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__40_chany_top_out[0] ,
    \sb_1__1__40_chany_top_out[1] ,
    \sb_1__1__40_chany_top_out[2] ,
    \sb_1__1__40_chany_top_out[3] ,
    \sb_1__1__40_chany_top_out[4] ,
    \sb_1__1__40_chany_top_out[5] ,
    \sb_1__1__40_chany_top_out[6] ,
    \sb_1__1__40_chany_top_out[7] ,
    \sb_1__1__40_chany_top_out[8] ,
    \sb_1__1__40_chany_top_out[9] ,
    \sb_1__1__40_chany_top_out[10] ,
    \sb_1__1__40_chany_top_out[11] ,
    \sb_1__1__40_chany_top_out[12] ,
    \sb_1__1__40_chany_top_out[13] ,
    \sb_1__1__40_chany_top_out[14] ,
    \sb_1__1__40_chany_top_out[15] ,
    \sb_1__1__40_chany_top_out[16] ,
    \sb_1__1__40_chany_top_out[17] ,
    \sb_1__1__40_chany_top_out[18] ,
    \sb_1__1__40_chany_top_out[19] }));
 sb_1__1_ sb_6__7_ (.bottom_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__48_ccff_tail),
    .ccff_tail(sb_1__1__41_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[170] ),
    .right_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__41_chanx_right_out[0] ,
    \cbx_1__1__41_chanx_right_out[1] ,
    \cbx_1__1__41_chanx_right_out[2] ,
    \cbx_1__1__41_chanx_right_out[3] ,
    \cbx_1__1__41_chanx_right_out[4] ,
    \cbx_1__1__41_chanx_right_out[5] ,
    \cbx_1__1__41_chanx_right_out[6] ,
    \cbx_1__1__41_chanx_right_out[7] ,
    \cbx_1__1__41_chanx_right_out[8] ,
    \cbx_1__1__41_chanx_right_out[9] ,
    \cbx_1__1__41_chanx_right_out[10] ,
    \cbx_1__1__41_chanx_right_out[11] ,
    \cbx_1__1__41_chanx_right_out[12] ,
    \cbx_1__1__41_chanx_right_out[13] ,
    \cbx_1__1__41_chanx_right_out[14] ,
    \cbx_1__1__41_chanx_right_out[15] ,
    \cbx_1__1__41_chanx_right_out[16] ,
    \cbx_1__1__41_chanx_right_out[17] ,
    \cbx_1__1__41_chanx_right_out[18] ,
    \cbx_1__1__41_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__41_chanx_left_out[0] ,
    \sb_1__1__41_chanx_left_out[1] ,
    \sb_1__1__41_chanx_left_out[2] ,
    \sb_1__1__41_chanx_left_out[3] ,
    \sb_1__1__41_chanx_left_out[4] ,
    \sb_1__1__41_chanx_left_out[5] ,
    \sb_1__1__41_chanx_left_out[6] ,
    \sb_1__1__41_chanx_left_out[7] ,
    \sb_1__1__41_chanx_left_out[8] ,
    \sb_1__1__41_chanx_left_out[9] ,
    \sb_1__1__41_chanx_left_out[10] ,
    \sb_1__1__41_chanx_left_out[11] ,
    \sb_1__1__41_chanx_left_out[12] ,
    \sb_1__1__41_chanx_left_out[13] ,
    \sb_1__1__41_chanx_left_out[14] ,
    \sb_1__1__41_chanx_left_out[15] ,
    \sb_1__1__41_chanx_left_out[16] ,
    \sb_1__1__41_chanx_left_out[17] ,
    \sb_1__1__41_chanx_left_out[18] ,
    \sb_1__1__41_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__48_chanx_left_out[0] ,
    \cbx_1__1__48_chanx_left_out[1] ,
    \cbx_1__1__48_chanx_left_out[2] ,
    \cbx_1__1__48_chanx_left_out[3] ,
    \cbx_1__1__48_chanx_left_out[4] ,
    \cbx_1__1__48_chanx_left_out[5] ,
    \cbx_1__1__48_chanx_left_out[6] ,
    \cbx_1__1__48_chanx_left_out[7] ,
    \cbx_1__1__48_chanx_left_out[8] ,
    \cbx_1__1__48_chanx_left_out[9] ,
    \cbx_1__1__48_chanx_left_out[10] ,
    \cbx_1__1__48_chanx_left_out[11] ,
    \cbx_1__1__48_chanx_left_out[12] ,
    \cbx_1__1__48_chanx_left_out[13] ,
    \cbx_1__1__48_chanx_left_out[14] ,
    \cbx_1__1__48_chanx_left_out[15] ,
    \cbx_1__1__48_chanx_left_out[16] ,
    \cbx_1__1__48_chanx_left_out[17] ,
    \cbx_1__1__48_chanx_left_out[18] ,
    \cbx_1__1__48_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__41_chanx_right_out[0] ,
    \sb_1__1__41_chanx_right_out[1] ,
    \sb_1__1__41_chanx_right_out[2] ,
    \sb_1__1__41_chanx_right_out[3] ,
    \sb_1__1__41_chanx_right_out[4] ,
    \sb_1__1__41_chanx_right_out[5] ,
    \sb_1__1__41_chanx_right_out[6] ,
    \sb_1__1__41_chanx_right_out[7] ,
    \sb_1__1__41_chanx_right_out[8] ,
    \sb_1__1__41_chanx_right_out[9] ,
    \sb_1__1__41_chanx_right_out[10] ,
    \sb_1__1__41_chanx_right_out[11] ,
    \sb_1__1__41_chanx_right_out[12] ,
    \sb_1__1__41_chanx_right_out[13] ,
    \sb_1__1__41_chanx_right_out[14] ,
    \sb_1__1__41_chanx_right_out[15] ,
    \sb_1__1__41_chanx_right_out[16] ,
    \sb_1__1__41_chanx_right_out[17] ,
    \sb_1__1__41_chanx_right_out[18] ,
    \sb_1__1__41_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__46_chany_top_out[0] ,
    \cby_1__1__46_chany_top_out[1] ,
    \cby_1__1__46_chany_top_out[2] ,
    \cby_1__1__46_chany_top_out[3] ,
    \cby_1__1__46_chany_top_out[4] ,
    \cby_1__1__46_chany_top_out[5] ,
    \cby_1__1__46_chany_top_out[6] ,
    \cby_1__1__46_chany_top_out[7] ,
    \cby_1__1__46_chany_top_out[8] ,
    \cby_1__1__46_chany_top_out[9] ,
    \cby_1__1__46_chany_top_out[10] ,
    \cby_1__1__46_chany_top_out[11] ,
    \cby_1__1__46_chany_top_out[12] ,
    \cby_1__1__46_chany_top_out[13] ,
    \cby_1__1__46_chany_top_out[14] ,
    \cby_1__1__46_chany_top_out[15] ,
    \cby_1__1__46_chany_top_out[16] ,
    \cby_1__1__46_chany_top_out[17] ,
    \cby_1__1__46_chany_top_out[18] ,
    \cby_1__1__46_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__41_chany_bottom_out[0] ,
    \sb_1__1__41_chany_bottom_out[1] ,
    \sb_1__1__41_chany_bottom_out[2] ,
    \sb_1__1__41_chany_bottom_out[3] ,
    \sb_1__1__41_chany_bottom_out[4] ,
    \sb_1__1__41_chany_bottom_out[5] ,
    \sb_1__1__41_chany_bottom_out[6] ,
    \sb_1__1__41_chany_bottom_out[7] ,
    \sb_1__1__41_chany_bottom_out[8] ,
    \sb_1__1__41_chany_bottom_out[9] ,
    \sb_1__1__41_chany_bottom_out[10] ,
    \sb_1__1__41_chany_bottom_out[11] ,
    \sb_1__1__41_chany_bottom_out[12] ,
    \sb_1__1__41_chany_bottom_out[13] ,
    \sb_1__1__41_chany_bottom_out[14] ,
    \sb_1__1__41_chany_bottom_out[15] ,
    \sb_1__1__41_chany_bottom_out[16] ,
    \sb_1__1__41_chany_bottom_out[17] ,
    \sb_1__1__41_chany_bottom_out[18] ,
    \sb_1__1__41_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__47_chany_bottom_out[0] ,
    \cby_1__1__47_chany_bottom_out[1] ,
    \cby_1__1__47_chany_bottom_out[2] ,
    \cby_1__1__47_chany_bottom_out[3] ,
    \cby_1__1__47_chany_bottom_out[4] ,
    \cby_1__1__47_chany_bottom_out[5] ,
    \cby_1__1__47_chany_bottom_out[6] ,
    \cby_1__1__47_chany_bottom_out[7] ,
    \cby_1__1__47_chany_bottom_out[8] ,
    \cby_1__1__47_chany_bottom_out[9] ,
    \cby_1__1__47_chany_bottom_out[10] ,
    \cby_1__1__47_chany_bottom_out[11] ,
    \cby_1__1__47_chany_bottom_out[12] ,
    \cby_1__1__47_chany_bottom_out[13] ,
    \cby_1__1__47_chany_bottom_out[14] ,
    \cby_1__1__47_chany_bottom_out[15] ,
    \cby_1__1__47_chany_bottom_out[16] ,
    \cby_1__1__47_chany_bottom_out[17] ,
    \cby_1__1__47_chany_bottom_out[18] ,
    \cby_1__1__47_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__41_chany_top_out[0] ,
    \sb_1__1__41_chany_top_out[1] ,
    \sb_1__1__41_chany_top_out[2] ,
    \sb_1__1__41_chany_top_out[3] ,
    \sb_1__1__41_chany_top_out[4] ,
    \sb_1__1__41_chany_top_out[5] ,
    \sb_1__1__41_chany_top_out[6] ,
    \sb_1__1__41_chany_top_out[7] ,
    \sb_1__1__41_chany_top_out[8] ,
    \sb_1__1__41_chany_top_out[9] ,
    \sb_1__1__41_chany_top_out[10] ,
    \sb_1__1__41_chany_top_out[11] ,
    \sb_1__1__41_chany_top_out[12] ,
    \sb_1__1__41_chany_top_out[13] ,
    \sb_1__1__41_chany_top_out[14] ,
    \sb_1__1__41_chany_top_out[15] ,
    \sb_1__1__41_chany_top_out[16] ,
    \sb_1__1__41_chany_top_out[17] ,
    \sb_1__1__41_chany_top_out[18] ,
    \sb_1__1__41_chany_top_out[19] }));
 sb_1__2_ sb_6__8_ (.SC_IN_BOT(\scff_Wires[110] ),
    .SC_OUT_BOT(\scff_Wires[111] ),
    .bottom_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_upper),
    .ccff_head(grid_io_top_6_ccff_tail),
    .ccff_tail(sb_1__8__5_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[172] ),
    .right_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__5_chanx_right_out[0] ,
    \cbx_1__8__5_chanx_right_out[1] ,
    \cbx_1__8__5_chanx_right_out[2] ,
    \cbx_1__8__5_chanx_right_out[3] ,
    \cbx_1__8__5_chanx_right_out[4] ,
    \cbx_1__8__5_chanx_right_out[5] ,
    \cbx_1__8__5_chanx_right_out[6] ,
    \cbx_1__8__5_chanx_right_out[7] ,
    \cbx_1__8__5_chanx_right_out[8] ,
    \cbx_1__8__5_chanx_right_out[9] ,
    \cbx_1__8__5_chanx_right_out[10] ,
    \cbx_1__8__5_chanx_right_out[11] ,
    \cbx_1__8__5_chanx_right_out[12] ,
    \cbx_1__8__5_chanx_right_out[13] ,
    \cbx_1__8__5_chanx_right_out[14] ,
    \cbx_1__8__5_chanx_right_out[15] ,
    \cbx_1__8__5_chanx_right_out[16] ,
    \cbx_1__8__5_chanx_right_out[17] ,
    \cbx_1__8__5_chanx_right_out[18] ,
    \cbx_1__8__5_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__8__5_chanx_left_out[0] ,
    \sb_1__8__5_chanx_left_out[1] ,
    \sb_1__8__5_chanx_left_out[2] ,
    \sb_1__8__5_chanx_left_out[3] ,
    \sb_1__8__5_chanx_left_out[4] ,
    \sb_1__8__5_chanx_left_out[5] ,
    \sb_1__8__5_chanx_left_out[6] ,
    \sb_1__8__5_chanx_left_out[7] ,
    \sb_1__8__5_chanx_left_out[8] ,
    \sb_1__8__5_chanx_left_out[9] ,
    \sb_1__8__5_chanx_left_out[10] ,
    \sb_1__8__5_chanx_left_out[11] ,
    \sb_1__8__5_chanx_left_out[12] ,
    \sb_1__8__5_chanx_left_out[13] ,
    \sb_1__8__5_chanx_left_out[14] ,
    \sb_1__8__5_chanx_left_out[15] ,
    \sb_1__8__5_chanx_left_out[16] ,
    \sb_1__8__5_chanx_left_out[17] ,
    \sb_1__8__5_chanx_left_out[18] ,
    \sb_1__8__5_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__8__6_chanx_left_out[0] ,
    \cbx_1__8__6_chanx_left_out[1] ,
    \cbx_1__8__6_chanx_left_out[2] ,
    \cbx_1__8__6_chanx_left_out[3] ,
    \cbx_1__8__6_chanx_left_out[4] ,
    \cbx_1__8__6_chanx_left_out[5] ,
    \cbx_1__8__6_chanx_left_out[6] ,
    \cbx_1__8__6_chanx_left_out[7] ,
    \cbx_1__8__6_chanx_left_out[8] ,
    \cbx_1__8__6_chanx_left_out[9] ,
    \cbx_1__8__6_chanx_left_out[10] ,
    \cbx_1__8__6_chanx_left_out[11] ,
    \cbx_1__8__6_chanx_left_out[12] ,
    \cbx_1__8__6_chanx_left_out[13] ,
    \cbx_1__8__6_chanx_left_out[14] ,
    \cbx_1__8__6_chanx_left_out[15] ,
    \cbx_1__8__6_chanx_left_out[16] ,
    \cbx_1__8__6_chanx_left_out[17] ,
    \cbx_1__8__6_chanx_left_out[18] ,
    \cbx_1__8__6_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__8__5_chanx_right_out[0] ,
    \sb_1__8__5_chanx_right_out[1] ,
    \sb_1__8__5_chanx_right_out[2] ,
    \sb_1__8__5_chanx_right_out[3] ,
    \sb_1__8__5_chanx_right_out[4] ,
    \sb_1__8__5_chanx_right_out[5] ,
    \sb_1__8__5_chanx_right_out[6] ,
    \sb_1__8__5_chanx_right_out[7] ,
    \sb_1__8__5_chanx_right_out[8] ,
    \sb_1__8__5_chanx_right_out[9] ,
    \sb_1__8__5_chanx_right_out[10] ,
    \sb_1__8__5_chanx_right_out[11] ,
    \sb_1__8__5_chanx_right_out[12] ,
    \sb_1__8__5_chanx_right_out[13] ,
    \sb_1__8__5_chanx_right_out[14] ,
    \sb_1__8__5_chanx_right_out[15] ,
    \sb_1__8__5_chanx_right_out[16] ,
    \sb_1__8__5_chanx_right_out[17] ,
    \sb_1__8__5_chanx_right_out[18] ,
    \sb_1__8__5_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__47_chany_top_out[0] ,
    \cby_1__1__47_chany_top_out[1] ,
    \cby_1__1__47_chany_top_out[2] ,
    \cby_1__1__47_chany_top_out[3] ,
    \cby_1__1__47_chany_top_out[4] ,
    \cby_1__1__47_chany_top_out[5] ,
    \cby_1__1__47_chany_top_out[6] ,
    \cby_1__1__47_chany_top_out[7] ,
    \cby_1__1__47_chany_top_out[8] ,
    \cby_1__1__47_chany_top_out[9] ,
    \cby_1__1__47_chany_top_out[10] ,
    \cby_1__1__47_chany_top_out[11] ,
    \cby_1__1__47_chany_top_out[12] ,
    \cby_1__1__47_chany_top_out[13] ,
    \cby_1__1__47_chany_top_out[14] ,
    \cby_1__1__47_chany_top_out[15] ,
    \cby_1__1__47_chany_top_out[16] ,
    \cby_1__1__47_chany_top_out[17] ,
    \cby_1__1__47_chany_top_out[18] ,
    \cby_1__1__47_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__8__5_chany_bottom_out[0] ,
    \sb_1__8__5_chany_bottom_out[1] ,
    \sb_1__8__5_chany_bottom_out[2] ,
    \sb_1__8__5_chany_bottom_out[3] ,
    \sb_1__8__5_chany_bottom_out[4] ,
    \sb_1__8__5_chany_bottom_out[5] ,
    \sb_1__8__5_chany_bottom_out[6] ,
    \sb_1__8__5_chany_bottom_out[7] ,
    \sb_1__8__5_chany_bottom_out[8] ,
    \sb_1__8__5_chany_bottom_out[9] ,
    \sb_1__8__5_chany_bottom_out[10] ,
    \sb_1__8__5_chany_bottom_out[11] ,
    \sb_1__8__5_chany_bottom_out[12] ,
    \sb_1__8__5_chany_bottom_out[13] ,
    \sb_1__8__5_chany_bottom_out[14] ,
    \sb_1__8__5_chany_bottom_out[15] ,
    \sb_1__8__5_chany_bottom_out[16] ,
    \sb_1__8__5_chany_bottom_out[17] ,
    \sb_1__8__5_chany_bottom_out[18] ,
    \sb_1__8__5_chany_bottom_out[19] }));
 sb_1__0_ sb_7__0_ (.SC_IN_TOP(\scff_Wires[129] ),
    .SC_OUT_TOP(\scff_Wires[130] ),
    .ccff_head(grid_io_bottom_0_ccff_tail),
    .ccff_tail(sb_1__0__6_ccff_tail),
    .left_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[175] ),
    .right_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_upper),
    .right_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_upper),
    .right_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_upper),
    .right_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_upper),
    .right_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_upper),
    .right_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_upper),
    .right_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_upper),
    .right_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_upper),
    .right_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_upper),
    .top_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__6_chanx_right_out[0] ,
    \cbx_1__0__6_chanx_right_out[1] ,
    \cbx_1__0__6_chanx_right_out[2] ,
    \cbx_1__0__6_chanx_right_out[3] ,
    \cbx_1__0__6_chanx_right_out[4] ,
    \cbx_1__0__6_chanx_right_out[5] ,
    \cbx_1__0__6_chanx_right_out[6] ,
    \cbx_1__0__6_chanx_right_out[7] ,
    \cbx_1__0__6_chanx_right_out[8] ,
    \cbx_1__0__6_chanx_right_out[9] ,
    \cbx_1__0__6_chanx_right_out[10] ,
    \cbx_1__0__6_chanx_right_out[11] ,
    \cbx_1__0__6_chanx_right_out[12] ,
    \cbx_1__0__6_chanx_right_out[13] ,
    \cbx_1__0__6_chanx_right_out[14] ,
    \cbx_1__0__6_chanx_right_out[15] ,
    \cbx_1__0__6_chanx_right_out[16] ,
    \cbx_1__0__6_chanx_right_out[17] ,
    \cbx_1__0__6_chanx_right_out[18] ,
    \cbx_1__0__6_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__0__6_chanx_left_out[0] ,
    \sb_1__0__6_chanx_left_out[1] ,
    \sb_1__0__6_chanx_left_out[2] ,
    \sb_1__0__6_chanx_left_out[3] ,
    \sb_1__0__6_chanx_left_out[4] ,
    \sb_1__0__6_chanx_left_out[5] ,
    \sb_1__0__6_chanx_left_out[6] ,
    \sb_1__0__6_chanx_left_out[7] ,
    \sb_1__0__6_chanx_left_out[8] ,
    \sb_1__0__6_chanx_left_out[9] ,
    \sb_1__0__6_chanx_left_out[10] ,
    \sb_1__0__6_chanx_left_out[11] ,
    \sb_1__0__6_chanx_left_out[12] ,
    \sb_1__0__6_chanx_left_out[13] ,
    \sb_1__0__6_chanx_left_out[14] ,
    \sb_1__0__6_chanx_left_out[15] ,
    \sb_1__0__6_chanx_left_out[16] ,
    \sb_1__0__6_chanx_left_out[17] ,
    \sb_1__0__6_chanx_left_out[18] ,
    \sb_1__0__6_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__0__7_chanx_left_out[0] ,
    \cbx_1__0__7_chanx_left_out[1] ,
    \cbx_1__0__7_chanx_left_out[2] ,
    \cbx_1__0__7_chanx_left_out[3] ,
    \cbx_1__0__7_chanx_left_out[4] ,
    \cbx_1__0__7_chanx_left_out[5] ,
    \cbx_1__0__7_chanx_left_out[6] ,
    \cbx_1__0__7_chanx_left_out[7] ,
    \cbx_1__0__7_chanx_left_out[8] ,
    \cbx_1__0__7_chanx_left_out[9] ,
    \cbx_1__0__7_chanx_left_out[10] ,
    \cbx_1__0__7_chanx_left_out[11] ,
    \cbx_1__0__7_chanx_left_out[12] ,
    \cbx_1__0__7_chanx_left_out[13] ,
    \cbx_1__0__7_chanx_left_out[14] ,
    \cbx_1__0__7_chanx_left_out[15] ,
    \cbx_1__0__7_chanx_left_out[16] ,
    \cbx_1__0__7_chanx_left_out[17] ,
    \cbx_1__0__7_chanx_left_out[18] ,
    \cbx_1__0__7_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__0__6_chanx_right_out[0] ,
    \sb_1__0__6_chanx_right_out[1] ,
    \sb_1__0__6_chanx_right_out[2] ,
    \sb_1__0__6_chanx_right_out[3] ,
    \sb_1__0__6_chanx_right_out[4] ,
    \sb_1__0__6_chanx_right_out[5] ,
    \sb_1__0__6_chanx_right_out[6] ,
    \sb_1__0__6_chanx_right_out[7] ,
    \sb_1__0__6_chanx_right_out[8] ,
    \sb_1__0__6_chanx_right_out[9] ,
    \sb_1__0__6_chanx_right_out[10] ,
    \sb_1__0__6_chanx_right_out[11] ,
    \sb_1__0__6_chanx_right_out[12] ,
    \sb_1__0__6_chanx_right_out[13] ,
    \sb_1__0__6_chanx_right_out[14] ,
    \sb_1__0__6_chanx_right_out[15] ,
    \sb_1__0__6_chanx_right_out[16] ,
    \sb_1__0__6_chanx_right_out[17] ,
    \sb_1__0__6_chanx_right_out[18] ,
    \sb_1__0__6_chanx_right_out[19] }),
    .chany_top_in({\cby_1__1__48_chany_bottom_out[0] ,
    \cby_1__1__48_chany_bottom_out[1] ,
    \cby_1__1__48_chany_bottom_out[2] ,
    \cby_1__1__48_chany_bottom_out[3] ,
    \cby_1__1__48_chany_bottom_out[4] ,
    \cby_1__1__48_chany_bottom_out[5] ,
    \cby_1__1__48_chany_bottom_out[6] ,
    \cby_1__1__48_chany_bottom_out[7] ,
    \cby_1__1__48_chany_bottom_out[8] ,
    \cby_1__1__48_chany_bottom_out[9] ,
    \cby_1__1__48_chany_bottom_out[10] ,
    \cby_1__1__48_chany_bottom_out[11] ,
    \cby_1__1__48_chany_bottom_out[12] ,
    \cby_1__1__48_chany_bottom_out[13] ,
    \cby_1__1__48_chany_bottom_out[14] ,
    \cby_1__1__48_chany_bottom_out[15] ,
    \cby_1__1__48_chany_bottom_out[16] ,
    \cby_1__1__48_chany_bottom_out[17] ,
    \cby_1__1__48_chany_bottom_out[18] ,
    \cby_1__1__48_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__0__6_chany_top_out[0] ,
    \sb_1__0__6_chany_top_out[1] ,
    \sb_1__0__6_chany_top_out[2] ,
    \sb_1__0__6_chany_top_out[3] ,
    \sb_1__0__6_chany_top_out[4] ,
    \sb_1__0__6_chany_top_out[5] ,
    \sb_1__0__6_chany_top_out[6] ,
    \sb_1__0__6_chany_top_out[7] ,
    \sb_1__0__6_chany_top_out[8] ,
    \sb_1__0__6_chany_top_out[9] ,
    \sb_1__0__6_chany_top_out[10] ,
    \sb_1__0__6_chany_top_out[11] ,
    \sb_1__0__6_chany_top_out[12] ,
    \sb_1__0__6_chany_top_out[13] ,
    \sb_1__0__6_chany_top_out[14] ,
    \sb_1__0__6_chany_top_out[15] ,
    \sb_1__0__6_chany_top_out[16] ,
    \sb_1__0__6_chany_top_out[17] ,
    \sb_1__0__6_chany_top_out[18] ,
    \sb_1__0__6_chany_top_out[19] }));
 sb_1__1_ sb_7__1_ (.bottom_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__49_ccff_tail),
    .ccff_tail(sb_1__1__42_ccff_tail),
    .clk_1_E_out(\clk_1_wires[85] ),
    .clk_1_N_in(\clk_2_wires[38] ),
    .clk_1_W_out(\clk_1_wires[86] ),
    .left_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[178] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[85] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[38] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[86] ),
    .right_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__42_chanx_right_out[0] ,
    \cbx_1__1__42_chanx_right_out[1] ,
    \cbx_1__1__42_chanx_right_out[2] ,
    \cbx_1__1__42_chanx_right_out[3] ,
    \cbx_1__1__42_chanx_right_out[4] ,
    \cbx_1__1__42_chanx_right_out[5] ,
    \cbx_1__1__42_chanx_right_out[6] ,
    \cbx_1__1__42_chanx_right_out[7] ,
    \cbx_1__1__42_chanx_right_out[8] ,
    \cbx_1__1__42_chanx_right_out[9] ,
    \cbx_1__1__42_chanx_right_out[10] ,
    \cbx_1__1__42_chanx_right_out[11] ,
    \cbx_1__1__42_chanx_right_out[12] ,
    \cbx_1__1__42_chanx_right_out[13] ,
    \cbx_1__1__42_chanx_right_out[14] ,
    \cbx_1__1__42_chanx_right_out[15] ,
    \cbx_1__1__42_chanx_right_out[16] ,
    \cbx_1__1__42_chanx_right_out[17] ,
    \cbx_1__1__42_chanx_right_out[18] ,
    \cbx_1__1__42_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__42_chanx_left_out[0] ,
    \sb_1__1__42_chanx_left_out[1] ,
    \sb_1__1__42_chanx_left_out[2] ,
    \sb_1__1__42_chanx_left_out[3] ,
    \sb_1__1__42_chanx_left_out[4] ,
    \sb_1__1__42_chanx_left_out[5] ,
    \sb_1__1__42_chanx_left_out[6] ,
    \sb_1__1__42_chanx_left_out[7] ,
    \sb_1__1__42_chanx_left_out[8] ,
    \sb_1__1__42_chanx_left_out[9] ,
    \sb_1__1__42_chanx_left_out[10] ,
    \sb_1__1__42_chanx_left_out[11] ,
    \sb_1__1__42_chanx_left_out[12] ,
    \sb_1__1__42_chanx_left_out[13] ,
    \sb_1__1__42_chanx_left_out[14] ,
    \sb_1__1__42_chanx_left_out[15] ,
    \sb_1__1__42_chanx_left_out[16] ,
    \sb_1__1__42_chanx_left_out[17] ,
    \sb_1__1__42_chanx_left_out[18] ,
    \sb_1__1__42_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__49_chanx_left_out[0] ,
    \cbx_1__1__49_chanx_left_out[1] ,
    \cbx_1__1__49_chanx_left_out[2] ,
    \cbx_1__1__49_chanx_left_out[3] ,
    \cbx_1__1__49_chanx_left_out[4] ,
    \cbx_1__1__49_chanx_left_out[5] ,
    \cbx_1__1__49_chanx_left_out[6] ,
    \cbx_1__1__49_chanx_left_out[7] ,
    \cbx_1__1__49_chanx_left_out[8] ,
    \cbx_1__1__49_chanx_left_out[9] ,
    \cbx_1__1__49_chanx_left_out[10] ,
    \cbx_1__1__49_chanx_left_out[11] ,
    \cbx_1__1__49_chanx_left_out[12] ,
    \cbx_1__1__49_chanx_left_out[13] ,
    \cbx_1__1__49_chanx_left_out[14] ,
    \cbx_1__1__49_chanx_left_out[15] ,
    \cbx_1__1__49_chanx_left_out[16] ,
    \cbx_1__1__49_chanx_left_out[17] ,
    \cbx_1__1__49_chanx_left_out[18] ,
    \cbx_1__1__49_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__42_chanx_right_out[0] ,
    \sb_1__1__42_chanx_right_out[1] ,
    \sb_1__1__42_chanx_right_out[2] ,
    \sb_1__1__42_chanx_right_out[3] ,
    \sb_1__1__42_chanx_right_out[4] ,
    \sb_1__1__42_chanx_right_out[5] ,
    \sb_1__1__42_chanx_right_out[6] ,
    \sb_1__1__42_chanx_right_out[7] ,
    \sb_1__1__42_chanx_right_out[8] ,
    \sb_1__1__42_chanx_right_out[9] ,
    \sb_1__1__42_chanx_right_out[10] ,
    \sb_1__1__42_chanx_right_out[11] ,
    \sb_1__1__42_chanx_right_out[12] ,
    \sb_1__1__42_chanx_right_out[13] ,
    \sb_1__1__42_chanx_right_out[14] ,
    \sb_1__1__42_chanx_right_out[15] ,
    \sb_1__1__42_chanx_right_out[16] ,
    \sb_1__1__42_chanx_right_out[17] ,
    \sb_1__1__42_chanx_right_out[18] ,
    \sb_1__1__42_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__48_chany_top_out[0] ,
    \cby_1__1__48_chany_top_out[1] ,
    \cby_1__1__48_chany_top_out[2] ,
    \cby_1__1__48_chany_top_out[3] ,
    \cby_1__1__48_chany_top_out[4] ,
    \cby_1__1__48_chany_top_out[5] ,
    \cby_1__1__48_chany_top_out[6] ,
    \cby_1__1__48_chany_top_out[7] ,
    \cby_1__1__48_chany_top_out[8] ,
    \cby_1__1__48_chany_top_out[9] ,
    \cby_1__1__48_chany_top_out[10] ,
    \cby_1__1__48_chany_top_out[11] ,
    \cby_1__1__48_chany_top_out[12] ,
    \cby_1__1__48_chany_top_out[13] ,
    \cby_1__1__48_chany_top_out[14] ,
    \cby_1__1__48_chany_top_out[15] ,
    \cby_1__1__48_chany_top_out[16] ,
    \cby_1__1__48_chany_top_out[17] ,
    \cby_1__1__48_chany_top_out[18] ,
    \cby_1__1__48_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__42_chany_bottom_out[0] ,
    \sb_1__1__42_chany_bottom_out[1] ,
    \sb_1__1__42_chany_bottom_out[2] ,
    \sb_1__1__42_chany_bottom_out[3] ,
    \sb_1__1__42_chany_bottom_out[4] ,
    \sb_1__1__42_chany_bottom_out[5] ,
    \sb_1__1__42_chany_bottom_out[6] ,
    \sb_1__1__42_chany_bottom_out[7] ,
    \sb_1__1__42_chany_bottom_out[8] ,
    \sb_1__1__42_chany_bottom_out[9] ,
    \sb_1__1__42_chany_bottom_out[10] ,
    \sb_1__1__42_chany_bottom_out[11] ,
    \sb_1__1__42_chany_bottom_out[12] ,
    \sb_1__1__42_chany_bottom_out[13] ,
    \sb_1__1__42_chany_bottom_out[14] ,
    \sb_1__1__42_chany_bottom_out[15] ,
    \sb_1__1__42_chany_bottom_out[16] ,
    \sb_1__1__42_chany_bottom_out[17] ,
    \sb_1__1__42_chany_bottom_out[18] ,
    \sb_1__1__42_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__49_chany_bottom_out[0] ,
    \cby_1__1__49_chany_bottom_out[1] ,
    \cby_1__1__49_chany_bottom_out[2] ,
    \cby_1__1__49_chany_bottom_out[3] ,
    \cby_1__1__49_chany_bottom_out[4] ,
    \cby_1__1__49_chany_bottom_out[5] ,
    \cby_1__1__49_chany_bottom_out[6] ,
    \cby_1__1__49_chany_bottom_out[7] ,
    \cby_1__1__49_chany_bottom_out[8] ,
    \cby_1__1__49_chany_bottom_out[9] ,
    \cby_1__1__49_chany_bottom_out[10] ,
    \cby_1__1__49_chany_bottom_out[11] ,
    \cby_1__1__49_chany_bottom_out[12] ,
    \cby_1__1__49_chany_bottom_out[13] ,
    \cby_1__1__49_chany_bottom_out[14] ,
    \cby_1__1__49_chany_bottom_out[15] ,
    \cby_1__1__49_chany_bottom_out[16] ,
    \cby_1__1__49_chany_bottom_out[17] ,
    \cby_1__1__49_chany_bottom_out[18] ,
    \cby_1__1__49_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__42_chany_top_out[0] ,
    \sb_1__1__42_chany_top_out[1] ,
    \sb_1__1__42_chany_top_out[2] ,
    \sb_1__1__42_chany_top_out[3] ,
    \sb_1__1__42_chany_top_out[4] ,
    \sb_1__1__42_chany_top_out[5] ,
    \sb_1__1__42_chany_top_out[6] ,
    \sb_1__1__42_chany_top_out[7] ,
    \sb_1__1__42_chany_top_out[8] ,
    \sb_1__1__42_chany_top_out[9] ,
    \sb_1__1__42_chany_top_out[10] ,
    \sb_1__1__42_chany_top_out[11] ,
    \sb_1__1__42_chany_top_out[12] ,
    \sb_1__1__42_chany_top_out[13] ,
    \sb_1__1__42_chany_top_out[14] ,
    \sb_1__1__42_chany_top_out[15] ,
    \sb_1__1__42_chany_top_out[16] ,
    \sb_1__1__42_chany_top_out[17] ,
    \sb_1__1__42_chany_top_out[18] ,
    \sb_1__1__42_chany_top_out[19] }));
 sb_1__1_ sb_7__2_ (.bottom_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__50_ccff_tail),
    .ccff_tail(sb_1__1__43_ccff_tail),
    .clk_2_N_in(\clk_2_wires[28] ),
    .clk_2_N_out(\clk_2_wires[35] ),
    .clk_2_S_out(\clk_2_wires[37] ),
    .left_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[181] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[28] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[35] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[37] ),
    .right_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__43_chanx_right_out[0] ,
    \cbx_1__1__43_chanx_right_out[1] ,
    \cbx_1__1__43_chanx_right_out[2] ,
    \cbx_1__1__43_chanx_right_out[3] ,
    \cbx_1__1__43_chanx_right_out[4] ,
    \cbx_1__1__43_chanx_right_out[5] ,
    \cbx_1__1__43_chanx_right_out[6] ,
    \cbx_1__1__43_chanx_right_out[7] ,
    \cbx_1__1__43_chanx_right_out[8] ,
    \cbx_1__1__43_chanx_right_out[9] ,
    \cbx_1__1__43_chanx_right_out[10] ,
    \cbx_1__1__43_chanx_right_out[11] ,
    \cbx_1__1__43_chanx_right_out[12] ,
    \cbx_1__1__43_chanx_right_out[13] ,
    \cbx_1__1__43_chanx_right_out[14] ,
    \cbx_1__1__43_chanx_right_out[15] ,
    \cbx_1__1__43_chanx_right_out[16] ,
    \cbx_1__1__43_chanx_right_out[17] ,
    \cbx_1__1__43_chanx_right_out[18] ,
    \cbx_1__1__43_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__43_chanx_left_out[0] ,
    \sb_1__1__43_chanx_left_out[1] ,
    \sb_1__1__43_chanx_left_out[2] ,
    \sb_1__1__43_chanx_left_out[3] ,
    \sb_1__1__43_chanx_left_out[4] ,
    \sb_1__1__43_chanx_left_out[5] ,
    \sb_1__1__43_chanx_left_out[6] ,
    \sb_1__1__43_chanx_left_out[7] ,
    \sb_1__1__43_chanx_left_out[8] ,
    \sb_1__1__43_chanx_left_out[9] ,
    \sb_1__1__43_chanx_left_out[10] ,
    \sb_1__1__43_chanx_left_out[11] ,
    \sb_1__1__43_chanx_left_out[12] ,
    \sb_1__1__43_chanx_left_out[13] ,
    \sb_1__1__43_chanx_left_out[14] ,
    \sb_1__1__43_chanx_left_out[15] ,
    \sb_1__1__43_chanx_left_out[16] ,
    \sb_1__1__43_chanx_left_out[17] ,
    \sb_1__1__43_chanx_left_out[18] ,
    \sb_1__1__43_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__50_chanx_left_out[0] ,
    \cbx_1__1__50_chanx_left_out[1] ,
    \cbx_1__1__50_chanx_left_out[2] ,
    \cbx_1__1__50_chanx_left_out[3] ,
    \cbx_1__1__50_chanx_left_out[4] ,
    \cbx_1__1__50_chanx_left_out[5] ,
    \cbx_1__1__50_chanx_left_out[6] ,
    \cbx_1__1__50_chanx_left_out[7] ,
    \cbx_1__1__50_chanx_left_out[8] ,
    \cbx_1__1__50_chanx_left_out[9] ,
    \cbx_1__1__50_chanx_left_out[10] ,
    \cbx_1__1__50_chanx_left_out[11] ,
    \cbx_1__1__50_chanx_left_out[12] ,
    \cbx_1__1__50_chanx_left_out[13] ,
    \cbx_1__1__50_chanx_left_out[14] ,
    \cbx_1__1__50_chanx_left_out[15] ,
    \cbx_1__1__50_chanx_left_out[16] ,
    \cbx_1__1__50_chanx_left_out[17] ,
    \cbx_1__1__50_chanx_left_out[18] ,
    \cbx_1__1__50_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__43_chanx_right_out[0] ,
    \sb_1__1__43_chanx_right_out[1] ,
    \sb_1__1__43_chanx_right_out[2] ,
    \sb_1__1__43_chanx_right_out[3] ,
    \sb_1__1__43_chanx_right_out[4] ,
    \sb_1__1__43_chanx_right_out[5] ,
    \sb_1__1__43_chanx_right_out[6] ,
    \sb_1__1__43_chanx_right_out[7] ,
    \sb_1__1__43_chanx_right_out[8] ,
    \sb_1__1__43_chanx_right_out[9] ,
    \sb_1__1__43_chanx_right_out[10] ,
    \sb_1__1__43_chanx_right_out[11] ,
    \sb_1__1__43_chanx_right_out[12] ,
    \sb_1__1__43_chanx_right_out[13] ,
    \sb_1__1__43_chanx_right_out[14] ,
    \sb_1__1__43_chanx_right_out[15] ,
    \sb_1__1__43_chanx_right_out[16] ,
    \sb_1__1__43_chanx_right_out[17] ,
    \sb_1__1__43_chanx_right_out[18] ,
    \sb_1__1__43_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__49_chany_top_out[0] ,
    \cby_1__1__49_chany_top_out[1] ,
    \cby_1__1__49_chany_top_out[2] ,
    \cby_1__1__49_chany_top_out[3] ,
    \cby_1__1__49_chany_top_out[4] ,
    \cby_1__1__49_chany_top_out[5] ,
    \cby_1__1__49_chany_top_out[6] ,
    \cby_1__1__49_chany_top_out[7] ,
    \cby_1__1__49_chany_top_out[8] ,
    \cby_1__1__49_chany_top_out[9] ,
    \cby_1__1__49_chany_top_out[10] ,
    \cby_1__1__49_chany_top_out[11] ,
    \cby_1__1__49_chany_top_out[12] ,
    \cby_1__1__49_chany_top_out[13] ,
    \cby_1__1__49_chany_top_out[14] ,
    \cby_1__1__49_chany_top_out[15] ,
    \cby_1__1__49_chany_top_out[16] ,
    \cby_1__1__49_chany_top_out[17] ,
    \cby_1__1__49_chany_top_out[18] ,
    \cby_1__1__49_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__43_chany_bottom_out[0] ,
    \sb_1__1__43_chany_bottom_out[1] ,
    \sb_1__1__43_chany_bottom_out[2] ,
    \sb_1__1__43_chany_bottom_out[3] ,
    \sb_1__1__43_chany_bottom_out[4] ,
    \sb_1__1__43_chany_bottom_out[5] ,
    \sb_1__1__43_chany_bottom_out[6] ,
    \sb_1__1__43_chany_bottom_out[7] ,
    \sb_1__1__43_chany_bottom_out[8] ,
    \sb_1__1__43_chany_bottom_out[9] ,
    \sb_1__1__43_chany_bottom_out[10] ,
    \sb_1__1__43_chany_bottom_out[11] ,
    \sb_1__1__43_chany_bottom_out[12] ,
    \sb_1__1__43_chany_bottom_out[13] ,
    \sb_1__1__43_chany_bottom_out[14] ,
    \sb_1__1__43_chany_bottom_out[15] ,
    \sb_1__1__43_chany_bottom_out[16] ,
    \sb_1__1__43_chany_bottom_out[17] ,
    \sb_1__1__43_chany_bottom_out[18] ,
    \sb_1__1__43_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__50_chany_bottom_out[0] ,
    \cby_1__1__50_chany_bottom_out[1] ,
    \cby_1__1__50_chany_bottom_out[2] ,
    \cby_1__1__50_chany_bottom_out[3] ,
    \cby_1__1__50_chany_bottom_out[4] ,
    \cby_1__1__50_chany_bottom_out[5] ,
    \cby_1__1__50_chany_bottom_out[6] ,
    \cby_1__1__50_chany_bottom_out[7] ,
    \cby_1__1__50_chany_bottom_out[8] ,
    \cby_1__1__50_chany_bottom_out[9] ,
    \cby_1__1__50_chany_bottom_out[10] ,
    \cby_1__1__50_chany_bottom_out[11] ,
    \cby_1__1__50_chany_bottom_out[12] ,
    \cby_1__1__50_chany_bottom_out[13] ,
    \cby_1__1__50_chany_bottom_out[14] ,
    \cby_1__1__50_chany_bottom_out[15] ,
    \cby_1__1__50_chany_bottom_out[16] ,
    \cby_1__1__50_chany_bottom_out[17] ,
    \cby_1__1__50_chany_bottom_out[18] ,
    \cby_1__1__50_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__43_chany_top_out[0] ,
    \sb_1__1__43_chany_top_out[1] ,
    \sb_1__1__43_chany_top_out[2] ,
    \sb_1__1__43_chany_top_out[3] ,
    \sb_1__1__43_chany_top_out[4] ,
    \sb_1__1__43_chany_top_out[5] ,
    \sb_1__1__43_chany_top_out[6] ,
    \sb_1__1__43_chany_top_out[7] ,
    \sb_1__1__43_chany_top_out[8] ,
    \sb_1__1__43_chany_top_out[9] ,
    \sb_1__1__43_chany_top_out[10] ,
    \sb_1__1__43_chany_top_out[11] ,
    \sb_1__1__43_chany_top_out[12] ,
    \sb_1__1__43_chany_top_out[13] ,
    \sb_1__1__43_chany_top_out[14] ,
    \sb_1__1__43_chany_top_out[15] ,
    \sb_1__1__43_chany_top_out[16] ,
    \sb_1__1__43_chany_top_out[17] ,
    \sb_1__1__43_chany_top_out[18] ,
    \sb_1__1__43_chany_top_out[19] }));
 sb_1__1_ sb_7__3_ (.bottom_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__51_ccff_tail),
    .ccff_tail(sb_1__1__44_ccff_tail),
    .clk_1_E_out(\clk_1_wires[92] ),
    .clk_1_N_in(\clk_2_wires[36] ),
    .clk_1_W_out(\clk_1_wires[93] ),
    .left_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[184] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[92] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[36] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[93] ),
    .right_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__44_chanx_right_out[0] ,
    \cbx_1__1__44_chanx_right_out[1] ,
    \cbx_1__1__44_chanx_right_out[2] ,
    \cbx_1__1__44_chanx_right_out[3] ,
    \cbx_1__1__44_chanx_right_out[4] ,
    \cbx_1__1__44_chanx_right_out[5] ,
    \cbx_1__1__44_chanx_right_out[6] ,
    \cbx_1__1__44_chanx_right_out[7] ,
    \cbx_1__1__44_chanx_right_out[8] ,
    \cbx_1__1__44_chanx_right_out[9] ,
    \cbx_1__1__44_chanx_right_out[10] ,
    \cbx_1__1__44_chanx_right_out[11] ,
    \cbx_1__1__44_chanx_right_out[12] ,
    \cbx_1__1__44_chanx_right_out[13] ,
    \cbx_1__1__44_chanx_right_out[14] ,
    \cbx_1__1__44_chanx_right_out[15] ,
    \cbx_1__1__44_chanx_right_out[16] ,
    \cbx_1__1__44_chanx_right_out[17] ,
    \cbx_1__1__44_chanx_right_out[18] ,
    \cbx_1__1__44_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__44_chanx_left_out[0] ,
    \sb_1__1__44_chanx_left_out[1] ,
    \sb_1__1__44_chanx_left_out[2] ,
    \sb_1__1__44_chanx_left_out[3] ,
    \sb_1__1__44_chanx_left_out[4] ,
    \sb_1__1__44_chanx_left_out[5] ,
    \sb_1__1__44_chanx_left_out[6] ,
    \sb_1__1__44_chanx_left_out[7] ,
    \sb_1__1__44_chanx_left_out[8] ,
    \sb_1__1__44_chanx_left_out[9] ,
    \sb_1__1__44_chanx_left_out[10] ,
    \sb_1__1__44_chanx_left_out[11] ,
    \sb_1__1__44_chanx_left_out[12] ,
    \sb_1__1__44_chanx_left_out[13] ,
    \sb_1__1__44_chanx_left_out[14] ,
    \sb_1__1__44_chanx_left_out[15] ,
    \sb_1__1__44_chanx_left_out[16] ,
    \sb_1__1__44_chanx_left_out[17] ,
    \sb_1__1__44_chanx_left_out[18] ,
    \sb_1__1__44_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__51_chanx_left_out[0] ,
    \cbx_1__1__51_chanx_left_out[1] ,
    \cbx_1__1__51_chanx_left_out[2] ,
    \cbx_1__1__51_chanx_left_out[3] ,
    \cbx_1__1__51_chanx_left_out[4] ,
    \cbx_1__1__51_chanx_left_out[5] ,
    \cbx_1__1__51_chanx_left_out[6] ,
    \cbx_1__1__51_chanx_left_out[7] ,
    \cbx_1__1__51_chanx_left_out[8] ,
    \cbx_1__1__51_chanx_left_out[9] ,
    \cbx_1__1__51_chanx_left_out[10] ,
    \cbx_1__1__51_chanx_left_out[11] ,
    \cbx_1__1__51_chanx_left_out[12] ,
    \cbx_1__1__51_chanx_left_out[13] ,
    \cbx_1__1__51_chanx_left_out[14] ,
    \cbx_1__1__51_chanx_left_out[15] ,
    \cbx_1__1__51_chanx_left_out[16] ,
    \cbx_1__1__51_chanx_left_out[17] ,
    \cbx_1__1__51_chanx_left_out[18] ,
    \cbx_1__1__51_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__44_chanx_right_out[0] ,
    \sb_1__1__44_chanx_right_out[1] ,
    \sb_1__1__44_chanx_right_out[2] ,
    \sb_1__1__44_chanx_right_out[3] ,
    \sb_1__1__44_chanx_right_out[4] ,
    \sb_1__1__44_chanx_right_out[5] ,
    \sb_1__1__44_chanx_right_out[6] ,
    \sb_1__1__44_chanx_right_out[7] ,
    \sb_1__1__44_chanx_right_out[8] ,
    \sb_1__1__44_chanx_right_out[9] ,
    \sb_1__1__44_chanx_right_out[10] ,
    \sb_1__1__44_chanx_right_out[11] ,
    \sb_1__1__44_chanx_right_out[12] ,
    \sb_1__1__44_chanx_right_out[13] ,
    \sb_1__1__44_chanx_right_out[14] ,
    \sb_1__1__44_chanx_right_out[15] ,
    \sb_1__1__44_chanx_right_out[16] ,
    \sb_1__1__44_chanx_right_out[17] ,
    \sb_1__1__44_chanx_right_out[18] ,
    \sb_1__1__44_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__50_chany_top_out[0] ,
    \cby_1__1__50_chany_top_out[1] ,
    \cby_1__1__50_chany_top_out[2] ,
    \cby_1__1__50_chany_top_out[3] ,
    \cby_1__1__50_chany_top_out[4] ,
    \cby_1__1__50_chany_top_out[5] ,
    \cby_1__1__50_chany_top_out[6] ,
    \cby_1__1__50_chany_top_out[7] ,
    \cby_1__1__50_chany_top_out[8] ,
    \cby_1__1__50_chany_top_out[9] ,
    \cby_1__1__50_chany_top_out[10] ,
    \cby_1__1__50_chany_top_out[11] ,
    \cby_1__1__50_chany_top_out[12] ,
    \cby_1__1__50_chany_top_out[13] ,
    \cby_1__1__50_chany_top_out[14] ,
    \cby_1__1__50_chany_top_out[15] ,
    \cby_1__1__50_chany_top_out[16] ,
    \cby_1__1__50_chany_top_out[17] ,
    \cby_1__1__50_chany_top_out[18] ,
    \cby_1__1__50_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__44_chany_bottom_out[0] ,
    \sb_1__1__44_chany_bottom_out[1] ,
    \sb_1__1__44_chany_bottom_out[2] ,
    \sb_1__1__44_chany_bottom_out[3] ,
    \sb_1__1__44_chany_bottom_out[4] ,
    \sb_1__1__44_chany_bottom_out[5] ,
    \sb_1__1__44_chany_bottom_out[6] ,
    \sb_1__1__44_chany_bottom_out[7] ,
    \sb_1__1__44_chany_bottom_out[8] ,
    \sb_1__1__44_chany_bottom_out[9] ,
    \sb_1__1__44_chany_bottom_out[10] ,
    \sb_1__1__44_chany_bottom_out[11] ,
    \sb_1__1__44_chany_bottom_out[12] ,
    \sb_1__1__44_chany_bottom_out[13] ,
    \sb_1__1__44_chany_bottom_out[14] ,
    \sb_1__1__44_chany_bottom_out[15] ,
    \sb_1__1__44_chany_bottom_out[16] ,
    \sb_1__1__44_chany_bottom_out[17] ,
    \sb_1__1__44_chany_bottom_out[18] ,
    \sb_1__1__44_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__51_chany_bottom_out[0] ,
    \cby_1__1__51_chany_bottom_out[1] ,
    \cby_1__1__51_chany_bottom_out[2] ,
    \cby_1__1__51_chany_bottom_out[3] ,
    \cby_1__1__51_chany_bottom_out[4] ,
    \cby_1__1__51_chany_bottom_out[5] ,
    \cby_1__1__51_chany_bottom_out[6] ,
    \cby_1__1__51_chany_bottom_out[7] ,
    \cby_1__1__51_chany_bottom_out[8] ,
    \cby_1__1__51_chany_bottom_out[9] ,
    \cby_1__1__51_chany_bottom_out[10] ,
    \cby_1__1__51_chany_bottom_out[11] ,
    \cby_1__1__51_chany_bottom_out[12] ,
    \cby_1__1__51_chany_bottom_out[13] ,
    \cby_1__1__51_chany_bottom_out[14] ,
    \cby_1__1__51_chany_bottom_out[15] ,
    \cby_1__1__51_chany_bottom_out[16] ,
    \cby_1__1__51_chany_bottom_out[17] ,
    \cby_1__1__51_chany_bottom_out[18] ,
    \cby_1__1__51_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__44_chany_top_out[0] ,
    \sb_1__1__44_chany_top_out[1] ,
    \sb_1__1__44_chany_top_out[2] ,
    \sb_1__1__44_chany_top_out[3] ,
    \sb_1__1__44_chany_top_out[4] ,
    \sb_1__1__44_chany_top_out[5] ,
    \sb_1__1__44_chany_top_out[6] ,
    \sb_1__1__44_chany_top_out[7] ,
    \sb_1__1__44_chany_top_out[8] ,
    \sb_1__1__44_chany_top_out[9] ,
    \sb_1__1__44_chany_top_out[10] ,
    \sb_1__1__44_chany_top_out[11] ,
    \sb_1__1__44_chany_top_out[12] ,
    \sb_1__1__44_chany_top_out[13] ,
    \sb_1__1__44_chany_top_out[14] ,
    \sb_1__1__44_chany_top_out[15] ,
    \sb_1__1__44_chany_top_out[16] ,
    \sb_1__1__44_chany_top_out[17] ,
    \sb_1__1__44_chany_top_out[18] ,
    \sb_1__1__44_chany_top_out[19] }));
 sb_1__1_ sb_7__4_ (.bottom_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__52_ccff_tail),
    .ccff_tail(sb_1__1__45_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[187] ),
    .right_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__45_chanx_right_out[0] ,
    \cbx_1__1__45_chanx_right_out[1] ,
    \cbx_1__1__45_chanx_right_out[2] ,
    \cbx_1__1__45_chanx_right_out[3] ,
    \cbx_1__1__45_chanx_right_out[4] ,
    \cbx_1__1__45_chanx_right_out[5] ,
    \cbx_1__1__45_chanx_right_out[6] ,
    \cbx_1__1__45_chanx_right_out[7] ,
    \cbx_1__1__45_chanx_right_out[8] ,
    \cbx_1__1__45_chanx_right_out[9] ,
    \cbx_1__1__45_chanx_right_out[10] ,
    \cbx_1__1__45_chanx_right_out[11] ,
    \cbx_1__1__45_chanx_right_out[12] ,
    \cbx_1__1__45_chanx_right_out[13] ,
    \cbx_1__1__45_chanx_right_out[14] ,
    \cbx_1__1__45_chanx_right_out[15] ,
    \cbx_1__1__45_chanx_right_out[16] ,
    \cbx_1__1__45_chanx_right_out[17] ,
    \cbx_1__1__45_chanx_right_out[18] ,
    \cbx_1__1__45_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__45_chanx_left_out[0] ,
    \sb_1__1__45_chanx_left_out[1] ,
    \sb_1__1__45_chanx_left_out[2] ,
    \sb_1__1__45_chanx_left_out[3] ,
    \sb_1__1__45_chanx_left_out[4] ,
    \sb_1__1__45_chanx_left_out[5] ,
    \sb_1__1__45_chanx_left_out[6] ,
    \sb_1__1__45_chanx_left_out[7] ,
    \sb_1__1__45_chanx_left_out[8] ,
    \sb_1__1__45_chanx_left_out[9] ,
    \sb_1__1__45_chanx_left_out[10] ,
    \sb_1__1__45_chanx_left_out[11] ,
    \sb_1__1__45_chanx_left_out[12] ,
    \sb_1__1__45_chanx_left_out[13] ,
    \sb_1__1__45_chanx_left_out[14] ,
    \sb_1__1__45_chanx_left_out[15] ,
    \sb_1__1__45_chanx_left_out[16] ,
    \sb_1__1__45_chanx_left_out[17] ,
    \sb_1__1__45_chanx_left_out[18] ,
    \sb_1__1__45_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__52_chanx_left_out[0] ,
    \cbx_1__1__52_chanx_left_out[1] ,
    \cbx_1__1__52_chanx_left_out[2] ,
    \cbx_1__1__52_chanx_left_out[3] ,
    \cbx_1__1__52_chanx_left_out[4] ,
    \cbx_1__1__52_chanx_left_out[5] ,
    \cbx_1__1__52_chanx_left_out[6] ,
    \cbx_1__1__52_chanx_left_out[7] ,
    \cbx_1__1__52_chanx_left_out[8] ,
    \cbx_1__1__52_chanx_left_out[9] ,
    \cbx_1__1__52_chanx_left_out[10] ,
    \cbx_1__1__52_chanx_left_out[11] ,
    \cbx_1__1__52_chanx_left_out[12] ,
    \cbx_1__1__52_chanx_left_out[13] ,
    \cbx_1__1__52_chanx_left_out[14] ,
    \cbx_1__1__52_chanx_left_out[15] ,
    \cbx_1__1__52_chanx_left_out[16] ,
    \cbx_1__1__52_chanx_left_out[17] ,
    \cbx_1__1__52_chanx_left_out[18] ,
    \cbx_1__1__52_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__45_chanx_right_out[0] ,
    \sb_1__1__45_chanx_right_out[1] ,
    \sb_1__1__45_chanx_right_out[2] ,
    \sb_1__1__45_chanx_right_out[3] ,
    \sb_1__1__45_chanx_right_out[4] ,
    \sb_1__1__45_chanx_right_out[5] ,
    \sb_1__1__45_chanx_right_out[6] ,
    \sb_1__1__45_chanx_right_out[7] ,
    \sb_1__1__45_chanx_right_out[8] ,
    \sb_1__1__45_chanx_right_out[9] ,
    \sb_1__1__45_chanx_right_out[10] ,
    \sb_1__1__45_chanx_right_out[11] ,
    \sb_1__1__45_chanx_right_out[12] ,
    \sb_1__1__45_chanx_right_out[13] ,
    \sb_1__1__45_chanx_right_out[14] ,
    \sb_1__1__45_chanx_right_out[15] ,
    \sb_1__1__45_chanx_right_out[16] ,
    \sb_1__1__45_chanx_right_out[17] ,
    \sb_1__1__45_chanx_right_out[18] ,
    \sb_1__1__45_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__51_chany_top_out[0] ,
    \cby_1__1__51_chany_top_out[1] ,
    \cby_1__1__51_chany_top_out[2] ,
    \cby_1__1__51_chany_top_out[3] ,
    \cby_1__1__51_chany_top_out[4] ,
    \cby_1__1__51_chany_top_out[5] ,
    \cby_1__1__51_chany_top_out[6] ,
    \cby_1__1__51_chany_top_out[7] ,
    \cby_1__1__51_chany_top_out[8] ,
    \cby_1__1__51_chany_top_out[9] ,
    \cby_1__1__51_chany_top_out[10] ,
    \cby_1__1__51_chany_top_out[11] ,
    \cby_1__1__51_chany_top_out[12] ,
    \cby_1__1__51_chany_top_out[13] ,
    \cby_1__1__51_chany_top_out[14] ,
    \cby_1__1__51_chany_top_out[15] ,
    \cby_1__1__51_chany_top_out[16] ,
    \cby_1__1__51_chany_top_out[17] ,
    \cby_1__1__51_chany_top_out[18] ,
    \cby_1__1__51_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__45_chany_bottom_out[0] ,
    \sb_1__1__45_chany_bottom_out[1] ,
    \sb_1__1__45_chany_bottom_out[2] ,
    \sb_1__1__45_chany_bottom_out[3] ,
    \sb_1__1__45_chany_bottom_out[4] ,
    \sb_1__1__45_chany_bottom_out[5] ,
    \sb_1__1__45_chany_bottom_out[6] ,
    \sb_1__1__45_chany_bottom_out[7] ,
    \sb_1__1__45_chany_bottom_out[8] ,
    \sb_1__1__45_chany_bottom_out[9] ,
    \sb_1__1__45_chany_bottom_out[10] ,
    \sb_1__1__45_chany_bottom_out[11] ,
    \sb_1__1__45_chany_bottom_out[12] ,
    \sb_1__1__45_chany_bottom_out[13] ,
    \sb_1__1__45_chany_bottom_out[14] ,
    \sb_1__1__45_chany_bottom_out[15] ,
    \sb_1__1__45_chany_bottom_out[16] ,
    \sb_1__1__45_chany_bottom_out[17] ,
    \sb_1__1__45_chany_bottom_out[18] ,
    \sb_1__1__45_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__52_chany_bottom_out[0] ,
    \cby_1__1__52_chany_bottom_out[1] ,
    \cby_1__1__52_chany_bottom_out[2] ,
    \cby_1__1__52_chany_bottom_out[3] ,
    \cby_1__1__52_chany_bottom_out[4] ,
    \cby_1__1__52_chany_bottom_out[5] ,
    \cby_1__1__52_chany_bottom_out[6] ,
    \cby_1__1__52_chany_bottom_out[7] ,
    \cby_1__1__52_chany_bottom_out[8] ,
    \cby_1__1__52_chany_bottom_out[9] ,
    \cby_1__1__52_chany_bottom_out[10] ,
    \cby_1__1__52_chany_bottom_out[11] ,
    \cby_1__1__52_chany_bottom_out[12] ,
    \cby_1__1__52_chany_bottom_out[13] ,
    \cby_1__1__52_chany_bottom_out[14] ,
    \cby_1__1__52_chany_bottom_out[15] ,
    \cby_1__1__52_chany_bottom_out[16] ,
    \cby_1__1__52_chany_bottom_out[17] ,
    \cby_1__1__52_chany_bottom_out[18] ,
    \cby_1__1__52_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__45_chany_top_out[0] ,
    \sb_1__1__45_chany_top_out[1] ,
    \sb_1__1__45_chany_top_out[2] ,
    \sb_1__1__45_chany_top_out[3] ,
    \sb_1__1__45_chany_top_out[4] ,
    \sb_1__1__45_chany_top_out[5] ,
    \sb_1__1__45_chany_top_out[6] ,
    \sb_1__1__45_chany_top_out[7] ,
    \sb_1__1__45_chany_top_out[8] ,
    \sb_1__1__45_chany_top_out[9] ,
    \sb_1__1__45_chany_top_out[10] ,
    \sb_1__1__45_chany_top_out[11] ,
    \sb_1__1__45_chany_top_out[12] ,
    \sb_1__1__45_chany_top_out[13] ,
    \sb_1__1__45_chany_top_out[14] ,
    \sb_1__1__45_chany_top_out[15] ,
    \sb_1__1__45_chany_top_out[16] ,
    \sb_1__1__45_chany_top_out[17] ,
    \sb_1__1__45_chany_top_out[18] ,
    \sb_1__1__45_chany_top_out[19] }));
 sb_1__1_ sb_7__5_ (.bottom_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__53_ccff_tail),
    .ccff_tail(sb_1__1__46_ccff_tail),
    .clk_1_E_out(\clk_1_wires[99] ),
    .clk_1_N_in(\clk_2_wires[51] ),
    .clk_1_W_out(\clk_1_wires[100] ),
    .left_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[190] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[99] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[51] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[100] ),
    .right_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__46_chanx_right_out[0] ,
    \cbx_1__1__46_chanx_right_out[1] ,
    \cbx_1__1__46_chanx_right_out[2] ,
    \cbx_1__1__46_chanx_right_out[3] ,
    \cbx_1__1__46_chanx_right_out[4] ,
    \cbx_1__1__46_chanx_right_out[5] ,
    \cbx_1__1__46_chanx_right_out[6] ,
    \cbx_1__1__46_chanx_right_out[7] ,
    \cbx_1__1__46_chanx_right_out[8] ,
    \cbx_1__1__46_chanx_right_out[9] ,
    \cbx_1__1__46_chanx_right_out[10] ,
    \cbx_1__1__46_chanx_right_out[11] ,
    \cbx_1__1__46_chanx_right_out[12] ,
    \cbx_1__1__46_chanx_right_out[13] ,
    \cbx_1__1__46_chanx_right_out[14] ,
    \cbx_1__1__46_chanx_right_out[15] ,
    \cbx_1__1__46_chanx_right_out[16] ,
    \cbx_1__1__46_chanx_right_out[17] ,
    \cbx_1__1__46_chanx_right_out[18] ,
    \cbx_1__1__46_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__46_chanx_left_out[0] ,
    \sb_1__1__46_chanx_left_out[1] ,
    \sb_1__1__46_chanx_left_out[2] ,
    \sb_1__1__46_chanx_left_out[3] ,
    \sb_1__1__46_chanx_left_out[4] ,
    \sb_1__1__46_chanx_left_out[5] ,
    \sb_1__1__46_chanx_left_out[6] ,
    \sb_1__1__46_chanx_left_out[7] ,
    \sb_1__1__46_chanx_left_out[8] ,
    \sb_1__1__46_chanx_left_out[9] ,
    \sb_1__1__46_chanx_left_out[10] ,
    \sb_1__1__46_chanx_left_out[11] ,
    \sb_1__1__46_chanx_left_out[12] ,
    \sb_1__1__46_chanx_left_out[13] ,
    \sb_1__1__46_chanx_left_out[14] ,
    \sb_1__1__46_chanx_left_out[15] ,
    \sb_1__1__46_chanx_left_out[16] ,
    \sb_1__1__46_chanx_left_out[17] ,
    \sb_1__1__46_chanx_left_out[18] ,
    \sb_1__1__46_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__53_chanx_left_out[0] ,
    \cbx_1__1__53_chanx_left_out[1] ,
    \cbx_1__1__53_chanx_left_out[2] ,
    \cbx_1__1__53_chanx_left_out[3] ,
    \cbx_1__1__53_chanx_left_out[4] ,
    \cbx_1__1__53_chanx_left_out[5] ,
    \cbx_1__1__53_chanx_left_out[6] ,
    \cbx_1__1__53_chanx_left_out[7] ,
    \cbx_1__1__53_chanx_left_out[8] ,
    \cbx_1__1__53_chanx_left_out[9] ,
    \cbx_1__1__53_chanx_left_out[10] ,
    \cbx_1__1__53_chanx_left_out[11] ,
    \cbx_1__1__53_chanx_left_out[12] ,
    \cbx_1__1__53_chanx_left_out[13] ,
    \cbx_1__1__53_chanx_left_out[14] ,
    \cbx_1__1__53_chanx_left_out[15] ,
    \cbx_1__1__53_chanx_left_out[16] ,
    \cbx_1__1__53_chanx_left_out[17] ,
    \cbx_1__1__53_chanx_left_out[18] ,
    \cbx_1__1__53_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__46_chanx_right_out[0] ,
    \sb_1__1__46_chanx_right_out[1] ,
    \sb_1__1__46_chanx_right_out[2] ,
    \sb_1__1__46_chanx_right_out[3] ,
    \sb_1__1__46_chanx_right_out[4] ,
    \sb_1__1__46_chanx_right_out[5] ,
    \sb_1__1__46_chanx_right_out[6] ,
    \sb_1__1__46_chanx_right_out[7] ,
    \sb_1__1__46_chanx_right_out[8] ,
    \sb_1__1__46_chanx_right_out[9] ,
    \sb_1__1__46_chanx_right_out[10] ,
    \sb_1__1__46_chanx_right_out[11] ,
    \sb_1__1__46_chanx_right_out[12] ,
    \sb_1__1__46_chanx_right_out[13] ,
    \sb_1__1__46_chanx_right_out[14] ,
    \sb_1__1__46_chanx_right_out[15] ,
    \sb_1__1__46_chanx_right_out[16] ,
    \sb_1__1__46_chanx_right_out[17] ,
    \sb_1__1__46_chanx_right_out[18] ,
    \sb_1__1__46_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__52_chany_top_out[0] ,
    \cby_1__1__52_chany_top_out[1] ,
    \cby_1__1__52_chany_top_out[2] ,
    \cby_1__1__52_chany_top_out[3] ,
    \cby_1__1__52_chany_top_out[4] ,
    \cby_1__1__52_chany_top_out[5] ,
    \cby_1__1__52_chany_top_out[6] ,
    \cby_1__1__52_chany_top_out[7] ,
    \cby_1__1__52_chany_top_out[8] ,
    \cby_1__1__52_chany_top_out[9] ,
    \cby_1__1__52_chany_top_out[10] ,
    \cby_1__1__52_chany_top_out[11] ,
    \cby_1__1__52_chany_top_out[12] ,
    \cby_1__1__52_chany_top_out[13] ,
    \cby_1__1__52_chany_top_out[14] ,
    \cby_1__1__52_chany_top_out[15] ,
    \cby_1__1__52_chany_top_out[16] ,
    \cby_1__1__52_chany_top_out[17] ,
    \cby_1__1__52_chany_top_out[18] ,
    \cby_1__1__52_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__46_chany_bottom_out[0] ,
    \sb_1__1__46_chany_bottom_out[1] ,
    \sb_1__1__46_chany_bottom_out[2] ,
    \sb_1__1__46_chany_bottom_out[3] ,
    \sb_1__1__46_chany_bottom_out[4] ,
    \sb_1__1__46_chany_bottom_out[5] ,
    \sb_1__1__46_chany_bottom_out[6] ,
    \sb_1__1__46_chany_bottom_out[7] ,
    \sb_1__1__46_chany_bottom_out[8] ,
    \sb_1__1__46_chany_bottom_out[9] ,
    \sb_1__1__46_chany_bottom_out[10] ,
    \sb_1__1__46_chany_bottom_out[11] ,
    \sb_1__1__46_chany_bottom_out[12] ,
    \sb_1__1__46_chany_bottom_out[13] ,
    \sb_1__1__46_chany_bottom_out[14] ,
    \sb_1__1__46_chany_bottom_out[15] ,
    \sb_1__1__46_chany_bottom_out[16] ,
    \sb_1__1__46_chany_bottom_out[17] ,
    \sb_1__1__46_chany_bottom_out[18] ,
    \sb_1__1__46_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__53_chany_bottom_out[0] ,
    \cby_1__1__53_chany_bottom_out[1] ,
    \cby_1__1__53_chany_bottom_out[2] ,
    \cby_1__1__53_chany_bottom_out[3] ,
    \cby_1__1__53_chany_bottom_out[4] ,
    \cby_1__1__53_chany_bottom_out[5] ,
    \cby_1__1__53_chany_bottom_out[6] ,
    \cby_1__1__53_chany_bottom_out[7] ,
    \cby_1__1__53_chany_bottom_out[8] ,
    \cby_1__1__53_chany_bottom_out[9] ,
    \cby_1__1__53_chany_bottom_out[10] ,
    \cby_1__1__53_chany_bottom_out[11] ,
    \cby_1__1__53_chany_bottom_out[12] ,
    \cby_1__1__53_chany_bottom_out[13] ,
    \cby_1__1__53_chany_bottom_out[14] ,
    \cby_1__1__53_chany_bottom_out[15] ,
    \cby_1__1__53_chany_bottom_out[16] ,
    \cby_1__1__53_chany_bottom_out[17] ,
    \cby_1__1__53_chany_bottom_out[18] ,
    \cby_1__1__53_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__46_chany_top_out[0] ,
    \sb_1__1__46_chany_top_out[1] ,
    \sb_1__1__46_chany_top_out[2] ,
    \sb_1__1__46_chany_top_out[3] ,
    \sb_1__1__46_chany_top_out[4] ,
    \sb_1__1__46_chany_top_out[5] ,
    \sb_1__1__46_chany_top_out[6] ,
    \sb_1__1__46_chany_top_out[7] ,
    \sb_1__1__46_chany_top_out[8] ,
    \sb_1__1__46_chany_top_out[9] ,
    \sb_1__1__46_chany_top_out[10] ,
    \sb_1__1__46_chany_top_out[11] ,
    \sb_1__1__46_chany_top_out[12] ,
    \sb_1__1__46_chany_top_out[13] ,
    \sb_1__1__46_chany_top_out[14] ,
    \sb_1__1__46_chany_top_out[15] ,
    \sb_1__1__46_chany_top_out[16] ,
    \sb_1__1__46_chany_top_out[17] ,
    \sb_1__1__46_chany_top_out[18] ,
    \sb_1__1__46_chany_top_out[19] }));
 sb_1__1_ sb_7__6_ (.bottom_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__54_ccff_tail),
    .ccff_tail(sb_1__1__47_ccff_tail),
    .clk_2_N_in(\clk_2_wires[41] ),
    .clk_2_N_out(\clk_2_wires[48] ),
    .clk_2_S_out(\clk_2_wires[50] ),
    .left_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[193] ),
    .prog_clk_2_N_in(\prog_clk_2_wires[41] ),
    .prog_clk_2_N_out(\prog_clk_2_wires[48] ),
    .prog_clk_2_S_out(\prog_clk_2_wires[50] ),
    .right_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__47_chanx_right_out[0] ,
    \cbx_1__1__47_chanx_right_out[1] ,
    \cbx_1__1__47_chanx_right_out[2] ,
    \cbx_1__1__47_chanx_right_out[3] ,
    \cbx_1__1__47_chanx_right_out[4] ,
    \cbx_1__1__47_chanx_right_out[5] ,
    \cbx_1__1__47_chanx_right_out[6] ,
    \cbx_1__1__47_chanx_right_out[7] ,
    \cbx_1__1__47_chanx_right_out[8] ,
    \cbx_1__1__47_chanx_right_out[9] ,
    \cbx_1__1__47_chanx_right_out[10] ,
    \cbx_1__1__47_chanx_right_out[11] ,
    \cbx_1__1__47_chanx_right_out[12] ,
    \cbx_1__1__47_chanx_right_out[13] ,
    \cbx_1__1__47_chanx_right_out[14] ,
    \cbx_1__1__47_chanx_right_out[15] ,
    \cbx_1__1__47_chanx_right_out[16] ,
    \cbx_1__1__47_chanx_right_out[17] ,
    \cbx_1__1__47_chanx_right_out[18] ,
    \cbx_1__1__47_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__47_chanx_left_out[0] ,
    \sb_1__1__47_chanx_left_out[1] ,
    \sb_1__1__47_chanx_left_out[2] ,
    \sb_1__1__47_chanx_left_out[3] ,
    \sb_1__1__47_chanx_left_out[4] ,
    \sb_1__1__47_chanx_left_out[5] ,
    \sb_1__1__47_chanx_left_out[6] ,
    \sb_1__1__47_chanx_left_out[7] ,
    \sb_1__1__47_chanx_left_out[8] ,
    \sb_1__1__47_chanx_left_out[9] ,
    \sb_1__1__47_chanx_left_out[10] ,
    \sb_1__1__47_chanx_left_out[11] ,
    \sb_1__1__47_chanx_left_out[12] ,
    \sb_1__1__47_chanx_left_out[13] ,
    \sb_1__1__47_chanx_left_out[14] ,
    \sb_1__1__47_chanx_left_out[15] ,
    \sb_1__1__47_chanx_left_out[16] ,
    \sb_1__1__47_chanx_left_out[17] ,
    \sb_1__1__47_chanx_left_out[18] ,
    \sb_1__1__47_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__54_chanx_left_out[0] ,
    \cbx_1__1__54_chanx_left_out[1] ,
    \cbx_1__1__54_chanx_left_out[2] ,
    \cbx_1__1__54_chanx_left_out[3] ,
    \cbx_1__1__54_chanx_left_out[4] ,
    \cbx_1__1__54_chanx_left_out[5] ,
    \cbx_1__1__54_chanx_left_out[6] ,
    \cbx_1__1__54_chanx_left_out[7] ,
    \cbx_1__1__54_chanx_left_out[8] ,
    \cbx_1__1__54_chanx_left_out[9] ,
    \cbx_1__1__54_chanx_left_out[10] ,
    \cbx_1__1__54_chanx_left_out[11] ,
    \cbx_1__1__54_chanx_left_out[12] ,
    \cbx_1__1__54_chanx_left_out[13] ,
    \cbx_1__1__54_chanx_left_out[14] ,
    \cbx_1__1__54_chanx_left_out[15] ,
    \cbx_1__1__54_chanx_left_out[16] ,
    \cbx_1__1__54_chanx_left_out[17] ,
    \cbx_1__1__54_chanx_left_out[18] ,
    \cbx_1__1__54_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__47_chanx_right_out[0] ,
    \sb_1__1__47_chanx_right_out[1] ,
    \sb_1__1__47_chanx_right_out[2] ,
    \sb_1__1__47_chanx_right_out[3] ,
    \sb_1__1__47_chanx_right_out[4] ,
    \sb_1__1__47_chanx_right_out[5] ,
    \sb_1__1__47_chanx_right_out[6] ,
    \sb_1__1__47_chanx_right_out[7] ,
    \sb_1__1__47_chanx_right_out[8] ,
    \sb_1__1__47_chanx_right_out[9] ,
    \sb_1__1__47_chanx_right_out[10] ,
    \sb_1__1__47_chanx_right_out[11] ,
    \sb_1__1__47_chanx_right_out[12] ,
    \sb_1__1__47_chanx_right_out[13] ,
    \sb_1__1__47_chanx_right_out[14] ,
    \sb_1__1__47_chanx_right_out[15] ,
    \sb_1__1__47_chanx_right_out[16] ,
    \sb_1__1__47_chanx_right_out[17] ,
    \sb_1__1__47_chanx_right_out[18] ,
    \sb_1__1__47_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__53_chany_top_out[0] ,
    \cby_1__1__53_chany_top_out[1] ,
    \cby_1__1__53_chany_top_out[2] ,
    \cby_1__1__53_chany_top_out[3] ,
    \cby_1__1__53_chany_top_out[4] ,
    \cby_1__1__53_chany_top_out[5] ,
    \cby_1__1__53_chany_top_out[6] ,
    \cby_1__1__53_chany_top_out[7] ,
    \cby_1__1__53_chany_top_out[8] ,
    \cby_1__1__53_chany_top_out[9] ,
    \cby_1__1__53_chany_top_out[10] ,
    \cby_1__1__53_chany_top_out[11] ,
    \cby_1__1__53_chany_top_out[12] ,
    \cby_1__1__53_chany_top_out[13] ,
    \cby_1__1__53_chany_top_out[14] ,
    \cby_1__1__53_chany_top_out[15] ,
    \cby_1__1__53_chany_top_out[16] ,
    \cby_1__1__53_chany_top_out[17] ,
    \cby_1__1__53_chany_top_out[18] ,
    \cby_1__1__53_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__47_chany_bottom_out[0] ,
    \sb_1__1__47_chany_bottom_out[1] ,
    \sb_1__1__47_chany_bottom_out[2] ,
    \sb_1__1__47_chany_bottom_out[3] ,
    \sb_1__1__47_chany_bottom_out[4] ,
    \sb_1__1__47_chany_bottom_out[5] ,
    \sb_1__1__47_chany_bottom_out[6] ,
    \sb_1__1__47_chany_bottom_out[7] ,
    \sb_1__1__47_chany_bottom_out[8] ,
    \sb_1__1__47_chany_bottom_out[9] ,
    \sb_1__1__47_chany_bottom_out[10] ,
    \sb_1__1__47_chany_bottom_out[11] ,
    \sb_1__1__47_chany_bottom_out[12] ,
    \sb_1__1__47_chany_bottom_out[13] ,
    \sb_1__1__47_chany_bottom_out[14] ,
    \sb_1__1__47_chany_bottom_out[15] ,
    \sb_1__1__47_chany_bottom_out[16] ,
    \sb_1__1__47_chany_bottom_out[17] ,
    \sb_1__1__47_chany_bottom_out[18] ,
    \sb_1__1__47_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__54_chany_bottom_out[0] ,
    \cby_1__1__54_chany_bottom_out[1] ,
    \cby_1__1__54_chany_bottom_out[2] ,
    \cby_1__1__54_chany_bottom_out[3] ,
    \cby_1__1__54_chany_bottom_out[4] ,
    \cby_1__1__54_chany_bottom_out[5] ,
    \cby_1__1__54_chany_bottom_out[6] ,
    \cby_1__1__54_chany_bottom_out[7] ,
    \cby_1__1__54_chany_bottom_out[8] ,
    \cby_1__1__54_chany_bottom_out[9] ,
    \cby_1__1__54_chany_bottom_out[10] ,
    \cby_1__1__54_chany_bottom_out[11] ,
    \cby_1__1__54_chany_bottom_out[12] ,
    \cby_1__1__54_chany_bottom_out[13] ,
    \cby_1__1__54_chany_bottom_out[14] ,
    \cby_1__1__54_chany_bottom_out[15] ,
    \cby_1__1__54_chany_bottom_out[16] ,
    \cby_1__1__54_chany_bottom_out[17] ,
    \cby_1__1__54_chany_bottom_out[18] ,
    \cby_1__1__54_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__47_chany_top_out[0] ,
    \sb_1__1__47_chany_top_out[1] ,
    \sb_1__1__47_chany_top_out[2] ,
    \sb_1__1__47_chany_top_out[3] ,
    \sb_1__1__47_chany_top_out[4] ,
    \sb_1__1__47_chany_top_out[5] ,
    \sb_1__1__47_chany_top_out[6] ,
    \sb_1__1__47_chany_top_out[7] ,
    \sb_1__1__47_chany_top_out[8] ,
    \sb_1__1__47_chany_top_out[9] ,
    \sb_1__1__47_chany_top_out[10] ,
    \sb_1__1__47_chany_top_out[11] ,
    \sb_1__1__47_chany_top_out[12] ,
    \sb_1__1__47_chany_top_out[13] ,
    \sb_1__1__47_chany_top_out[14] ,
    \sb_1__1__47_chany_top_out[15] ,
    \sb_1__1__47_chany_top_out[16] ,
    \sb_1__1__47_chany_top_out[17] ,
    \sb_1__1__47_chany_top_out[18] ,
    \sb_1__1__47_chany_top_out[19] }));
 sb_1__1_ sb_7__7_ (.bottom_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_upper),
    .ccff_head(cbx_1__1__55_ccff_tail),
    .ccff_tail(sb_1__1__48_ccff_tail),
    .clk_1_E_out(\clk_1_wires[106] ),
    .clk_1_N_in(\clk_2_wires[49] ),
    .clk_1_W_out(\clk_1_wires[107] ),
    .left_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[196] ),
    .prog_clk_1_E_out(\prog_clk_1_wires[106] ),
    .prog_clk_1_N_in(\prog_clk_2_wires[49] ),
    .prog_clk_1_W_out(\prog_clk_1_wires[107] ),
    .right_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_upper),
    .top_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__48_chanx_right_out[0] ,
    \cbx_1__1__48_chanx_right_out[1] ,
    \cbx_1__1__48_chanx_right_out[2] ,
    \cbx_1__1__48_chanx_right_out[3] ,
    \cbx_1__1__48_chanx_right_out[4] ,
    \cbx_1__1__48_chanx_right_out[5] ,
    \cbx_1__1__48_chanx_right_out[6] ,
    \cbx_1__1__48_chanx_right_out[7] ,
    \cbx_1__1__48_chanx_right_out[8] ,
    \cbx_1__1__48_chanx_right_out[9] ,
    \cbx_1__1__48_chanx_right_out[10] ,
    \cbx_1__1__48_chanx_right_out[11] ,
    \cbx_1__1__48_chanx_right_out[12] ,
    \cbx_1__1__48_chanx_right_out[13] ,
    \cbx_1__1__48_chanx_right_out[14] ,
    \cbx_1__1__48_chanx_right_out[15] ,
    \cbx_1__1__48_chanx_right_out[16] ,
    \cbx_1__1__48_chanx_right_out[17] ,
    \cbx_1__1__48_chanx_right_out[18] ,
    \cbx_1__1__48_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__1__48_chanx_left_out[0] ,
    \sb_1__1__48_chanx_left_out[1] ,
    \sb_1__1__48_chanx_left_out[2] ,
    \sb_1__1__48_chanx_left_out[3] ,
    \sb_1__1__48_chanx_left_out[4] ,
    \sb_1__1__48_chanx_left_out[5] ,
    \sb_1__1__48_chanx_left_out[6] ,
    \sb_1__1__48_chanx_left_out[7] ,
    \sb_1__1__48_chanx_left_out[8] ,
    \sb_1__1__48_chanx_left_out[9] ,
    \sb_1__1__48_chanx_left_out[10] ,
    \sb_1__1__48_chanx_left_out[11] ,
    \sb_1__1__48_chanx_left_out[12] ,
    \sb_1__1__48_chanx_left_out[13] ,
    \sb_1__1__48_chanx_left_out[14] ,
    \sb_1__1__48_chanx_left_out[15] ,
    \sb_1__1__48_chanx_left_out[16] ,
    \sb_1__1__48_chanx_left_out[17] ,
    \sb_1__1__48_chanx_left_out[18] ,
    \sb_1__1__48_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__1__55_chanx_left_out[0] ,
    \cbx_1__1__55_chanx_left_out[1] ,
    \cbx_1__1__55_chanx_left_out[2] ,
    \cbx_1__1__55_chanx_left_out[3] ,
    \cbx_1__1__55_chanx_left_out[4] ,
    \cbx_1__1__55_chanx_left_out[5] ,
    \cbx_1__1__55_chanx_left_out[6] ,
    \cbx_1__1__55_chanx_left_out[7] ,
    \cbx_1__1__55_chanx_left_out[8] ,
    \cbx_1__1__55_chanx_left_out[9] ,
    \cbx_1__1__55_chanx_left_out[10] ,
    \cbx_1__1__55_chanx_left_out[11] ,
    \cbx_1__1__55_chanx_left_out[12] ,
    \cbx_1__1__55_chanx_left_out[13] ,
    \cbx_1__1__55_chanx_left_out[14] ,
    \cbx_1__1__55_chanx_left_out[15] ,
    \cbx_1__1__55_chanx_left_out[16] ,
    \cbx_1__1__55_chanx_left_out[17] ,
    \cbx_1__1__55_chanx_left_out[18] ,
    \cbx_1__1__55_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__1__48_chanx_right_out[0] ,
    \sb_1__1__48_chanx_right_out[1] ,
    \sb_1__1__48_chanx_right_out[2] ,
    \sb_1__1__48_chanx_right_out[3] ,
    \sb_1__1__48_chanx_right_out[4] ,
    \sb_1__1__48_chanx_right_out[5] ,
    \sb_1__1__48_chanx_right_out[6] ,
    \sb_1__1__48_chanx_right_out[7] ,
    \sb_1__1__48_chanx_right_out[8] ,
    \sb_1__1__48_chanx_right_out[9] ,
    \sb_1__1__48_chanx_right_out[10] ,
    \sb_1__1__48_chanx_right_out[11] ,
    \sb_1__1__48_chanx_right_out[12] ,
    \sb_1__1__48_chanx_right_out[13] ,
    \sb_1__1__48_chanx_right_out[14] ,
    \sb_1__1__48_chanx_right_out[15] ,
    \sb_1__1__48_chanx_right_out[16] ,
    \sb_1__1__48_chanx_right_out[17] ,
    \sb_1__1__48_chanx_right_out[18] ,
    \sb_1__1__48_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__54_chany_top_out[0] ,
    \cby_1__1__54_chany_top_out[1] ,
    \cby_1__1__54_chany_top_out[2] ,
    \cby_1__1__54_chany_top_out[3] ,
    \cby_1__1__54_chany_top_out[4] ,
    \cby_1__1__54_chany_top_out[5] ,
    \cby_1__1__54_chany_top_out[6] ,
    \cby_1__1__54_chany_top_out[7] ,
    \cby_1__1__54_chany_top_out[8] ,
    \cby_1__1__54_chany_top_out[9] ,
    \cby_1__1__54_chany_top_out[10] ,
    \cby_1__1__54_chany_top_out[11] ,
    \cby_1__1__54_chany_top_out[12] ,
    \cby_1__1__54_chany_top_out[13] ,
    \cby_1__1__54_chany_top_out[14] ,
    \cby_1__1__54_chany_top_out[15] ,
    \cby_1__1__54_chany_top_out[16] ,
    \cby_1__1__54_chany_top_out[17] ,
    \cby_1__1__54_chany_top_out[18] ,
    \cby_1__1__54_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__1__48_chany_bottom_out[0] ,
    \sb_1__1__48_chany_bottom_out[1] ,
    \sb_1__1__48_chany_bottom_out[2] ,
    \sb_1__1__48_chany_bottom_out[3] ,
    \sb_1__1__48_chany_bottom_out[4] ,
    \sb_1__1__48_chany_bottom_out[5] ,
    \sb_1__1__48_chany_bottom_out[6] ,
    \sb_1__1__48_chany_bottom_out[7] ,
    \sb_1__1__48_chany_bottom_out[8] ,
    \sb_1__1__48_chany_bottom_out[9] ,
    \sb_1__1__48_chany_bottom_out[10] ,
    \sb_1__1__48_chany_bottom_out[11] ,
    \sb_1__1__48_chany_bottom_out[12] ,
    \sb_1__1__48_chany_bottom_out[13] ,
    \sb_1__1__48_chany_bottom_out[14] ,
    \sb_1__1__48_chany_bottom_out[15] ,
    \sb_1__1__48_chany_bottom_out[16] ,
    \sb_1__1__48_chany_bottom_out[17] ,
    \sb_1__1__48_chany_bottom_out[18] ,
    \sb_1__1__48_chany_bottom_out[19] }),
    .chany_top_in({\cby_1__1__55_chany_bottom_out[0] ,
    \cby_1__1__55_chany_bottom_out[1] ,
    \cby_1__1__55_chany_bottom_out[2] ,
    \cby_1__1__55_chany_bottom_out[3] ,
    \cby_1__1__55_chany_bottom_out[4] ,
    \cby_1__1__55_chany_bottom_out[5] ,
    \cby_1__1__55_chany_bottom_out[6] ,
    \cby_1__1__55_chany_bottom_out[7] ,
    \cby_1__1__55_chany_bottom_out[8] ,
    \cby_1__1__55_chany_bottom_out[9] ,
    \cby_1__1__55_chany_bottom_out[10] ,
    \cby_1__1__55_chany_bottom_out[11] ,
    \cby_1__1__55_chany_bottom_out[12] ,
    \cby_1__1__55_chany_bottom_out[13] ,
    \cby_1__1__55_chany_bottom_out[14] ,
    \cby_1__1__55_chany_bottom_out[15] ,
    \cby_1__1__55_chany_bottom_out[16] ,
    \cby_1__1__55_chany_bottom_out[17] ,
    \cby_1__1__55_chany_bottom_out[18] ,
    \cby_1__1__55_chany_bottom_out[19] }),
    .chany_top_out({\sb_1__1__48_chany_top_out[0] ,
    \sb_1__1__48_chany_top_out[1] ,
    \sb_1__1__48_chany_top_out[2] ,
    \sb_1__1__48_chany_top_out[3] ,
    \sb_1__1__48_chany_top_out[4] ,
    \sb_1__1__48_chany_top_out[5] ,
    \sb_1__1__48_chany_top_out[6] ,
    \sb_1__1__48_chany_top_out[7] ,
    \sb_1__1__48_chany_top_out[8] ,
    \sb_1__1__48_chany_top_out[9] ,
    \sb_1__1__48_chany_top_out[10] ,
    \sb_1__1__48_chany_top_out[11] ,
    \sb_1__1__48_chany_top_out[12] ,
    \sb_1__1__48_chany_top_out[13] ,
    \sb_1__1__48_chany_top_out[14] ,
    \sb_1__1__48_chany_top_out[15] ,
    \sb_1__1__48_chany_top_out[16] ,
    \sb_1__1__48_chany_top_out[17] ,
    \sb_1__1__48_chany_top_out[18] ,
    \sb_1__1__48_chany_top_out[19] }));
 sb_1__2_ sb_7__8_ (.bottom_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_upper),
    .ccff_head(grid_io_top_7_ccff_tail),
    .ccff_tail(sb_1__8__6_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[198] ),
    .right_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_upper),
    .right_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_upper),
    .right_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_upper),
    .right_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_upper),
    .right_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_upper),
    .right_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_upper),
    .right_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_upper),
    .right_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_upper),
    .right_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_upper),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__6_chanx_right_out[0] ,
    \cbx_1__8__6_chanx_right_out[1] ,
    \cbx_1__8__6_chanx_right_out[2] ,
    \cbx_1__8__6_chanx_right_out[3] ,
    \cbx_1__8__6_chanx_right_out[4] ,
    \cbx_1__8__6_chanx_right_out[5] ,
    \cbx_1__8__6_chanx_right_out[6] ,
    \cbx_1__8__6_chanx_right_out[7] ,
    \cbx_1__8__6_chanx_right_out[8] ,
    \cbx_1__8__6_chanx_right_out[9] ,
    \cbx_1__8__6_chanx_right_out[10] ,
    \cbx_1__8__6_chanx_right_out[11] ,
    \cbx_1__8__6_chanx_right_out[12] ,
    \cbx_1__8__6_chanx_right_out[13] ,
    \cbx_1__8__6_chanx_right_out[14] ,
    \cbx_1__8__6_chanx_right_out[15] ,
    \cbx_1__8__6_chanx_right_out[16] ,
    \cbx_1__8__6_chanx_right_out[17] ,
    \cbx_1__8__6_chanx_right_out[18] ,
    \cbx_1__8__6_chanx_right_out[19] }),
    .chanx_left_out({\sb_1__8__6_chanx_left_out[0] ,
    \sb_1__8__6_chanx_left_out[1] ,
    \sb_1__8__6_chanx_left_out[2] ,
    \sb_1__8__6_chanx_left_out[3] ,
    \sb_1__8__6_chanx_left_out[4] ,
    \sb_1__8__6_chanx_left_out[5] ,
    \sb_1__8__6_chanx_left_out[6] ,
    \sb_1__8__6_chanx_left_out[7] ,
    \sb_1__8__6_chanx_left_out[8] ,
    \sb_1__8__6_chanx_left_out[9] ,
    \sb_1__8__6_chanx_left_out[10] ,
    \sb_1__8__6_chanx_left_out[11] ,
    \sb_1__8__6_chanx_left_out[12] ,
    \sb_1__8__6_chanx_left_out[13] ,
    \sb_1__8__6_chanx_left_out[14] ,
    \sb_1__8__6_chanx_left_out[15] ,
    \sb_1__8__6_chanx_left_out[16] ,
    \sb_1__8__6_chanx_left_out[17] ,
    \sb_1__8__6_chanx_left_out[18] ,
    \sb_1__8__6_chanx_left_out[19] }),
    .chanx_right_in({\cbx_1__8__7_chanx_left_out[0] ,
    \cbx_1__8__7_chanx_left_out[1] ,
    \cbx_1__8__7_chanx_left_out[2] ,
    \cbx_1__8__7_chanx_left_out[3] ,
    \cbx_1__8__7_chanx_left_out[4] ,
    \cbx_1__8__7_chanx_left_out[5] ,
    \cbx_1__8__7_chanx_left_out[6] ,
    \cbx_1__8__7_chanx_left_out[7] ,
    \cbx_1__8__7_chanx_left_out[8] ,
    \cbx_1__8__7_chanx_left_out[9] ,
    \cbx_1__8__7_chanx_left_out[10] ,
    \cbx_1__8__7_chanx_left_out[11] ,
    \cbx_1__8__7_chanx_left_out[12] ,
    \cbx_1__8__7_chanx_left_out[13] ,
    \cbx_1__8__7_chanx_left_out[14] ,
    \cbx_1__8__7_chanx_left_out[15] ,
    \cbx_1__8__7_chanx_left_out[16] ,
    \cbx_1__8__7_chanx_left_out[17] ,
    \cbx_1__8__7_chanx_left_out[18] ,
    \cbx_1__8__7_chanx_left_out[19] }),
    .chanx_right_out({\sb_1__8__6_chanx_right_out[0] ,
    \sb_1__8__6_chanx_right_out[1] ,
    \sb_1__8__6_chanx_right_out[2] ,
    \sb_1__8__6_chanx_right_out[3] ,
    \sb_1__8__6_chanx_right_out[4] ,
    \sb_1__8__6_chanx_right_out[5] ,
    \sb_1__8__6_chanx_right_out[6] ,
    \sb_1__8__6_chanx_right_out[7] ,
    \sb_1__8__6_chanx_right_out[8] ,
    \sb_1__8__6_chanx_right_out[9] ,
    \sb_1__8__6_chanx_right_out[10] ,
    \sb_1__8__6_chanx_right_out[11] ,
    \sb_1__8__6_chanx_right_out[12] ,
    \sb_1__8__6_chanx_right_out[13] ,
    \sb_1__8__6_chanx_right_out[14] ,
    \sb_1__8__6_chanx_right_out[15] ,
    \sb_1__8__6_chanx_right_out[16] ,
    \sb_1__8__6_chanx_right_out[17] ,
    \sb_1__8__6_chanx_right_out[18] ,
    \sb_1__8__6_chanx_right_out[19] }),
    .chany_bottom_in({\cby_1__1__55_chany_top_out[0] ,
    \cby_1__1__55_chany_top_out[1] ,
    \cby_1__1__55_chany_top_out[2] ,
    \cby_1__1__55_chany_top_out[3] ,
    \cby_1__1__55_chany_top_out[4] ,
    \cby_1__1__55_chany_top_out[5] ,
    \cby_1__1__55_chany_top_out[6] ,
    \cby_1__1__55_chany_top_out[7] ,
    \cby_1__1__55_chany_top_out[8] ,
    \cby_1__1__55_chany_top_out[9] ,
    \cby_1__1__55_chany_top_out[10] ,
    \cby_1__1__55_chany_top_out[11] ,
    \cby_1__1__55_chany_top_out[12] ,
    \cby_1__1__55_chany_top_out[13] ,
    \cby_1__1__55_chany_top_out[14] ,
    \cby_1__1__55_chany_top_out[15] ,
    \cby_1__1__55_chany_top_out[16] ,
    \cby_1__1__55_chany_top_out[17] ,
    \cby_1__1__55_chany_top_out[18] ,
    \cby_1__1__55_chany_top_out[19] }),
    .chany_bottom_out({\sb_1__8__6_chany_bottom_out[0] ,
    \sb_1__8__6_chany_bottom_out[1] ,
    \sb_1__8__6_chany_bottom_out[2] ,
    \sb_1__8__6_chany_bottom_out[3] ,
    \sb_1__8__6_chany_bottom_out[4] ,
    \sb_1__8__6_chany_bottom_out[5] ,
    \sb_1__8__6_chany_bottom_out[6] ,
    \sb_1__8__6_chany_bottom_out[7] ,
    \sb_1__8__6_chany_bottom_out[8] ,
    \sb_1__8__6_chany_bottom_out[9] ,
    \sb_1__8__6_chany_bottom_out[10] ,
    \sb_1__8__6_chany_bottom_out[11] ,
    \sb_1__8__6_chany_bottom_out[12] ,
    \sb_1__8__6_chany_bottom_out[13] ,
    \sb_1__8__6_chany_bottom_out[14] ,
    \sb_1__8__6_chany_bottom_out[15] ,
    \sb_1__8__6_chany_bottom_out[16] ,
    \sb_1__8__6_chany_bottom_out[17] ,
    \sb_1__8__6_chany_bottom_out[18] ,
    \sb_1__8__6_chany_bottom_out[19] }));
 sb_2__0_ sb_8__0_ (.ccff_head(grid_io_right_7_ccff_tail),
    .ccff_tail(sb_8__0__0_ccff_tail),
    .left_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_lower),
    .left_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_lower),
    .left_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_lower),
    .left_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_lower),
    .left_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_lower),
    .left_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_lower),
    .left_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_lower),
    .left_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_lower),
    .left_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[201] ),
    .top_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__0__7_chanx_right_out[0] ,
    \cbx_1__0__7_chanx_right_out[1] ,
    \cbx_1__0__7_chanx_right_out[2] ,
    \cbx_1__0__7_chanx_right_out[3] ,
    \cbx_1__0__7_chanx_right_out[4] ,
    \cbx_1__0__7_chanx_right_out[5] ,
    \cbx_1__0__7_chanx_right_out[6] ,
    \cbx_1__0__7_chanx_right_out[7] ,
    \cbx_1__0__7_chanx_right_out[8] ,
    \cbx_1__0__7_chanx_right_out[9] ,
    \cbx_1__0__7_chanx_right_out[10] ,
    \cbx_1__0__7_chanx_right_out[11] ,
    \cbx_1__0__7_chanx_right_out[12] ,
    \cbx_1__0__7_chanx_right_out[13] ,
    \cbx_1__0__7_chanx_right_out[14] ,
    \cbx_1__0__7_chanx_right_out[15] ,
    \cbx_1__0__7_chanx_right_out[16] ,
    \cbx_1__0__7_chanx_right_out[17] ,
    \cbx_1__0__7_chanx_right_out[18] ,
    \cbx_1__0__7_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__0__0_chanx_left_out[0] ,
    \sb_8__0__0_chanx_left_out[1] ,
    \sb_8__0__0_chanx_left_out[2] ,
    \sb_8__0__0_chanx_left_out[3] ,
    \sb_8__0__0_chanx_left_out[4] ,
    \sb_8__0__0_chanx_left_out[5] ,
    \sb_8__0__0_chanx_left_out[6] ,
    \sb_8__0__0_chanx_left_out[7] ,
    \sb_8__0__0_chanx_left_out[8] ,
    \sb_8__0__0_chanx_left_out[9] ,
    \sb_8__0__0_chanx_left_out[10] ,
    \sb_8__0__0_chanx_left_out[11] ,
    \sb_8__0__0_chanx_left_out[12] ,
    \sb_8__0__0_chanx_left_out[13] ,
    \sb_8__0__0_chanx_left_out[14] ,
    \sb_8__0__0_chanx_left_out[15] ,
    \sb_8__0__0_chanx_left_out[16] ,
    \sb_8__0__0_chanx_left_out[17] ,
    \sb_8__0__0_chanx_left_out[18] ,
    \sb_8__0__0_chanx_left_out[19] }),
    .chany_top_in({\cby_8__1__0_chany_bottom_out[0] ,
    \cby_8__1__0_chany_bottom_out[1] ,
    \cby_8__1__0_chany_bottom_out[2] ,
    \cby_8__1__0_chany_bottom_out[3] ,
    \cby_8__1__0_chany_bottom_out[4] ,
    \cby_8__1__0_chany_bottom_out[5] ,
    \cby_8__1__0_chany_bottom_out[6] ,
    \cby_8__1__0_chany_bottom_out[7] ,
    \cby_8__1__0_chany_bottom_out[8] ,
    \cby_8__1__0_chany_bottom_out[9] ,
    \cby_8__1__0_chany_bottom_out[10] ,
    \cby_8__1__0_chany_bottom_out[11] ,
    \cby_8__1__0_chany_bottom_out[12] ,
    \cby_8__1__0_chany_bottom_out[13] ,
    \cby_8__1__0_chany_bottom_out[14] ,
    \cby_8__1__0_chany_bottom_out[15] ,
    \cby_8__1__0_chany_bottom_out[16] ,
    \cby_8__1__0_chany_bottom_out[17] ,
    \cby_8__1__0_chany_bottom_out[18] ,
    \cby_8__1__0_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__0__0_chany_top_out[0] ,
    \sb_8__0__0_chany_top_out[1] ,
    \sb_8__0__0_chany_top_out[2] ,
    \sb_8__0__0_chany_top_out[3] ,
    \sb_8__0__0_chany_top_out[4] ,
    \sb_8__0__0_chany_top_out[5] ,
    \sb_8__0__0_chany_top_out[6] ,
    \sb_8__0__0_chany_top_out[7] ,
    \sb_8__0__0_chany_top_out[8] ,
    \sb_8__0__0_chany_top_out[9] ,
    \sb_8__0__0_chany_top_out[10] ,
    \sb_8__0__0_chany_top_out[11] ,
    \sb_8__0__0_chany_top_out[12] ,
    \sb_8__0__0_chany_top_out[13] ,
    \sb_8__0__0_chany_top_out[14] ,
    \sb_8__0__0_chany_top_out[15] ,
    \sb_8__0__0_chany_top_out[16] ,
    \sb_8__0__0_chany_top_out[17] ,
    \sb_8__0__0_chany_top_out[18] ,
    \sb_8__0__0_chany_top_out[19] }));
 sb_2__1_ sb_8__1_ (.bottom_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_right_6_ccff_tail),
    .ccff_tail(sb_8__1__0_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[204] ),
    .top_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__49_chanx_right_out[0] ,
    \cbx_1__1__49_chanx_right_out[1] ,
    \cbx_1__1__49_chanx_right_out[2] ,
    \cbx_1__1__49_chanx_right_out[3] ,
    \cbx_1__1__49_chanx_right_out[4] ,
    \cbx_1__1__49_chanx_right_out[5] ,
    \cbx_1__1__49_chanx_right_out[6] ,
    \cbx_1__1__49_chanx_right_out[7] ,
    \cbx_1__1__49_chanx_right_out[8] ,
    \cbx_1__1__49_chanx_right_out[9] ,
    \cbx_1__1__49_chanx_right_out[10] ,
    \cbx_1__1__49_chanx_right_out[11] ,
    \cbx_1__1__49_chanx_right_out[12] ,
    \cbx_1__1__49_chanx_right_out[13] ,
    \cbx_1__1__49_chanx_right_out[14] ,
    \cbx_1__1__49_chanx_right_out[15] ,
    \cbx_1__1__49_chanx_right_out[16] ,
    \cbx_1__1__49_chanx_right_out[17] ,
    \cbx_1__1__49_chanx_right_out[18] ,
    \cbx_1__1__49_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__1__0_chanx_left_out[0] ,
    \sb_8__1__0_chanx_left_out[1] ,
    \sb_8__1__0_chanx_left_out[2] ,
    \sb_8__1__0_chanx_left_out[3] ,
    \sb_8__1__0_chanx_left_out[4] ,
    \sb_8__1__0_chanx_left_out[5] ,
    \sb_8__1__0_chanx_left_out[6] ,
    \sb_8__1__0_chanx_left_out[7] ,
    \sb_8__1__0_chanx_left_out[8] ,
    \sb_8__1__0_chanx_left_out[9] ,
    \sb_8__1__0_chanx_left_out[10] ,
    \sb_8__1__0_chanx_left_out[11] ,
    \sb_8__1__0_chanx_left_out[12] ,
    \sb_8__1__0_chanx_left_out[13] ,
    \sb_8__1__0_chanx_left_out[14] ,
    \sb_8__1__0_chanx_left_out[15] ,
    \sb_8__1__0_chanx_left_out[16] ,
    \sb_8__1__0_chanx_left_out[17] ,
    \sb_8__1__0_chanx_left_out[18] ,
    \sb_8__1__0_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__0_chany_top_out[0] ,
    \cby_8__1__0_chany_top_out[1] ,
    \cby_8__1__0_chany_top_out[2] ,
    \cby_8__1__0_chany_top_out[3] ,
    \cby_8__1__0_chany_top_out[4] ,
    \cby_8__1__0_chany_top_out[5] ,
    \cby_8__1__0_chany_top_out[6] ,
    \cby_8__1__0_chany_top_out[7] ,
    \cby_8__1__0_chany_top_out[8] ,
    \cby_8__1__0_chany_top_out[9] ,
    \cby_8__1__0_chany_top_out[10] ,
    \cby_8__1__0_chany_top_out[11] ,
    \cby_8__1__0_chany_top_out[12] ,
    \cby_8__1__0_chany_top_out[13] ,
    \cby_8__1__0_chany_top_out[14] ,
    \cby_8__1__0_chany_top_out[15] ,
    \cby_8__1__0_chany_top_out[16] ,
    \cby_8__1__0_chany_top_out[17] ,
    \cby_8__1__0_chany_top_out[18] ,
    \cby_8__1__0_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__1__0_chany_bottom_out[0] ,
    \sb_8__1__0_chany_bottom_out[1] ,
    \sb_8__1__0_chany_bottom_out[2] ,
    \sb_8__1__0_chany_bottom_out[3] ,
    \sb_8__1__0_chany_bottom_out[4] ,
    \sb_8__1__0_chany_bottom_out[5] ,
    \sb_8__1__0_chany_bottom_out[6] ,
    \sb_8__1__0_chany_bottom_out[7] ,
    \sb_8__1__0_chany_bottom_out[8] ,
    \sb_8__1__0_chany_bottom_out[9] ,
    \sb_8__1__0_chany_bottom_out[10] ,
    \sb_8__1__0_chany_bottom_out[11] ,
    \sb_8__1__0_chany_bottom_out[12] ,
    \sb_8__1__0_chany_bottom_out[13] ,
    \sb_8__1__0_chany_bottom_out[14] ,
    \sb_8__1__0_chany_bottom_out[15] ,
    \sb_8__1__0_chany_bottom_out[16] ,
    \sb_8__1__0_chany_bottom_out[17] ,
    \sb_8__1__0_chany_bottom_out[18] ,
    \sb_8__1__0_chany_bottom_out[19] }),
    .chany_top_in({\cby_8__1__1_chany_bottom_out[0] ,
    \cby_8__1__1_chany_bottom_out[1] ,
    \cby_8__1__1_chany_bottom_out[2] ,
    \cby_8__1__1_chany_bottom_out[3] ,
    \cby_8__1__1_chany_bottom_out[4] ,
    \cby_8__1__1_chany_bottom_out[5] ,
    \cby_8__1__1_chany_bottom_out[6] ,
    \cby_8__1__1_chany_bottom_out[7] ,
    \cby_8__1__1_chany_bottom_out[8] ,
    \cby_8__1__1_chany_bottom_out[9] ,
    \cby_8__1__1_chany_bottom_out[10] ,
    \cby_8__1__1_chany_bottom_out[11] ,
    \cby_8__1__1_chany_bottom_out[12] ,
    \cby_8__1__1_chany_bottom_out[13] ,
    \cby_8__1__1_chany_bottom_out[14] ,
    \cby_8__1__1_chany_bottom_out[15] ,
    \cby_8__1__1_chany_bottom_out[16] ,
    \cby_8__1__1_chany_bottom_out[17] ,
    \cby_8__1__1_chany_bottom_out[18] ,
    \cby_8__1__1_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__1__0_chany_top_out[0] ,
    \sb_8__1__0_chany_top_out[1] ,
    \sb_8__1__0_chany_top_out[2] ,
    \sb_8__1__0_chany_top_out[3] ,
    \sb_8__1__0_chany_top_out[4] ,
    \sb_8__1__0_chany_top_out[5] ,
    \sb_8__1__0_chany_top_out[6] ,
    \sb_8__1__0_chany_top_out[7] ,
    \sb_8__1__0_chany_top_out[8] ,
    \sb_8__1__0_chany_top_out[9] ,
    \sb_8__1__0_chany_top_out[10] ,
    \sb_8__1__0_chany_top_out[11] ,
    \sb_8__1__0_chany_top_out[12] ,
    \sb_8__1__0_chany_top_out[13] ,
    \sb_8__1__0_chany_top_out[14] ,
    \sb_8__1__0_chany_top_out[15] ,
    \sb_8__1__0_chany_top_out[16] ,
    \sb_8__1__0_chany_top_out[17] ,
    \sb_8__1__0_chany_top_out[18] ,
    \sb_8__1__0_chany_top_out[19] }));
 sb_2__1_ sb_8__2_ (.bottom_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_right_5_ccff_tail),
    .ccff_tail(sb_8__1__1_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[207] ),
    .top_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__50_chanx_right_out[0] ,
    \cbx_1__1__50_chanx_right_out[1] ,
    \cbx_1__1__50_chanx_right_out[2] ,
    \cbx_1__1__50_chanx_right_out[3] ,
    \cbx_1__1__50_chanx_right_out[4] ,
    \cbx_1__1__50_chanx_right_out[5] ,
    \cbx_1__1__50_chanx_right_out[6] ,
    \cbx_1__1__50_chanx_right_out[7] ,
    \cbx_1__1__50_chanx_right_out[8] ,
    \cbx_1__1__50_chanx_right_out[9] ,
    \cbx_1__1__50_chanx_right_out[10] ,
    \cbx_1__1__50_chanx_right_out[11] ,
    \cbx_1__1__50_chanx_right_out[12] ,
    \cbx_1__1__50_chanx_right_out[13] ,
    \cbx_1__1__50_chanx_right_out[14] ,
    \cbx_1__1__50_chanx_right_out[15] ,
    \cbx_1__1__50_chanx_right_out[16] ,
    \cbx_1__1__50_chanx_right_out[17] ,
    \cbx_1__1__50_chanx_right_out[18] ,
    \cbx_1__1__50_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__1__1_chanx_left_out[0] ,
    \sb_8__1__1_chanx_left_out[1] ,
    \sb_8__1__1_chanx_left_out[2] ,
    \sb_8__1__1_chanx_left_out[3] ,
    \sb_8__1__1_chanx_left_out[4] ,
    \sb_8__1__1_chanx_left_out[5] ,
    \sb_8__1__1_chanx_left_out[6] ,
    \sb_8__1__1_chanx_left_out[7] ,
    \sb_8__1__1_chanx_left_out[8] ,
    \sb_8__1__1_chanx_left_out[9] ,
    \sb_8__1__1_chanx_left_out[10] ,
    \sb_8__1__1_chanx_left_out[11] ,
    \sb_8__1__1_chanx_left_out[12] ,
    \sb_8__1__1_chanx_left_out[13] ,
    \sb_8__1__1_chanx_left_out[14] ,
    \sb_8__1__1_chanx_left_out[15] ,
    \sb_8__1__1_chanx_left_out[16] ,
    \sb_8__1__1_chanx_left_out[17] ,
    \sb_8__1__1_chanx_left_out[18] ,
    \sb_8__1__1_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__1_chany_top_out[0] ,
    \cby_8__1__1_chany_top_out[1] ,
    \cby_8__1__1_chany_top_out[2] ,
    \cby_8__1__1_chany_top_out[3] ,
    \cby_8__1__1_chany_top_out[4] ,
    \cby_8__1__1_chany_top_out[5] ,
    \cby_8__1__1_chany_top_out[6] ,
    \cby_8__1__1_chany_top_out[7] ,
    \cby_8__1__1_chany_top_out[8] ,
    \cby_8__1__1_chany_top_out[9] ,
    \cby_8__1__1_chany_top_out[10] ,
    \cby_8__1__1_chany_top_out[11] ,
    \cby_8__1__1_chany_top_out[12] ,
    \cby_8__1__1_chany_top_out[13] ,
    \cby_8__1__1_chany_top_out[14] ,
    \cby_8__1__1_chany_top_out[15] ,
    \cby_8__1__1_chany_top_out[16] ,
    \cby_8__1__1_chany_top_out[17] ,
    \cby_8__1__1_chany_top_out[18] ,
    \cby_8__1__1_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__1__1_chany_bottom_out[0] ,
    \sb_8__1__1_chany_bottom_out[1] ,
    \sb_8__1__1_chany_bottom_out[2] ,
    \sb_8__1__1_chany_bottom_out[3] ,
    \sb_8__1__1_chany_bottom_out[4] ,
    \sb_8__1__1_chany_bottom_out[5] ,
    \sb_8__1__1_chany_bottom_out[6] ,
    \sb_8__1__1_chany_bottom_out[7] ,
    \sb_8__1__1_chany_bottom_out[8] ,
    \sb_8__1__1_chany_bottom_out[9] ,
    \sb_8__1__1_chany_bottom_out[10] ,
    \sb_8__1__1_chany_bottom_out[11] ,
    \sb_8__1__1_chany_bottom_out[12] ,
    \sb_8__1__1_chany_bottom_out[13] ,
    \sb_8__1__1_chany_bottom_out[14] ,
    \sb_8__1__1_chany_bottom_out[15] ,
    \sb_8__1__1_chany_bottom_out[16] ,
    \sb_8__1__1_chany_bottom_out[17] ,
    \sb_8__1__1_chany_bottom_out[18] ,
    \sb_8__1__1_chany_bottom_out[19] }),
    .chany_top_in({\cby_8__1__2_chany_bottom_out[0] ,
    \cby_8__1__2_chany_bottom_out[1] ,
    \cby_8__1__2_chany_bottom_out[2] ,
    \cby_8__1__2_chany_bottom_out[3] ,
    \cby_8__1__2_chany_bottom_out[4] ,
    \cby_8__1__2_chany_bottom_out[5] ,
    \cby_8__1__2_chany_bottom_out[6] ,
    \cby_8__1__2_chany_bottom_out[7] ,
    \cby_8__1__2_chany_bottom_out[8] ,
    \cby_8__1__2_chany_bottom_out[9] ,
    \cby_8__1__2_chany_bottom_out[10] ,
    \cby_8__1__2_chany_bottom_out[11] ,
    \cby_8__1__2_chany_bottom_out[12] ,
    \cby_8__1__2_chany_bottom_out[13] ,
    \cby_8__1__2_chany_bottom_out[14] ,
    \cby_8__1__2_chany_bottom_out[15] ,
    \cby_8__1__2_chany_bottom_out[16] ,
    \cby_8__1__2_chany_bottom_out[17] ,
    \cby_8__1__2_chany_bottom_out[18] ,
    \cby_8__1__2_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__1__1_chany_top_out[0] ,
    \sb_8__1__1_chany_top_out[1] ,
    \sb_8__1__1_chany_top_out[2] ,
    \sb_8__1__1_chany_top_out[3] ,
    \sb_8__1__1_chany_top_out[4] ,
    \sb_8__1__1_chany_top_out[5] ,
    \sb_8__1__1_chany_top_out[6] ,
    \sb_8__1__1_chany_top_out[7] ,
    \sb_8__1__1_chany_top_out[8] ,
    \sb_8__1__1_chany_top_out[9] ,
    \sb_8__1__1_chany_top_out[10] ,
    \sb_8__1__1_chany_top_out[11] ,
    \sb_8__1__1_chany_top_out[12] ,
    \sb_8__1__1_chany_top_out[13] ,
    \sb_8__1__1_chany_top_out[14] ,
    \sb_8__1__1_chany_top_out[15] ,
    \sb_8__1__1_chany_top_out[16] ,
    \sb_8__1__1_chany_top_out[17] ,
    \sb_8__1__1_chany_top_out[18] ,
    \sb_8__1__1_chany_top_out[19] }));
 sb_2__1_ sb_8__3_ (.bottom_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_right_4_ccff_tail),
    .ccff_tail(sb_8__1__2_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[210] ),
    .top_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__51_chanx_right_out[0] ,
    \cbx_1__1__51_chanx_right_out[1] ,
    \cbx_1__1__51_chanx_right_out[2] ,
    \cbx_1__1__51_chanx_right_out[3] ,
    \cbx_1__1__51_chanx_right_out[4] ,
    \cbx_1__1__51_chanx_right_out[5] ,
    \cbx_1__1__51_chanx_right_out[6] ,
    \cbx_1__1__51_chanx_right_out[7] ,
    \cbx_1__1__51_chanx_right_out[8] ,
    \cbx_1__1__51_chanx_right_out[9] ,
    \cbx_1__1__51_chanx_right_out[10] ,
    \cbx_1__1__51_chanx_right_out[11] ,
    \cbx_1__1__51_chanx_right_out[12] ,
    \cbx_1__1__51_chanx_right_out[13] ,
    \cbx_1__1__51_chanx_right_out[14] ,
    \cbx_1__1__51_chanx_right_out[15] ,
    \cbx_1__1__51_chanx_right_out[16] ,
    \cbx_1__1__51_chanx_right_out[17] ,
    \cbx_1__1__51_chanx_right_out[18] ,
    \cbx_1__1__51_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__1__2_chanx_left_out[0] ,
    \sb_8__1__2_chanx_left_out[1] ,
    \sb_8__1__2_chanx_left_out[2] ,
    \sb_8__1__2_chanx_left_out[3] ,
    \sb_8__1__2_chanx_left_out[4] ,
    \sb_8__1__2_chanx_left_out[5] ,
    \sb_8__1__2_chanx_left_out[6] ,
    \sb_8__1__2_chanx_left_out[7] ,
    \sb_8__1__2_chanx_left_out[8] ,
    \sb_8__1__2_chanx_left_out[9] ,
    \sb_8__1__2_chanx_left_out[10] ,
    \sb_8__1__2_chanx_left_out[11] ,
    \sb_8__1__2_chanx_left_out[12] ,
    \sb_8__1__2_chanx_left_out[13] ,
    \sb_8__1__2_chanx_left_out[14] ,
    \sb_8__1__2_chanx_left_out[15] ,
    \sb_8__1__2_chanx_left_out[16] ,
    \sb_8__1__2_chanx_left_out[17] ,
    \sb_8__1__2_chanx_left_out[18] ,
    \sb_8__1__2_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__2_chany_top_out[0] ,
    \cby_8__1__2_chany_top_out[1] ,
    \cby_8__1__2_chany_top_out[2] ,
    \cby_8__1__2_chany_top_out[3] ,
    \cby_8__1__2_chany_top_out[4] ,
    \cby_8__1__2_chany_top_out[5] ,
    \cby_8__1__2_chany_top_out[6] ,
    \cby_8__1__2_chany_top_out[7] ,
    \cby_8__1__2_chany_top_out[8] ,
    \cby_8__1__2_chany_top_out[9] ,
    \cby_8__1__2_chany_top_out[10] ,
    \cby_8__1__2_chany_top_out[11] ,
    \cby_8__1__2_chany_top_out[12] ,
    \cby_8__1__2_chany_top_out[13] ,
    \cby_8__1__2_chany_top_out[14] ,
    \cby_8__1__2_chany_top_out[15] ,
    \cby_8__1__2_chany_top_out[16] ,
    \cby_8__1__2_chany_top_out[17] ,
    \cby_8__1__2_chany_top_out[18] ,
    \cby_8__1__2_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__1__2_chany_bottom_out[0] ,
    \sb_8__1__2_chany_bottom_out[1] ,
    \sb_8__1__2_chany_bottom_out[2] ,
    \sb_8__1__2_chany_bottom_out[3] ,
    \sb_8__1__2_chany_bottom_out[4] ,
    \sb_8__1__2_chany_bottom_out[5] ,
    \sb_8__1__2_chany_bottom_out[6] ,
    \sb_8__1__2_chany_bottom_out[7] ,
    \sb_8__1__2_chany_bottom_out[8] ,
    \sb_8__1__2_chany_bottom_out[9] ,
    \sb_8__1__2_chany_bottom_out[10] ,
    \sb_8__1__2_chany_bottom_out[11] ,
    \sb_8__1__2_chany_bottom_out[12] ,
    \sb_8__1__2_chany_bottom_out[13] ,
    \sb_8__1__2_chany_bottom_out[14] ,
    \sb_8__1__2_chany_bottom_out[15] ,
    \sb_8__1__2_chany_bottom_out[16] ,
    \sb_8__1__2_chany_bottom_out[17] ,
    \sb_8__1__2_chany_bottom_out[18] ,
    \sb_8__1__2_chany_bottom_out[19] }),
    .chany_top_in({\cby_8__1__3_chany_bottom_out[0] ,
    \cby_8__1__3_chany_bottom_out[1] ,
    \cby_8__1__3_chany_bottom_out[2] ,
    \cby_8__1__3_chany_bottom_out[3] ,
    \cby_8__1__3_chany_bottom_out[4] ,
    \cby_8__1__3_chany_bottom_out[5] ,
    \cby_8__1__3_chany_bottom_out[6] ,
    \cby_8__1__3_chany_bottom_out[7] ,
    \cby_8__1__3_chany_bottom_out[8] ,
    \cby_8__1__3_chany_bottom_out[9] ,
    \cby_8__1__3_chany_bottom_out[10] ,
    \cby_8__1__3_chany_bottom_out[11] ,
    \cby_8__1__3_chany_bottom_out[12] ,
    \cby_8__1__3_chany_bottom_out[13] ,
    \cby_8__1__3_chany_bottom_out[14] ,
    \cby_8__1__3_chany_bottom_out[15] ,
    \cby_8__1__3_chany_bottom_out[16] ,
    \cby_8__1__3_chany_bottom_out[17] ,
    \cby_8__1__3_chany_bottom_out[18] ,
    \cby_8__1__3_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__1__2_chany_top_out[0] ,
    \sb_8__1__2_chany_top_out[1] ,
    \sb_8__1__2_chany_top_out[2] ,
    \sb_8__1__2_chany_top_out[3] ,
    \sb_8__1__2_chany_top_out[4] ,
    \sb_8__1__2_chany_top_out[5] ,
    \sb_8__1__2_chany_top_out[6] ,
    \sb_8__1__2_chany_top_out[7] ,
    \sb_8__1__2_chany_top_out[8] ,
    \sb_8__1__2_chany_top_out[9] ,
    \sb_8__1__2_chany_top_out[10] ,
    \sb_8__1__2_chany_top_out[11] ,
    \sb_8__1__2_chany_top_out[12] ,
    \sb_8__1__2_chany_top_out[13] ,
    \sb_8__1__2_chany_top_out[14] ,
    \sb_8__1__2_chany_top_out[15] ,
    \sb_8__1__2_chany_top_out[16] ,
    \sb_8__1__2_chany_top_out[17] ,
    \sb_8__1__2_chany_top_out[18] ,
    \sb_8__1__2_chany_top_out[19] }));
 sb_2__1_ sb_8__4_ (.bottom_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_right_3_ccff_tail),
    .ccff_tail(sb_8__1__3_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[213] ),
    .top_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__52_chanx_right_out[0] ,
    \cbx_1__1__52_chanx_right_out[1] ,
    \cbx_1__1__52_chanx_right_out[2] ,
    \cbx_1__1__52_chanx_right_out[3] ,
    \cbx_1__1__52_chanx_right_out[4] ,
    \cbx_1__1__52_chanx_right_out[5] ,
    \cbx_1__1__52_chanx_right_out[6] ,
    \cbx_1__1__52_chanx_right_out[7] ,
    \cbx_1__1__52_chanx_right_out[8] ,
    \cbx_1__1__52_chanx_right_out[9] ,
    \cbx_1__1__52_chanx_right_out[10] ,
    \cbx_1__1__52_chanx_right_out[11] ,
    \cbx_1__1__52_chanx_right_out[12] ,
    \cbx_1__1__52_chanx_right_out[13] ,
    \cbx_1__1__52_chanx_right_out[14] ,
    \cbx_1__1__52_chanx_right_out[15] ,
    \cbx_1__1__52_chanx_right_out[16] ,
    \cbx_1__1__52_chanx_right_out[17] ,
    \cbx_1__1__52_chanx_right_out[18] ,
    \cbx_1__1__52_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__1__3_chanx_left_out[0] ,
    \sb_8__1__3_chanx_left_out[1] ,
    \sb_8__1__3_chanx_left_out[2] ,
    \sb_8__1__3_chanx_left_out[3] ,
    \sb_8__1__3_chanx_left_out[4] ,
    \sb_8__1__3_chanx_left_out[5] ,
    \sb_8__1__3_chanx_left_out[6] ,
    \sb_8__1__3_chanx_left_out[7] ,
    \sb_8__1__3_chanx_left_out[8] ,
    \sb_8__1__3_chanx_left_out[9] ,
    \sb_8__1__3_chanx_left_out[10] ,
    \sb_8__1__3_chanx_left_out[11] ,
    \sb_8__1__3_chanx_left_out[12] ,
    \sb_8__1__3_chanx_left_out[13] ,
    \sb_8__1__3_chanx_left_out[14] ,
    \sb_8__1__3_chanx_left_out[15] ,
    \sb_8__1__3_chanx_left_out[16] ,
    \sb_8__1__3_chanx_left_out[17] ,
    \sb_8__1__3_chanx_left_out[18] ,
    \sb_8__1__3_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__3_chany_top_out[0] ,
    \cby_8__1__3_chany_top_out[1] ,
    \cby_8__1__3_chany_top_out[2] ,
    \cby_8__1__3_chany_top_out[3] ,
    \cby_8__1__3_chany_top_out[4] ,
    \cby_8__1__3_chany_top_out[5] ,
    \cby_8__1__3_chany_top_out[6] ,
    \cby_8__1__3_chany_top_out[7] ,
    \cby_8__1__3_chany_top_out[8] ,
    \cby_8__1__3_chany_top_out[9] ,
    \cby_8__1__3_chany_top_out[10] ,
    \cby_8__1__3_chany_top_out[11] ,
    \cby_8__1__3_chany_top_out[12] ,
    \cby_8__1__3_chany_top_out[13] ,
    \cby_8__1__3_chany_top_out[14] ,
    \cby_8__1__3_chany_top_out[15] ,
    \cby_8__1__3_chany_top_out[16] ,
    \cby_8__1__3_chany_top_out[17] ,
    \cby_8__1__3_chany_top_out[18] ,
    \cby_8__1__3_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__1__3_chany_bottom_out[0] ,
    \sb_8__1__3_chany_bottom_out[1] ,
    \sb_8__1__3_chany_bottom_out[2] ,
    \sb_8__1__3_chany_bottom_out[3] ,
    \sb_8__1__3_chany_bottom_out[4] ,
    \sb_8__1__3_chany_bottom_out[5] ,
    \sb_8__1__3_chany_bottom_out[6] ,
    \sb_8__1__3_chany_bottom_out[7] ,
    \sb_8__1__3_chany_bottom_out[8] ,
    \sb_8__1__3_chany_bottom_out[9] ,
    \sb_8__1__3_chany_bottom_out[10] ,
    \sb_8__1__3_chany_bottom_out[11] ,
    \sb_8__1__3_chany_bottom_out[12] ,
    \sb_8__1__3_chany_bottom_out[13] ,
    \sb_8__1__3_chany_bottom_out[14] ,
    \sb_8__1__3_chany_bottom_out[15] ,
    \sb_8__1__3_chany_bottom_out[16] ,
    \sb_8__1__3_chany_bottom_out[17] ,
    \sb_8__1__3_chany_bottom_out[18] ,
    \sb_8__1__3_chany_bottom_out[19] }),
    .chany_top_in({\cby_8__1__4_chany_bottom_out[0] ,
    \cby_8__1__4_chany_bottom_out[1] ,
    \cby_8__1__4_chany_bottom_out[2] ,
    \cby_8__1__4_chany_bottom_out[3] ,
    \cby_8__1__4_chany_bottom_out[4] ,
    \cby_8__1__4_chany_bottom_out[5] ,
    \cby_8__1__4_chany_bottom_out[6] ,
    \cby_8__1__4_chany_bottom_out[7] ,
    \cby_8__1__4_chany_bottom_out[8] ,
    \cby_8__1__4_chany_bottom_out[9] ,
    \cby_8__1__4_chany_bottom_out[10] ,
    \cby_8__1__4_chany_bottom_out[11] ,
    \cby_8__1__4_chany_bottom_out[12] ,
    \cby_8__1__4_chany_bottom_out[13] ,
    \cby_8__1__4_chany_bottom_out[14] ,
    \cby_8__1__4_chany_bottom_out[15] ,
    \cby_8__1__4_chany_bottom_out[16] ,
    \cby_8__1__4_chany_bottom_out[17] ,
    \cby_8__1__4_chany_bottom_out[18] ,
    \cby_8__1__4_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__1__3_chany_top_out[0] ,
    \sb_8__1__3_chany_top_out[1] ,
    \sb_8__1__3_chany_top_out[2] ,
    \sb_8__1__3_chany_top_out[3] ,
    \sb_8__1__3_chany_top_out[4] ,
    \sb_8__1__3_chany_top_out[5] ,
    \sb_8__1__3_chany_top_out[6] ,
    \sb_8__1__3_chany_top_out[7] ,
    \sb_8__1__3_chany_top_out[8] ,
    \sb_8__1__3_chany_top_out[9] ,
    \sb_8__1__3_chany_top_out[10] ,
    \sb_8__1__3_chany_top_out[11] ,
    \sb_8__1__3_chany_top_out[12] ,
    \sb_8__1__3_chany_top_out[13] ,
    \sb_8__1__3_chany_top_out[14] ,
    \sb_8__1__3_chany_top_out[15] ,
    \sb_8__1__3_chany_top_out[16] ,
    \sb_8__1__3_chany_top_out[17] ,
    \sb_8__1__3_chany_top_out[18] ,
    \sb_8__1__3_chany_top_out[19] }));
 sb_2__1_ sb_8__5_ (.bottom_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_right_2_ccff_tail),
    .ccff_tail(sb_8__1__4_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[216] ),
    .top_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__53_chanx_right_out[0] ,
    \cbx_1__1__53_chanx_right_out[1] ,
    \cbx_1__1__53_chanx_right_out[2] ,
    \cbx_1__1__53_chanx_right_out[3] ,
    \cbx_1__1__53_chanx_right_out[4] ,
    \cbx_1__1__53_chanx_right_out[5] ,
    \cbx_1__1__53_chanx_right_out[6] ,
    \cbx_1__1__53_chanx_right_out[7] ,
    \cbx_1__1__53_chanx_right_out[8] ,
    \cbx_1__1__53_chanx_right_out[9] ,
    \cbx_1__1__53_chanx_right_out[10] ,
    \cbx_1__1__53_chanx_right_out[11] ,
    \cbx_1__1__53_chanx_right_out[12] ,
    \cbx_1__1__53_chanx_right_out[13] ,
    \cbx_1__1__53_chanx_right_out[14] ,
    \cbx_1__1__53_chanx_right_out[15] ,
    \cbx_1__1__53_chanx_right_out[16] ,
    \cbx_1__1__53_chanx_right_out[17] ,
    \cbx_1__1__53_chanx_right_out[18] ,
    \cbx_1__1__53_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__1__4_chanx_left_out[0] ,
    \sb_8__1__4_chanx_left_out[1] ,
    \sb_8__1__4_chanx_left_out[2] ,
    \sb_8__1__4_chanx_left_out[3] ,
    \sb_8__1__4_chanx_left_out[4] ,
    \sb_8__1__4_chanx_left_out[5] ,
    \sb_8__1__4_chanx_left_out[6] ,
    \sb_8__1__4_chanx_left_out[7] ,
    \sb_8__1__4_chanx_left_out[8] ,
    \sb_8__1__4_chanx_left_out[9] ,
    \sb_8__1__4_chanx_left_out[10] ,
    \sb_8__1__4_chanx_left_out[11] ,
    \sb_8__1__4_chanx_left_out[12] ,
    \sb_8__1__4_chanx_left_out[13] ,
    \sb_8__1__4_chanx_left_out[14] ,
    \sb_8__1__4_chanx_left_out[15] ,
    \sb_8__1__4_chanx_left_out[16] ,
    \sb_8__1__4_chanx_left_out[17] ,
    \sb_8__1__4_chanx_left_out[18] ,
    \sb_8__1__4_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__4_chany_top_out[0] ,
    \cby_8__1__4_chany_top_out[1] ,
    \cby_8__1__4_chany_top_out[2] ,
    \cby_8__1__4_chany_top_out[3] ,
    \cby_8__1__4_chany_top_out[4] ,
    \cby_8__1__4_chany_top_out[5] ,
    \cby_8__1__4_chany_top_out[6] ,
    \cby_8__1__4_chany_top_out[7] ,
    \cby_8__1__4_chany_top_out[8] ,
    \cby_8__1__4_chany_top_out[9] ,
    \cby_8__1__4_chany_top_out[10] ,
    \cby_8__1__4_chany_top_out[11] ,
    \cby_8__1__4_chany_top_out[12] ,
    \cby_8__1__4_chany_top_out[13] ,
    \cby_8__1__4_chany_top_out[14] ,
    \cby_8__1__4_chany_top_out[15] ,
    \cby_8__1__4_chany_top_out[16] ,
    \cby_8__1__4_chany_top_out[17] ,
    \cby_8__1__4_chany_top_out[18] ,
    \cby_8__1__4_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__1__4_chany_bottom_out[0] ,
    \sb_8__1__4_chany_bottom_out[1] ,
    \sb_8__1__4_chany_bottom_out[2] ,
    \sb_8__1__4_chany_bottom_out[3] ,
    \sb_8__1__4_chany_bottom_out[4] ,
    \sb_8__1__4_chany_bottom_out[5] ,
    \sb_8__1__4_chany_bottom_out[6] ,
    \sb_8__1__4_chany_bottom_out[7] ,
    \sb_8__1__4_chany_bottom_out[8] ,
    \sb_8__1__4_chany_bottom_out[9] ,
    \sb_8__1__4_chany_bottom_out[10] ,
    \sb_8__1__4_chany_bottom_out[11] ,
    \sb_8__1__4_chany_bottom_out[12] ,
    \sb_8__1__4_chany_bottom_out[13] ,
    \sb_8__1__4_chany_bottom_out[14] ,
    \sb_8__1__4_chany_bottom_out[15] ,
    \sb_8__1__4_chany_bottom_out[16] ,
    \sb_8__1__4_chany_bottom_out[17] ,
    \sb_8__1__4_chany_bottom_out[18] ,
    \sb_8__1__4_chany_bottom_out[19] }),
    .chany_top_in({\cby_8__1__5_chany_bottom_out[0] ,
    \cby_8__1__5_chany_bottom_out[1] ,
    \cby_8__1__5_chany_bottom_out[2] ,
    \cby_8__1__5_chany_bottom_out[3] ,
    \cby_8__1__5_chany_bottom_out[4] ,
    \cby_8__1__5_chany_bottom_out[5] ,
    \cby_8__1__5_chany_bottom_out[6] ,
    \cby_8__1__5_chany_bottom_out[7] ,
    \cby_8__1__5_chany_bottom_out[8] ,
    \cby_8__1__5_chany_bottom_out[9] ,
    \cby_8__1__5_chany_bottom_out[10] ,
    \cby_8__1__5_chany_bottom_out[11] ,
    \cby_8__1__5_chany_bottom_out[12] ,
    \cby_8__1__5_chany_bottom_out[13] ,
    \cby_8__1__5_chany_bottom_out[14] ,
    \cby_8__1__5_chany_bottom_out[15] ,
    \cby_8__1__5_chany_bottom_out[16] ,
    \cby_8__1__5_chany_bottom_out[17] ,
    \cby_8__1__5_chany_bottom_out[18] ,
    \cby_8__1__5_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__1__4_chany_top_out[0] ,
    \sb_8__1__4_chany_top_out[1] ,
    \sb_8__1__4_chany_top_out[2] ,
    \sb_8__1__4_chany_top_out[3] ,
    \sb_8__1__4_chany_top_out[4] ,
    \sb_8__1__4_chany_top_out[5] ,
    \sb_8__1__4_chany_top_out[6] ,
    \sb_8__1__4_chany_top_out[7] ,
    \sb_8__1__4_chany_top_out[8] ,
    \sb_8__1__4_chany_top_out[9] ,
    \sb_8__1__4_chany_top_out[10] ,
    \sb_8__1__4_chany_top_out[11] ,
    \sb_8__1__4_chany_top_out[12] ,
    \sb_8__1__4_chany_top_out[13] ,
    \sb_8__1__4_chany_top_out[14] ,
    \sb_8__1__4_chany_top_out[15] ,
    \sb_8__1__4_chany_top_out[16] ,
    \sb_8__1__4_chany_top_out[17] ,
    \sb_8__1__4_chany_top_out[18] ,
    \sb_8__1__4_chany_top_out[19] }));
 sb_2__1_ sb_8__6_ (.bottom_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_right_1_ccff_tail),
    .ccff_tail(sb_8__1__5_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[219] ),
    .top_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__54_chanx_right_out[0] ,
    \cbx_1__1__54_chanx_right_out[1] ,
    \cbx_1__1__54_chanx_right_out[2] ,
    \cbx_1__1__54_chanx_right_out[3] ,
    \cbx_1__1__54_chanx_right_out[4] ,
    \cbx_1__1__54_chanx_right_out[5] ,
    \cbx_1__1__54_chanx_right_out[6] ,
    \cbx_1__1__54_chanx_right_out[7] ,
    \cbx_1__1__54_chanx_right_out[8] ,
    \cbx_1__1__54_chanx_right_out[9] ,
    \cbx_1__1__54_chanx_right_out[10] ,
    \cbx_1__1__54_chanx_right_out[11] ,
    \cbx_1__1__54_chanx_right_out[12] ,
    \cbx_1__1__54_chanx_right_out[13] ,
    \cbx_1__1__54_chanx_right_out[14] ,
    \cbx_1__1__54_chanx_right_out[15] ,
    \cbx_1__1__54_chanx_right_out[16] ,
    \cbx_1__1__54_chanx_right_out[17] ,
    \cbx_1__1__54_chanx_right_out[18] ,
    \cbx_1__1__54_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__1__5_chanx_left_out[0] ,
    \sb_8__1__5_chanx_left_out[1] ,
    \sb_8__1__5_chanx_left_out[2] ,
    \sb_8__1__5_chanx_left_out[3] ,
    \sb_8__1__5_chanx_left_out[4] ,
    \sb_8__1__5_chanx_left_out[5] ,
    \sb_8__1__5_chanx_left_out[6] ,
    \sb_8__1__5_chanx_left_out[7] ,
    \sb_8__1__5_chanx_left_out[8] ,
    \sb_8__1__5_chanx_left_out[9] ,
    \sb_8__1__5_chanx_left_out[10] ,
    \sb_8__1__5_chanx_left_out[11] ,
    \sb_8__1__5_chanx_left_out[12] ,
    \sb_8__1__5_chanx_left_out[13] ,
    \sb_8__1__5_chanx_left_out[14] ,
    \sb_8__1__5_chanx_left_out[15] ,
    \sb_8__1__5_chanx_left_out[16] ,
    \sb_8__1__5_chanx_left_out[17] ,
    \sb_8__1__5_chanx_left_out[18] ,
    \sb_8__1__5_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__5_chany_top_out[0] ,
    \cby_8__1__5_chany_top_out[1] ,
    \cby_8__1__5_chany_top_out[2] ,
    \cby_8__1__5_chany_top_out[3] ,
    \cby_8__1__5_chany_top_out[4] ,
    \cby_8__1__5_chany_top_out[5] ,
    \cby_8__1__5_chany_top_out[6] ,
    \cby_8__1__5_chany_top_out[7] ,
    \cby_8__1__5_chany_top_out[8] ,
    \cby_8__1__5_chany_top_out[9] ,
    \cby_8__1__5_chany_top_out[10] ,
    \cby_8__1__5_chany_top_out[11] ,
    \cby_8__1__5_chany_top_out[12] ,
    \cby_8__1__5_chany_top_out[13] ,
    \cby_8__1__5_chany_top_out[14] ,
    \cby_8__1__5_chany_top_out[15] ,
    \cby_8__1__5_chany_top_out[16] ,
    \cby_8__1__5_chany_top_out[17] ,
    \cby_8__1__5_chany_top_out[18] ,
    \cby_8__1__5_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__1__5_chany_bottom_out[0] ,
    \sb_8__1__5_chany_bottom_out[1] ,
    \sb_8__1__5_chany_bottom_out[2] ,
    \sb_8__1__5_chany_bottom_out[3] ,
    \sb_8__1__5_chany_bottom_out[4] ,
    \sb_8__1__5_chany_bottom_out[5] ,
    \sb_8__1__5_chany_bottom_out[6] ,
    \sb_8__1__5_chany_bottom_out[7] ,
    \sb_8__1__5_chany_bottom_out[8] ,
    \sb_8__1__5_chany_bottom_out[9] ,
    \sb_8__1__5_chany_bottom_out[10] ,
    \sb_8__1__5_chany_bottom_out[11] ,
    \sb_8__1__5_chany_bottom_out[12] ,
    \sb_8__1__5_chany_bottom_out[13] ,
    \sb_8__1__5_chany_bottom_out[14] ,
    \sb_8__1__5_chany_bottom_out[15] ,
    \sb_8__1__5_chany_bottom_out[16] ,
    \sb_8__1__5_chany_bottom_out[17] ,
    \sb_8__1__5_chany_bottom_out[18] ,
    \sb_8__1__5_chany_bottom_out[19] }),
    .chany_top_in({\cby_8__1__6_chany_bottom_out[0] ,
    \cby_8__1__6_chany_bottom_out[1] ,
    \cby_8__1__6_chany_bottom_out[2] ,
    \cby_8__1__6_chany_bottom_out[3] ,
    \cby_8__1__6_chany_bottom_out[4] ,
    \cby_8__1__6_chany_bottom_out[5] ,
    \cby_8__1__6_chany_bottom_out[6] ,
    \cby_8__1__6_chany_bottom_out[7] ,
    \cby_8__1__6_chany_bottom_out[8] ,
    \cby_8__1__6_chany_bottom_out[9] ,
    \cby_8__1__6_chany_bottom_out[10] ,
    \cby_8__1__6_chany_bottom_out[11] ,
    \cby_8__1__6_chany_bottom_out[12] ,
    \cby_8__1__6_chany_bottom_out[13] ,
    \cby_8__1__6_chany_bottom_out[14] ,
    \cby_8__1__6_chany_bottom_out[15] ,
    \cby_8__1__6_chany_bottom_out[16] ,
    \cby_8__1__6_chany_bottom_out[17] ,
    \cby_8__1__6_chany_bottom_out[18] ,
    \cby_8__1__6_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__1__5_chany_top_out[0] ,
    \sb_8__1__5_chany_top_out[1] ,
    \sb_8__1__5_chany_top_out[2] ,
    \sb_8__1__5_chany_top_out[3] ,
    \sb_8__1__5_chany_top_out[4] ,
    \sb_8__1__5_chany_top_out[5] ,
    \sb_8__1__5_chany_top_out[6] ,
    \sb_8__1__5_chany_top_out[7] ,
    \sb_8__1__5_chany_top_out[8] ,
    \sb_8__1__5_chany_top_out[9] ,
    \sb_8__1__5_chany_top_out[10] ,
    \sb_8__1__5_chany_top_out[11] ,
    \sb_8__1__5_chany_top_out[12] ,
    \sb_8__1__5_chany_top_out[13] ,
    \sb_8__1__5_chany_top_out[14] ,
    \sb_8__1__5_chany_top_out[15] ,
    \sb_8__1__5_chany_top_out[16] ,
    \sb_8__1__5_chany_top_out[17] ,
    \sb_8__1__5_chany_top_out[18] ,
    \sb_8__1__5_chany_top_out[19] }));
 sb_2__1_ sb_8__7_ (.bottom_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_upper),
    .ccff_head(grid_io_right_0_ccff_tail),
    .ccff_tail(sb_8__1__6_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_lower),
    .prog_clk_0_N_in(\prog_clk_0_wires[222] ),
    .top_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_lower),
    .top_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_lower),
    .top_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_lower),
    .top_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_lower),
    .top_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_lower),
    .top_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_lower),
    .top_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_lower),
    .top_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_lower),
    .top_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_lower),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__1__55_chanx_right_out[0] ,
    \cbx_1__1__55_chanx_right_out[1] ,
    \cbx_1__1__55_chanx_right_out[2] ,
    \cbx_1__1__55_chanx_right_out[3] ,
    \cbx_1__1__55_chanx_right_out[4] ,
    \cbx_1__1__55_chanx_right_out[5] ,
    \cbx_1__1__55_chanx_right_out[6] ,
    \cbx_1__1__55_chanx_right_out[7] ,
    \cbx_1__1__55_chanx_right_out[8] ,
    \cbx_1__1__55_chanx_right_out[9] ,
    \cbx_1__1__55_chanx_right_out[10] ,
    \cbx_1__1__55_chanx_right_out[11] ,
    \cbx_1__1__55_chanx_right_out[12] ,
    \cbx_1__1__55_chanx_right_out[13] ,
    \cbx_1__1__55_chanx_right_out[14] ,
    \cbx_1__1__55_chanx_right_out[15] ,
    \cbx_1__1__55_chanx_right_out[16] ,
    \cbx_1__1__55_chanx_right_out[17] ,
    \cbx_1__1__55_chanx_right_out[18] ,
    \cbx_1__1__55_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__1__6_chanx_left_out[0] ,
    \sb_8__1__6_chanx_left_out[1] ,
    \sb_8__1__6_chanx_left_out[2] ,
    \sb_8__1__6_chanx_left_out[3] ,
    \sb_8__1__6_chanx_left_out[4] ,
    \sb_8__1__6_chanx_left_out[5] ,
    \sb_8__1__6_chanx_left_out[6] ,
    \sb_8__1__6_chanx_left_out[7] ,
    \sb_8__1__6_chanx_left_out[8] ,
    \sb_8__1__6_chanx_left_out[9] ,
    \sb_8__1__6_chanx_left_out[10] ,
    \sb_8__1__6_chanx_left_out[11] ,
    \sb_8__1__6_chanx_left_out[12] ,
    \sb_8__1__6_chanx_left_out[13] ,
    \sb_8__1__6_chanx_left_out[14] ,
    \sb_8__1__6_chanx_left_out[15] ,
    \sb_8__1__6_chanx_left_out[16] ,
    \sb_8__1__6_chanx_left_out[17] ,
    \sb_8__1__6_chanx_left_out[18] ,
    \sb_8__1__6_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__6_chany_top_out[0] ,
    \cby_8__1__6_chany_top_out[1] ,
    \cby_8__1__6_chany_top_out[2] ,
    \cby_8__1__6_chany_top_out[3] ,
    \cby_8__1__6_chany_top_out[4] ,
    \cby_8__1__6_chany_top_out[5] ,
    \cby_8__1__6_chany_top_out[6] ,
    \cby_8__1__6_chany_top_out[7] ,
    \cby_8__1__6_chany_top_out[8] ,
    \cby_8__1__6_chany_top_out[9] ,
    \cby_8__1__6_chany_top_out[10] ,
    \cby_8__1__6_chany_top_out[11] ,
    \cby_8__1__6_chany_top_out[12] ,
    \cby_8__1__6_chany_top_out[13] ,
    \cby_8__1__6_chany_top_out[14] ,
    \cby_8__1__6_chany_top_out[15] ,
    \cby_8__1__6_chany_top_out[16] ,
    \cby_8__1__6_chany_top_out[17] ,
    \cby_8__1__6_chany_top_out[18] ,
    \cby_8__1__6_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__1__6_chany_bottom_out[0] ,
    \sb_8__1__6_chany_bottom_out[1] ,
    \sb_8__1__6_chany_bottom_out[2] ,
    \sb_8__1__6_chany_bottom_out[3] ,
    \sb_8__1__6_chany_bottom_out[4] ,
    \sb_8__1__6_chany_bottom_out[5] ,
    \sb_8__1__6_chany_bottom_out[6] ,
    \sb_8__1__6_chany_bottom_out[7] ,
    \sb_8__1__6_chany_bottom_out[8] ,
    \sb_8__1__6_chany_bottom_out[9] ,
    \sb_8__1__6_chany_bottom_out[10] ,
    \sb_8__1__6_chany_bottom_out[11] ,
    \sb_8__1__6_chany_bottom_out[12] ,
    \sb_8__1__6_chany_bottom_out[13] ,
    \sb_8__1__6_chany_bottom_out[14] ,
    \sb_8__1__6_chany_bottom_out[15] ,
    \sb_8__1__6_chany_bottom_out[16] ,
    \sb_8__1__6_chany_bottom_out[17] ,
    \sb_8__1__6_chany_bottom_out[18] ,
    \sb_8__1__6_chany_bottom_out[19] }),
    .chany_top_in({\cby_8__1__7_chany_bottom_out[0] ,
    \cby_8__1__7_chany_bottom_out[1] ,
    \cby_8__1__7_chany_bottom_out[2] ,
    \cby_8__1__7_chany_bottom_out[3] ,
    \cby_8__1__7_chany_bottom_out[4] ,
    \cby_8__1__7_chany_bottom_out[5] ,
    \cby_8__1__7_chany_bottom_out[6] ,
    \cby_8__1__7_chany_bottom_out[7] ,
    \cby_8__1__7_chany_bottom_out[8] ,
    \cby_8__1__7_chany_bottom_out[9] ,
    \cby_8__1__7_chany_bottom_out[10] ,
    \cby_8__1__7_chany_bottom_out[11] ,
    \cby_8__1__7_chany_bottom_out[12] ,
    \cby_8__1__7_chany_bottom_out[13] ,
    \cby_8__1__7_chany_bottom_out[14] ,
    \cby_8__1__7_chany_bottom_out[15] ,
    \cby_8__1__7_chany_bottom_out[16] ,
    \cby_8__1__7_chany_bottom_out[17] ,
    \cby_8__1__7_chany_bottom_out[18] ,
    \cby_8__1__7_chany_bottom_out[19] }),
    .chany_top_out({\sb_8__1__6_chany_top_out[0] ,
    \sb_8__1__6_chany_top_out[1] ,
    \sb_8__1__6_chany_top_out[2] ,
    \sb_8__1__6_chany_top_out[3] ,
    \sb_8__1__6_chany_top_out[4] ,
    \sb_8__1__6_chany_top_out[5] ,
    \sb_8__1__6_chany_top_out[6] ,
    \sb_8__1__6_chany_top_out[7] ,
    \sb_8__1__6_chany_top_out[8] ,
    \sb_8__1__6_chany_top_out[9] ,
    \sb_8__1__6_chany_top_out[10] ,
    \sb_8__1__6_chany_top_out[11] ,
    \sb_8__1__6_chany_top_out[12] ,
    \sb_8__1__6_chany_top_out[13] ,
    \sb_8__1__6_chany_top_out[14] ,
    \sb_8__1__6_chany_top_out[15] ,
    \sb_8__1__6_chany_top_out[16] ,
    \sb_8__1__6_chany_top_out[17] ,
    \sb_8__1__6_chany_top_out[18] ,
    \sb_8__1__6_chany_top_out[19] }));
 sb_2__2_ sb_8__8_ (.SC_IN_BOT(\scff_Wires[147] ),
    .SC_OUT_BOT(sc_tail),
    .bottom_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_upper),
    .bottom_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_upper),
    .bottom_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_upper),
    .bottom_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_upper),
    .bottom_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_upper),
    .bottom_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_upper),
    .bottom_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_upper),
    .bottom_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_upper),
    .bottom_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_upper),
    .ccff_head(ccff_head),
    .ccff_tail(sb_8__8__0_ccff_tail),
    .left_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_lower),
    .left_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_lower),
    .left_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_lower),
    .left_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_lower),
    .left_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_lower),
    .left_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_lower),
    .left_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_lower),
    .left_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_lower),
    .left_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_lower),
    .prog_clk_0_S_in(\prog_clk_0_wires[224] ),
    .VPWR(VPWR),
    .VGND(VGND),
    .chanx_left_in({\cbx_1__8__7_chanx_right_out[0] ,
    \cbx_1__8__7_chanx_right_out[1] ,
    \cbx_1__8__7_chanx_right_out[2] ,
    \cbx_1__8__7_chanx_right_out[3] ,
    \cbx_1__8__7_chanx_right_out[4] ,
    \cbx_1__8__7_chanx_right_out[5] ,
    \cbx_1__8__7_chanx_right_out[6] ,
    \cbx_1__8__7_chanx_right_out[7] ,
    \cbx_1__8__7_chanx_right_out[8] ,
    \cbx_1__8__7_chanx_right_out[9] ,
    \cbx_1__8__7_chanx_right_out[10] ,
    \cbx_1__8__7_chanx_right_out[11] ,
    \cbx_1__8__7_chanx_right_out[12] ,
    \cbx_1__8__7_chanx_right_out[13] ,
    \cbx_1__8__7_chanx_right_out[14] ,
    \cbx_1__8__7_chanx_right_out[15] ,
    \cbx_1__8__7_chanx_right_out[16] ,
    \cbx_1__8__7_chanx_right_out[17] ,
    \cbx_1__8__7_chanx_right_out[18] ,
    \cbx_1__8__7_chanx_right_out[19] }),
    .chanx_left_out({\sb_8__8__0_chanx_left_out[0] ,
    \sb_8__8__0_chanx_left_out[1] ,
    \sb_8__8__0_chanx_left_out[2] ,
    \sb_8__8__0_chanx_left_out[3] ,
    \sb_8__8__0_chanx_left_out[4] ,
    \sb_8__8__0_chanx_left_out[5] ,
    \sb_8__8__0_chanx_left_out[6] ,
    \sb_8__8__0_chanx_left_out[7] ,
    \sb_8__8__0_chanx_left_out[8] ,
    \sb_8__8__0_chanx_left_out[9] ,
    \sb_8__8__0_chanx_left_out[10] ,
    \sb_8__8__0_chanx_left_out[11] ,
    \sb_8__8__0_chanx_left_out[12] ,
    \sb_8__8__0_chanx_left_out[13] ,
    \sb_8__8__0_chanx_left_out[14] ,
    \sb_8__8__0_chanx_left_out[15] ,
    \sb_8__8__0_chanx_left_out[16] ,
    \sb_8__8__0_chanx_left_out[17] ,
    \sb_8__8__0_chanx_left_out[18] ,
    \sb_8__8__0_chanx_left_out[19] }),
    .chany_bottom_in({\cby_8__1__7_chany_top_out[0] ,
    \cby_8__1__7_chany_top_out[1] ,
    \cby_8__1__7_chany_top_out[2] ,
    \cby_8__1__7_chany_top_out[3] ,
    \cby_8__1__7_chany_top_out[4] ,
    \cby_8__1__7_chany_top_out[5] ,
    \cby_8__1__7_chany_top_out[6] ,
    \cby_8__1__7_chany_top_out[7] ,
    \cby_8__1__7_chany_top_out[8] ,
    \cby_8__1__7_chany_top_out[9] ,
    \cby_8__1__7_chany_top_out[10] ,
    \cby_8__1__7_chany_top_out[11] ,
    \cby_8__1__7_chany_top_out[12] ,
    \cby_8__1__7_chany_top_out[13] ,
    \cby_8__1__7_chany_top_out[14] ,
    \cby_8__1__7_chany_top_out[15] ,
    \cby_8__1__7_chany_top_out[16] ,
    \cby_8__1__7_chany_top_out[17] ,
    \cby_8__1__7_chany_top_out[18] ,
    \cby_8__1__7_chany_top_out[19] }),
    .chany_bottom_out({\sb_8__8__0_chany_bottom_out[0] ,
    \sb_8__8__0_chany_bottom_out[1] ,
    \sb_8__8__0_chany_bottom_out[2] ,
    \sb_8__8__0_chany_bottom_out[3] ,
    \sb_8__8__0_chany_bottom_out[4] ,
    \sb_8__8__0_chany_bottom_out[5] ,
    \sb_8__8__0_chany_bottom_out[6] ,
    \sb_8__8__0_chany_bottom_out[7] ,
    \sb_8__8__0_chany_bottom_out[8] ,
    \sb_8__8__0_chany_bottom_out[9] ,
    \sb_8__8__0_chany_bottom_out[10] ,
    \sb_8__8__0_chany_bottom_out[11] ,
    \sb_8__8__0_chany_bottom_out[12] ,
    \sb_8__8__0_chany_bottom_out[13] ,
    \sb_8__8__0_chany_bottom_out[14] ,
    \sb_8__8__0_chany_bottom_out[15] ,
    \sb_8__8__0_chany_bottom_out[16] ,
    \sb_8__8__0_chany_bottom_out[17] ,
    \sb_8__8__0_chany_bottom_out[18] ,
    \sb_8__8__0_chany_bottom_out[19] }));
 tie_array tie_array (.VPWR(VPWR),
    .VGND(VGND),
    .x({\logic_zero_tie[7] ,
    \logic_zero_tie[6] ,
    \logic_zero_tie[5] ,
    \logic_zero_tie[4] ,
    \logic_zero_tie[3] ,
    \logic_zero_tie[2] ,
    \logic_zero_tie[1] ,
    \logic_zero_tie[0] }));
endmodule
