VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2475.000 BY 2715.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -12.760 -3.720 -7.960 2718.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 -3.720 2487.560 1.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2713.480 2487.560 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2482.760 -3.720 2487.560 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.920 -3.720 13.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 -3.720 70.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 171.365 70.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 477.540 70.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 792.540 70.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 1107.540 70.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 1422.540 70.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 1737.540 70.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 2052.540 70.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 2367.540 70.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 2682.540 70.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 -3.720 127.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 171.365 127.120 199.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 475.085 127.120 514.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 790.085 127.120 829.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 1105.085 127.120 1144.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 1420.085 127.120 1459.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 1735.085 127.120 1774.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 2050.085 127.120 2089.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 2365.085 127.120 2402.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 2618.885 127.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.920 -3.720 184.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 -3.720 241.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 454.005 241.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 769.005 241.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 1084.005 241.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 1399.005 241.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 1714.005 241.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 2029.005 241.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 2344.005 241.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 2656.285 241.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 -3.720 298.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 165.245 298.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 454.005 298.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 769.005 298.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 1084.005 298.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 1399.005 298.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 1714.005 298.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 2029.005 298.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 2344.005 298.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 2656.285 298.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 -3.720 355.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 165.245 355.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 454.005 355.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 769.005 355.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 1084.005 355.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 1399.005 355.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 1714.005 355.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 2029.005 355.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 2344.005 355.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 2656.285 355.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 -3.720 412.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 162.940 412.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 477.540 412.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 792.540 412.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 1107.540 412.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 1422.540 412.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 1737.540 412.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 2052.540 412.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 2367.540 412.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 2682.540 412.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.920 -3.720 469.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 -3.720 526.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 454.005 526.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 769.005 526.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 1084.005 526.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 1399.005 526.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 1714.005 526.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 2029.005 526.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 2344.005 526.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 2656.285 526.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 -3.720 583.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 165.245 583.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 454.005 583.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 769.005 583.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 1084.005 583.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 1399.005 583.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 1714.005 583.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 2029.005 583.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 2344.005 583.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 2656.285 583.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 -3.720 640.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 165.245 640.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 454.005 640.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 769.005 640.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 1084.005 640.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 1399.005 640.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 1714.005 640.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 2029.005 640.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 2344.005 640.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 2656.285 640.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 -3.720 697.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 162.940 697.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 477.540 697.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 792.540 697.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 1107.540 697.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 1422.540 697.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 1737.540 697.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 2052.540 697.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 2367.540 697.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 2682.540 697.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.920 -3.720 754.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 -3.720 811.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 454.005 811.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 769.005 811.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 1084.005 811.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 1399.005 811.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 1714.005 811.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 2029.005 811.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 2344.005 811.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 2656.285 811.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 -3.720 868.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 165.245 868.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 454.005 868.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 769.005 868.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 1084.005 868.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 1399.005 868.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 1714.005 868.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 2029.005 868.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 2344.005 868.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 2656.285 868.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 -3.720 925.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 165.245 925.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 454.005 925.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 769.005 925.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 1084.005 925.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 1399.005 925.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 1714.005 925.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 2029.005 925.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 2344.005 925.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 2656.285 925.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 -3.720 982.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 162.940 982.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 477.540 982.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 792.540 982.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 1107.540 982.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 1422.540 982.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 1737.540 982.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 2052.540 982.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 2367.540 982.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 2682.540 982.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.920 -3.720 1039.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 -3.720 1096.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 454.005 1096.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 769.005 1096.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 1084.005 1096.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 1399.005 1096.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 1714.005 1096.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 2029.005 1096.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 2344.005 1096.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 2656.285 1096.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 -3.720 1153.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 165.245 1153.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 454.005 1153.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 769.005 1153.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 1084.005 1153.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 1399.005 1153.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 1714.005 1153.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 2029.005 1153.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 2344.005 1153.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 2656.285 1153.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 -3.720 1210.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 165.245 1210.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 454.005 1210.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 769.005 1210.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 1084.005 1210.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 1399.005 1210.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 1714.005 1210.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 2029.005 1210.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 2344.005 1210.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 2656.285 1210.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 -3.720 1267.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 162.940 1267.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 477.540 1267.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 792.540 1267.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 1107.540 1267.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 1422.540 1267.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 1737.540 1267.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 2052.540 1267.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 2367.540 1267.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 2682.540 1267.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1320.920 -3.720 1324.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 -3.720 1381.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 454.005 1381.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 769.005 1381.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 1084.005 1381.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 1399.005 1381.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 1714.005 1381.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 2029.005 1381.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 2344.005 1381.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 2656.285 1381.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 -3.720 1438.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 165.245 1438.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 454.005 1438.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 769.005 1438.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 1084.005 1438.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 1399.005 1438.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 1714.005 1438.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 2029.005 1438.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 2344.005 1438.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 2656.285 1438.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 -3.720 1495.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 165.245 1495.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 454.005 1495.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 769.005 1495.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 1084.005 1495.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 1399.005 1495.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 1714.005 1495.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 2029.005 1495.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 2344.005 1495.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 2656.285 1495.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 -3.720 1552.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 162.940 1552.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 477.540 1552.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 792.540 1552.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 1107.540 1552.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 1422.540 1552.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 1737.540 1552.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 2052.540 1552.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 2367.540 1552.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 2682.540 1552.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1605.920 -3.720 1609.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 -3.720 1666.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 454.005 1666.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 769.005 1666.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 1084.005 1666.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 1399.005 1666.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 1714.005 1666.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 2029.005 1666.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 2344.005 1666.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 2656.285 1666.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 -3.720 1723.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 165.245 1723.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 454.005 1723.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 769.005 1723.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 1084.005 1723.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 1399.005 1723.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 1714.005 1723.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 2029.005 1723.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 2344.005 1723.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 2656.285 1723.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 -3.720 1780.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 165.245 1780.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 454.005 1780.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 769.005 1780.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 1084.005 1780.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 1399.005 1780.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 1714.005 1780.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 2029.005 1780.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 2344.005 1780.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 2656.285 1780.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 -3.720 1837.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 162.940 1837.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 477.540 1837.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 792.540 1837.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 1107.540 1837.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 1422.540 1837.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 1737.540 1837.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 2052.540 1837.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 2367.540 1837.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 2682.540 1837.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1890.920 -3.720 1894.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 -3.720 1951.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 454.005 1951.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 769.005 1951.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 1084.005 1951.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 1399.005 1951.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 1714.005 1951.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 2029.005 1951.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 2344.005 1951.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 2656.285 1951.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 -3.720 2008.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 165.245 2008.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 454.005 2008.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 769.005 2008.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 1084.005 2008.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 1399.005 2008.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 1714.005 2008.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 2029.005 2008.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 2344.005 2008.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 2656.285 2008.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 -3.720 2065.120 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 165.245 2065.120 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 454.005 2065.120 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 769.005 2065.120 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 1084.005 2065.120 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 1399.005 2065.120 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 1714.005 2065.120 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 2029.005 2065.120 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 2344.005 2065.120 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 2656.285 2065.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 -3.720 2122.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 162.940 2122.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 477.540 2122.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 792.540 2122.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 1107.540 2122.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 1422.540 2122.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 1737.540 2122.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 2052.540 2122.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 2367.540 2122.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 2682.540 2122.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.920 -3.720 2179.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 -3.720 2236.120 60.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 161.165 2236.120 196.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 475.085 2236.120 511.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 790.085 2236.120 826.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 1105.085 2236.120 1141.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 1420.085 2236.120 1456.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 1735.085 2236.120 1771.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 2050.085 2236.120 2086.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 2365.085 2236.120 2406.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 2680.085 2236.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 -3.720 2293.120 60.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 161.165 2293.120 196.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 475.085 2293.120 511.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 790.085 2293.120 826.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 1105.085 2293.120 1141.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 1420.085 2293.120 1456.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 1735.085 2293.120 1771.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 2050.085 2293.120 2086.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 2365.085 2293.120 2406.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 2680.085 2293.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 -3.720 2350.120 196.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 475.085 2350.120 511.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 790.085 2350.120 826.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 1105.085 2350.120 1141.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 1420.085 2350.120 1456.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 1735.085 2350.120 1771.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 2050.085 2350.120 2086.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 2365.085 2350.120 2406.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 2680.085 2350.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 -3.720 2407.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 162.940 2407.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 477.540 2407.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 792.540 2407.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 1107.540 2407.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 1422.540 2407.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 1737.540 2407.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 2052.540 2407.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 2367.540 2407.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 2682.540 2407.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2460.920 -3.720 2464.120 2718.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 25.680 2487.560 28.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 78.180 2487.560 81.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 130.680 2487.560 133.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 183.180 2487.560 186.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 235.680 2487.560 238.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 288.180 2487.560 291.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 340.680 2487.560 343.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 393.180 2487.560 396.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 445.680 2487.560 448.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 498.180 2487.560 501.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 550.680 2487.560 553.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 603.180 2487.560 606.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 655.680 2487.560 658.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 708.180 2487.560 711.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 760.680 2487.560 763.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 813.180 2487.560 816.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 865.680 2487.560 868.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 918.180 2487.560 921.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 970.680 2487.560 973.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1023.180 2487.560 1026.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1075.680 2487.560 1078.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1128.180 2487.560 1131.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1180.680 2487.560 1183.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1233.180 2487.560 1236.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1285.680 2487.560 1288.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1338.180 2487.560 1341.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1390.680 2487.560 1393.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1443.180 2487.560 1446.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1495.680 2487.560 1498.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1548.180 2487.560 1551.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1600.680 2487.560 1603.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1653.180 2487.560 1656.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1705.680 2487.560 1708.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1758.180 2487.560 1761.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1810.680 2487.560 1813.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1863.180 2487.560 1866.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1915.680 2487.560 1918.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1968.180 2487.560 1971.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2020.680 2487.560 2023.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2073.180 2487.560 2076.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2125.680 2487.560 2128.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2178.180 2487.560 2181.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2230.680 2487.560 2233.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2283.180 2487.560 2286.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2335.680 2487.560 2338.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2388.180 2487.560 2391.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2440.680 2487.560 2443.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2493.180 2487.560 2496.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2545.680 2487.560 2548.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2598.180 2487.560 2601.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2650.680 2487.560 2653.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -5.960 3.080 -1.160 2711.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.960 3.080 2480.760 7.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.960 2706.680 2480.760 2711.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.960 3.080 2480.760 2711.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.120 -3.720 8.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.120 -3.720 65.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.120 171.365 65.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 -3.720 122.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 171.365 122.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 477.540 122.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 792.540 122.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 1107.540 122.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 1422.540 122.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 1737.540 122.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 2052.540 122.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 2367.540 122.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 2682.540 122.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 176.120 -3.720 179.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 -3.720 236.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 162.940 236.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 477.540 236.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 792.540 236.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 1107.540 236.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 1422.540 236.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 1737.540 236.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 2052.540 236.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 2367.540 236.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 2682.540 236.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 -3.720 293.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 165.245 293.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 454.005 293.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 769.005 293.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 1084.005 293.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 1399.005 293.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 1714.005 293.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 2029.005 293.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 2344.005 293.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 2656.285 293.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 -3.720 350.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 165.245 350.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 454.005 350.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 769.005 350.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 1084.005 350.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 1399.005 350.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 1714.005 350.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 2029.005 350.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 2344.005 350.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 2656.285 350.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 -3.720 407.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 454.005 407.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 769.005 407.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 1084.005 407.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 1399.005 407.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 1714.005 407.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 2029.005 407.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 2344.005 407.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 2656.285 407.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.120 -3.720 464.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 -3.720 521.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 162.940 521.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 477.540 521.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 792.540 521.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 1107.540 521.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 1422.540 521.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 1737.540 521.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 2052.540 521.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 2367.540 521.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 2682.540 521.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 -3.720 578.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 165.245 578.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 454.005 578.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 769.005 578.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 1084.005 578.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 1399.005 578.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 1714.005 578.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 2029.005 578.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 2344.005 578.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 2656.285 578.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 -3.720 635.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 165.245 635.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 454.005 635.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 769.005 635.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 1084.005 635.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 1399.005 635.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 1714.005 635.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 2029.005 635.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 2344.005 635.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 2656.285 635.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 -3.720 692.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 454.005 692.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 769.005 692.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 1084.005 692.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 1399.005 692.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 1714.005 692.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 2029.005 692.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 2344.005 692.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 2656.285 692.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.120 -3.720 749.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 -3.720 806.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 162.940 806.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 477.540 806.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 792.540 806.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 1107.540 806.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 1422.540 806.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 1737.540 806.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 2052.540 806.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 2367.540 806.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 2682.540 806.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 -3.720 863.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 165.245 863.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 454.005 863.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 769.005 863.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 1084.005 863.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 1399.005 863.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 1714.005 863.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 2029.005 863.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 2344.005 863.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 2656.285 863.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 -3.720 920.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 165.245 920.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 454.005 920.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 769.005 920.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 1084.005 920.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 1399.005 920.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 1714.005 920.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 2029.005 920.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 2344.005 920.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 2656.285 920.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 -3.720 977.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 454.005 977.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 769.005 977.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 1084.005 977.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 1399.005 977.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 1714.005 977.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 2029.005 977.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 2344.005 977.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 2656.285 977.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1031.120 -3.720 1034.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 -3.720 1091.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 162.940 1091.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 477.540 1091.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 792.540 1091.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 1107.540 1091.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 1422.540 1091.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 1737.540 1091.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 2052.540 1091.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 2367.540 1091.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 2682.540 1091.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 -3.720 1148.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 165.245 1148.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 454.005 1148.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 769.005 1148.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 1084.005 1148.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 1399.005 1148.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 1714.005 1148.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 2029.005 1148.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 2344.005 1148.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 2656.285 1148.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 -3.720 1205.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 165.245 1205.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 454.005 1205.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 769.005 1205.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 1084.005 1205.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 1399.005 1205.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 1714.005 1205.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 2029.005 1205.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 2344.005 1205.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 2656.285 1205.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 -3.720 1262.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 454.005 1262.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 769.005 1262.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 1084.005 1262.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 1399.005 1262.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 1714.005 1262.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 2029.005 1262.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 2344.005 1262.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 2656.285 1262.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1316.120 -3.720 1319.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 -3.720 1376.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 162.940 1376.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 477.540 1376.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 792.540 1376.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 1107.540 1376.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 1422.540 1376.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 1737.540 1376.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 2052.540 1376.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 2367.540 1376.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 2682.540 1376.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 -3.720 1433.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 165.245 1433.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 454.005 1433.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 769.005 1433.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 1084.005 1433.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 1399.005 1433.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 1714.005 1433.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 2029.005 1433.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 2344.005 1433.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 2656.285 1433.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 -3.720 1490.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 165.245 1490.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 454.005 1490.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 769.005 1490.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 1084.005 1490.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 1399.005 1490.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 1714.005 1490.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 2029.005 1490.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 2344.005 1490.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 2656.285 1490.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 -3.720 1547.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 454.005 1547.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 769.005 1547.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 1084.005 1547.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 1399.005 1547.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 1714.005 1547.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 2029.005 1547.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 2344.005 1547.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 2656.285 1547.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1601.120 -3.720 1604.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 -3.720 1661.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 162.940 1661.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 477.540 1661.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 792.540 1661.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 1107.540 1661.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 1422.540 1661.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 1737.540 1661.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 2052.540 1661.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 2367.540 1661.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 2682.540 1661.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 -3.720 1718.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 165.245 1718.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 454.005 1718.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 769.005 1718.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 1084.005 1718.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 1399.005 1718.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 1714.005 1718.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 2029.005 1718.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 2344.005 1718.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 2656.285 1718.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 -3.720 1775.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 165.245 1775.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 454.005 1775.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 769.005 1775.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 1084.005 1775.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 1399.005 1775.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 1714.005 1775.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 2029.005 1775.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 2344.005 1775.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 2656.285 1775.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 -3.720 1832.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 454.005 1832.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 769.005 1832.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 1084.005 1832.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 1399.005 1832.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 1714.005 1832.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 2029.005 1832.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 2344.005 1832.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 2656.285 1832.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1886.120 -3.720 1889.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 -3.720 1946.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 162.940 1946.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 477.540 1946.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 792.540 1946.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 1107.540 1946.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 1422.540 1946.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 1737.540 1946.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 2052.540 1946.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 2367.540 1946.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 2682.540 1946.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 -3.720 2003.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 165.245 2003.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 454.005 2003.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 769.005 2003.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 1084.005 2003.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 1399.005 2003.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 1714.005 2003.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 2029.005 2003.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 2344.005 2003.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 2656.285 2003.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 -3.720 2060.320 67.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 165.245 2060.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 454.005 2060.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 769.005 2060.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 1084.005 2060.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 1399.005 2060.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 1714.005 2060.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 2029.005 2060.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 2344.005 2060.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 2656.285 2060.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 -3.720 2117.320 222.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 454.005 2117.320 537.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 769.005 2117.320 852.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 1084.005 2117.320 1167.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 1399.005 2117.320 1482.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 1714.005 2117.320 1797.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 2029.005 2117.320 2112.955 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 2344.005 2117.320 2421.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 2656.285 2117.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.120 -3.720 2174.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 -3.720 2231.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 162.940 2231.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 477.540 2231.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 792.540 2231.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 1107.540 2231.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 1422.540 2231.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 1737.540 2231.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 2052.540 2231.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 2367.540 2231.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 2682.540 2231.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 -3.720 2288.320 60.675 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 161.165 2288.320 196.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 475.085 2288.320 511.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 790.085 2288.320 826.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 1105.085 2288.320 1141.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 1420.085 2288.320 1456.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 1735.085 2288.320 1771.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 2050.085 2288.320 2086.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 2365.085 2288.320 2406.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 2680.085 2288.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 -3.720 2345.320 196.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 475.085 2345.320 511.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 790.085 2345.320 826.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 1105.085 2345.320 1141.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 1420.085 2345.320 1456.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 1735.085 2345.320 1771.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 2050.085 2345.320 2086.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 2365.085 2345.320 2406.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 2680.085 2345.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 -3.720 2402.320 196.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 475.085 2402.320 511.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 790.085 2402.320 826.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 1105.085 2402.320 1141.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 1420.085 2402.320 1456.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 1735.085 2402.320 1771.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 2050.085 2402.320 2086.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 2365.085 2402.320 2406.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 2680.085 2402.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2456.120 -3.720 2459.320 2718.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 19.280 2487.560 22.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 71.780 2487.560 74.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 124.280 2487.560 127.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 176.780 2487.560 179.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 229.280 2487.560 232.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 281.780 2487.560 284.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 334.280 2487.560 337.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 386.780 2487.560 389.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 439.280 2487.560 442.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 491.780 2487.560 494.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 544.280 2487.560 547.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 596.780 2487.560 599.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 649.280 2487.560 652.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 701.780 2487.560 704.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 754.280 2487.560 757.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 806.780 2487.560 809.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 859.280 2487.560 862.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 911.780 2487.560 914.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 964.280 2487.560 967.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1016.780 2487.560 1019.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1069.280 2487.560 1072.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1121.780 2487.560 1124.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1174.280 2487.560 1177.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1226.780 2487.560 1229.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1279.280 2487.560 1282.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1331.780 2487.560 1334.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1384.280 2487.560 1387.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1436.780 2487.560 1439.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1489.280 2487.560 1492.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1541.780 2487.560 1544.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1594.280 2487.560 1597.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1646.780 2487.560 1649.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1699.280 2487.560 1702.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1751.780 2487.560 1754.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1804.280 2487.560 1807.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1856.780 2487.560 1859.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1909.280 2487.560 1912.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1961.780 2487.560 1964.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2014.280 2487.560 2017.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2066.780 2487.560 2069.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2119.280 2487.560 2122.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2171.780 2487.560 2174.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2224.280 2487.560 2227.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2276.780 2487.560 2279.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2329.280 2487.560 2332.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2381.780 2487.560 2384.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2434.280 2487.560 2437.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2486.780 2487.560 2489.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2539.280 2487.560 2542.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2591.780 2487.560 2594.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2644.280 2487.560 2647.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2696.780 2487.560 2699.980 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END clk
  PIN gfpga_pad_io_soc_dir[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 2711.000 65.230 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[0]
  PIN gfpga_pad_io_soc_dir[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END gfpga_pad_io_soc_dir[100]
  PIN gfpga_pad_io_soc_dir[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END gfpga_pad_io_soc_dir[101]
  PIN gfpga_pad_io_soc_dir[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END gfpga_pad_io_soc_dir[102]
  PIN gfpga_pad_io_soc_dir[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END gfpga_pad_io_soc_dir[103]
  PIN gfpga_pad_io_soc_dir[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END gfpga_pad_io_soc_dir[104]
  PIN gfpga_pad_io_soc_dir[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END gfpga_pad_io_soc_dir[105]
  PIN gfpga_pad_io_soc_dir[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END gfpga_pad_io_soc_dir[106]
  PIN gfpga_pad_io_soc_dir[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END gfpga_pad_io_soc_dir[107]
  PIN gfpga_pad_io_soc_dir[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END gfpga_pad_io_soc_dir[108]
  PIN gfpga_pad_io_soc_dir[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END gfpga_pad_io_soc_dir[109]
  PIN gfpga_pad_io_soc_dir[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 2711.000 763.970 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[10]
  PIN gfpga_pad_io_soc_dir[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END gfpga_pad_io_soc_dir[110]
  PIN gfpga_pad_io_soc_dir[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END gfpga_pad_io_soc_dir[111]
  PIN gfpga_pad_io_soc_dir[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END gfpga_pad_io_soc_dir[112]
  PIN gfpga_pad_io_soc_dir[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END gfpga_pad_io_soc_dir[113]
  PIN gfpga_pad_io_soc_dir[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1628.640 4.000 1629.240 ;
    END
  END gfpga_pad_io_soc_dir[114]
  PIN gfpga_pad_io_soc_dir[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END gfpga_pad_io_soc_dir[115]
  PIN gfpga_pad_io_soc_dir[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.840 4.000 1792.440 ;
    END
  END gfpga_pad_io_soc_dir[116]
  PIN gfpga_pad_io_soc_dir[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1873.440 4.000 1874.040 ;
    END
  END gfpga_pad_io_soc_dir[117]
  PIN gfpga_pad_io_soc_dir[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1955.040 4.000 1955.640 ;
    END
  END gfpga_pad_io_soc_dir[118]
  PIN gfpga_pad_io_soc_dir[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2036.640 4.000 2037.240 ;
    END
  END gfpga_pad_io_soc_dir[119]
  PIN gfpga_pad_io_soc_dir[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 2711.000 831.590 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[11]
  PIN gfpga_pad_io_soc_dir[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.240 4.000 2118.840 ;
    END
  END gfpga_pad_io_soc_dir[120]
  PIN gfpga_pad_io_soc_dir[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2199.840 4.000 2200.440 ;
    END
  END gfpga_pad_io_soc_dir[121]
  PIN gfpga_pad_io_soc_dir[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2281.440 4.000 2282.040 ;
    END
  END gfpga_pad_io_soc_dir[122]
  PIN gfpga_pad_io_soc_dir[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2363.040 4.000 2363.640 ;
    END
  END gfpga_pad_io_soc_dir[123]
  PIN gfpga_pad_io_soc_dir[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2444.640 4.000 2445.240 ;
    END
  END gfpga_pad_io_soc_dir[124]
  PIN gfpga_pad_io_soc_dir[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2526.240 4.000 2526.840 ;
    END
  END gfpga_pad_io_soc_dir[125]
  PIN gfpga_pad_io_soc_dir[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2607.840 4.000 2608.440 ;
    END
  END gfpga_pad_io_soc_dir[126]
  PIN gfpga_pad_io_soc_dir[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2689.440 4.000 2690.040 ;
    END
  END gfpga_pad_io_soc_dir[127]
  PIN gfpga_pad_io_soc_dir[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 2711.000 899.210 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[12]
  PIN gfpga_pad_io_soc_dir[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 2711.000 966.830 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[13]
  PIN gfpga_pad_io_soc_dir[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 2711.000 1034.450 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[14]
  PIN gfpga_pad_io_soc_dir[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 2711.000 1102.070 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[15]
  PIN gfpga_pad_io_soc_dir[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 2711.000 1169.690 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[16]
  PIN gfpga_pad_io_soc_dir[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 2711.000 1237.310 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[17]
  PIN gfpga_pad_io_soc_dir[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.650 2711.000 1304.930 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[18]
  PIN gfpga_pad_io_soc_dir[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.270 2711.000 1372.550 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[19]
  PIN gfpga_pad_io_soc_dir[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 2711.000 132.850 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[1]
  PIN gfpga_pad_io_soc_dir[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 2711.000 1440.170 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[20]
  PIN gfpga_pad_io_soc_dir[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 2711.000 1507.790 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[21]
  PIN gfpga_pad_io_soc_dir[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 2711.000 1575.410 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[22]
  PIN gfpga_pad_io_soc_dir[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.750 2711.000 1643.030 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[23]
  PIN gfpga_pad_io_soc_dir[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.370 2711.000 1710.650 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[24]
  PIN gfpga_pad_io_soc_dir[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.990 2711.000 1778.270 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[25]
  PIN gfpga_pad_io_soc_dir[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.610 2711.000 1845.890 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[26]
  PIN gfpga_pad_io_soc_dir[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.230 2711.000 1913.510 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[27]
  PIN gfpga_pad_io_soc_dir[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.850 2711.000 1981.130 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[28]
  PIN gfpga_pad_io_soc_dir[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.470 2711.000 2048.750 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[29]
  PIN gfpga_pad_io_soc_dir[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 2711.000 200.470 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[2]
  PIN gfpga_pad_io_soc_dir[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2116.090 2711.000 2116.370 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[30]
  PIN gfpga_pad_io_soc_dir[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.710 2711.000 2183.990 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[31]
  PIN gfpga_pad_io_soc_dir[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.330 2711.000 2251.610 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[32]
  PIN gfpga_pad_io_soc_dir[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.950 2711.000 2319.230 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[33]
  PIN gfpga_pad_io_soc_dir[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.570 2711.000 2386.850 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[34]
  PIN gfpga_pad_io_soc_dir[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.190 2711.000 2454.470 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[35]
  PIN gfpga_pad_io_soc_dir[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2603.080 2475.000 2603.680 ;
    END
  END gfpga_pad_io_soc_dir[36]
  PIN gfpga_pad_io_soc_dir[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2523.520 2475.000 2524.120 ;
    END
  END gfpga_pad_io_soc_dir[37]
  PIN gfpga_pad_io_soc_dir[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2443.960 2475.000 2444.560 ;
    END
  END gfpga_pad_io_soc_dir[38]
  PIN gfpga_pad_io_soc_dir[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2364.400 2475.000 2365.000 ;
    END
  END gfpga_pad_io_soc_dir[39]
  PIN gfpga_pad_io_soc_dir[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 2711.000 268.090 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[3]
  PIN gfpga_pad_io_soc_dir[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2284.840 2475.000 2285.440 ;
    END
  END gfpga_pad_io_soc_dir[40]
  PIN gfpga_pad_io_soc_dir[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2205.280 2475.000 2205.880 ;
    END
  END gfpga_pad_io_soc_dir[41]
  PIN gfpga_pad_io_soc_dir[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2125.720 2475.000 2126.320 ;
    END
  END gfpga_pad_io_soc_dir[42]
  PIN gfpga_pad_io_soc_dir[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2046.160 2475.000 2046.760 ;
    END
  END gfpga_pad_io_soc_dir[43]
  PIN gfpga_pad_io_soc_dir[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1966.600 2475.000 1967.200 ;
    END
  END gfpga_pad_io_soc_dir[44]
  PIN gfpga_pad_io_soc_dir[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1887.040 2475.000 1887.640 ;
    END
  END gfpga_pad_io_soc_dir[45]
  PIN gfpga_pad_io_soc_dir[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1807.480 2475.000 1808.080 ;
    END
  END gfpga_pad_io_soc_dir[46]
  PIN gfpga_pad_io_soc_dir[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1727.920 2475.000 1728.520 ;
    END
  END gfpga_pad_io_soc_dir[47]
  PIN gfpga_pad_io_soc_dir[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1648.360 2475.000 1648.960 ;
    END
  END gfpga_pad_io_soc_dir[48]
  PIN gfpga_pad_io_soc_dir[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1568.800 2475.000 1569.400 ;
    END
  END gfpga_pad_io_soc_dir[49]
  PIN gfpga_pad_io_soc_dir[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 2711.000 358.250 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[4]
  PIN gfpga_pad_io_soc_dir[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1489.240 2475.000 1489.840 ;
    END
  END gfpga_pad_io_soc_dir[50]
  PIN gfpga_pad_io_soc_dir[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1409.680 2475.000 1410.280 ;
    END
  END gfpga_pad_io_soc_dir[51]
  PIN gfpga_pad_io_soc_dir[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1330.120 2475.000 1330.720 ;
    END
  END gfpga_pad_io_soc_dir[52]
  PIN gfpga_pad_io_soc_dir[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1250.560 2475.000 1251.160 ;
    END
  END gfpga_pad_io_soc_dir[53]
  PIN gfpga_pad_io_soc_dir[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1171.000 2475.000 1171.600 ;
    END
  END gfpga_pad_io_soc_dir[54]
  PIN gfpga_pad_io_soc_dir[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1091.440 2475.000 1092.040 ;
    END
  END gfpga_pad_io_soc_dir[55]
  PIN gfpga_pad_io_soc_dir[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1011.880 2475.000 1012.480 ;
    END
  END gfpga_pad_io_soc_dir[56]
  PIN gfpga_pad_io_soc_dir[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 932.320 2475.000 932.920 ;
    END
  END gfpga_pad_io_soc_dir[57]
  PIN gfpga_pad_io_soc_dir[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 852.760 2475.000 853.360 ;
    END
  END gfpga_pad_io_soc_dir[58]
  PIN gfpga_pad_io_soc_dir[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 773.200 2475.000 773.800 ;
    END
  END gfpga_pad_io_soc_dir[59]
  PIN gfpga_pad_io_soc_dir[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 2711.000 425.870 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[5]
  PIN gfpga_pad_io_soc_dir[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 693.640 2475.000 694.240 ;
    END
  END gfpga_pad_io_soc_dir[60]
  PIN gfpga_pad_io_soc_dir[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 614.080 2475.000 614.680 ;
    END
  END gfpga_pad_io_soc_dir[61]
  PIN gfpga_pad_io_soc_dir[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 534.520 2475.000 535.120 ;
    END
  END gfpga_pad_io_soc_dir[62]
  PIN gfpga_pad_io_soc_dir[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 454.960 2475.000 455.560 ;
    END
  END gfpga_pad_io_soc_dir[63]
  PIN gfpga_pad_io_soc_dir[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 375.400 2475.000 376.000 ;
    END
  END gfpga_pad_io_soc_dir[64]
  PIN gfpga_pad_io_soc_dir[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 295.840 2475.000 296.440 ;
    END
  END gfpga_pad_io_soc_dir[65]
  PIN gfpga_pad_io_soc_dir[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 216.280 2475.000 216.880 ;
    END
  END gfpga_pad_io_soc_dir[66]
  PIN gfpga_pad_io_soc_dir[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 136.720 2475.000 137.320 ;
    END
  END gfpga_pad_io_soc_dir[67]
  PIN gfpga_pad_io_soc_dir[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.230 0.000 2396.510 4.000 ;
    END
  END gfpga_pad_io_soc_dir[68]
  PIN gfpga_pad_io_soc_dir[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2309.290 0.000 2309.570 4.000 ;
    END
  END gfpga_pad_io_soc_dir[69]
  PIN gfpga_pad_io_soc_dir[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 2711.000 493.490 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[6]
  PIN gfpga_pad_io_soc_dir[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2222.350 0.000 2222.630 4.000 ;
    END
  END gfpga_pad_io_soc_dir[70]
  PIN gfpga_pad_io_soc_dir[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.410 0.000 2135.690 4.000 ;
    END
  END gfpga_pad_io_soc_dir[71]
  PIN gfpga_pad_io_soc_dir[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.470 0.000 2048.750 4.000 ;
    END
  END gfpga_pad_io_soc_dir[72]
  PIN gfpga_pad_io_soc_dir[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.530 0.000 1961.810 4.000 ;
    END
  END gfpga_pad_io_soc_dir[73]
  PIN gfpga_pad_io_soc_dir[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.590 0.000 1874.870 4.000 ;
    END
  END gfpga_pad_io_soc_dir[74]
  PIN gfpga_pad_io_soc_dir[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.650 0.000 1787.930 4.000 ;
    END
  END gfpga_pad_io_soc_dir[75]
  PIN gfpga_pad_io_soc_dir[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.710 0.000 1700.990 4.000 ;
    END
  END gfpga_pad_io_soc_dir[76]
  PIN gfpga_pad_io_soc_dir[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.770 0.000 1614.050 4.000 ;
    END
  END gfpga_pad_io_soc_dir[77]
  PIN gfpga_pad_io_soc_dir[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.830 0.000 1527.110 4.000 ;
    END
  END gfpga_pad_io_soc_dir[78]
  PIN gfpga_pad_io_soc_dir[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 4.000 ;
    END
  END gfpga_pad_io_soc_dir[79]
  PIN gfpga_pad_io_soc_dir[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 2711.000 561.110 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[7]
  PIN gfpga_pad_io_soc_dir[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END gfpga_pad_io_soc_dir[80]
  PIN gfpga_pad_io_soc_dir[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END gfpga_pad_io_soc_dir[81]
  PIN gfpga_pad_io_soc_dir[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.070 0.000 1179.350 4.000 ;
    END
  END gfpga_pad_io_soc_dir[82]
  PIN gfpga_pad_io_soc_dir[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END gfpga_pad_io_soc_dir[83]
  PIN gfpga_pad_io_soc_dir[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END gfpga_pad_io_soc_dir[84]
  PIN gfpga_pad_io_soc_dir[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 0.000 918.530 4.000 ;
    END
  END gfpga_pad_io_soc_dir[85]
  PIN gfpga_pad_io_soc_dir[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END gfpga_pad_io_soc_dir[86]
  PIN gfpga_pad_io_soc_dir[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END gfpga_pad_io_soc_dir[87]
  PIN gfpga_pad_io_soc_dir[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END gfpga_pad_io_soc_dir[88]
  PIN gfpga_pad_io_soc_dir[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END gfpga_pad_io_soc_dir[89]
  PIN gfpga_pad_io_soc_dir[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 2711.000 628.730 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[8]
  PIN gfpga_pad_io_soc_dir[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END gfpga_pad_io_soc_dir[90]
  PIN gfpga_pad_io_soc_dir[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END gfpga_pad_io_soc_dir[91]
  PIN gfpga_pad_io_soc_dir[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END gfpga_pad_io_soc_dir[92]
  PIN gfpga_pad_io_soc_dir[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END gfpga_pad_io_soc_dir[93]
  PIN gfpga_pad_io_soc_dir[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END gfpga_pad_io_soc_dir[94]
  PIN gfpga_pad_io_soc_dir[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END gfpga_pad_io_soc_dir[95]
  PIN gfpga_pad_io_soc_dir[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END gfpga_pad_io_soc_dir[96]
  PIN gfpga_pad_io_soc_dir[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END gfpga_pad_io_soc_dir[97]
  PIN gfpga_pad_io_soc_dir[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END gfpga_pad_io_soc_dir[98]
  PIN gfpga_pad_io_soc_dir[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END gfpga_pad_io_soc_dir[99]
  PIN gfpga_pad_io_soc_dir[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 2711.000 696.350 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[9]
  PIN gfpga_pad_io_soc_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 2711.000 20.150 2715.000 ;
    END
  END gfpga_pad_io_soc_in[0]
  PIN gfpga_pad_io_soc_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END gfpga_pad_io_soc_in[100]
  PIN gfpga_pad_io_soc_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END gfpga_pad_io_soc_in[101]
  PIN gfpga_pad_io_soc_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END gfpga_pad_io_soc_in[102]
  PIN gfpga_pad_io_soc_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END gfpga_pad_io_soc_in[103]
  PIN gfpga_pad_io_soc_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END gfpga_pad_io_soc_in[104]
  PIN gfpga_pad_io_soc_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END gfpga_pad_io_soc_in[105]
  PIN gfpga_pad_io_soc_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END gfpga_pad_io_soc_in[106]
  PIN gfpga_pad_io_soc_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END gfpga_pad_io_soc_in[107]
  PIN gfpga_pad_io_soc_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END gfpga_pad_io_soc_in[108]
  PIN gfpga_pad_io_soc_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END gfpga_pad_io_soc_in[109]
  PIN gfpga_pad_io_soc_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 2711.000 718.890 2715.000 ;
    END
  END gfpga_pad_io_soc_in[10]
  PIN gfpga_pad_io_soc_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END gfpga_pad_io_soc_in[110]
  PIN gfpga_pad_io_soc_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END gfpga_pad_io_soc_in[111]
  PIN gfpga_pad_io_soc_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END gfpga_pad_io_soc_in[112]
  PIN gfpga_pad_io_soc_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END gfpga_pad_io_soc_in[113]
  PIN gfpga_pad_io_soc_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.240 4.000 1574.840 ;
    END
  END gfpga_pad_io_soc_in[114]
  PIN gfpga_pad_io_soc_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1655.840 4.000 1656.440 ;
    END
  END gfpga_pad_io_soc_in[115]
  PIN gfpga_pad_io_soc_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1737.440 4.000 1738.040 ;
    END
  END gfpga_pad_io_soc_in[116]
  PIN gfpga_pad_io_soc_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1819.040 4.000 1819.640 ;
    END
  END gfpga_pad_io_soc_in[117]
  PIN gfpga_pad_io_soc_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1900.640 4.000 1901.240 ;
    END
  END gfpga_pad_io_soc_in[118]
  PIN gfpga_pad_io_soc_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1982.240 4.000 1982.840 ;
    END
  END gfpga_pad_io_soc_in[119]
  PIN gfpga_pad_io_soc_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 2711.000 786.510 2715.000 ;
    END
  END gfpga_pad_io_soc_in[11]
  PIN gfpga_pad_io_soc_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2063.840 4.000 2064.440 ;
    END
  END gfpga_pad_io_soc_in[120]
  PIN gfpga_pad_io_soc_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2145.440 4.000 2146.040 ;
    END
  END gfpga_pad_io_soc_in[121]
  PIN gfpga_pad_io_soc_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2227.040 4.000 2227.640 ;
    END
  END gfpga_pad_io_soc_in[122]
  PIN gfpga_pad_io_soc_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2308.640 4.000 2309.240 ;
    END
  END gfpga_pad_io_soc_in[123]
  PIN gfpga_pad_io_soc_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2390.240 4.000 2390.840 ;
    END
  END gfpga_pad_io_soc_in[124]
  PIN gfpga_pad_io_soc_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2471.840 4.000 2472.440 ;
    END
  END gfpga_pad_io_soc_in[125]
  PIN gfpga_pad_io_soc_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2553.440 4.000 2554.040 ;
    END
  END gfpga_pad_io_soc_in[126]
  PIN gfpga_pad_io_soc_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2635.040 4.000 2635.640 ;
    END
  END gfpga_pad_io_soc_in[127]
  PIN gfpga_pad_io_soc_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 2711.000 854.130 2715.000 ;
    END
  END gfpga_pad_io_soc_in[12]
  PIN gfpga_pad_io_soc_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 2711.000 921.750 2715.000 ;
    END
  END gfpga_pad_io_soc_in[13]
  PIN gfpga_pad_io_soc_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 2711.000 989.370 2715.000 ;
    END
  END gfpga_pad_io_soc_in[14]
  PIN gfpga_pad_io_soc_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 2711.000 1056.990 2715.000 ;
    END
  END gfpga_pad_io_soc_in[15]
  PIN gfpga_pad_io_soc_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 2711.000 1124.610 2715.000 ;
    END
  END gfpga_pad_io_soc_in[16]
  PIN gfpga_pad_io_soc_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 2711.000 1192.230 2715.000 ;
    END
  END gfpga_pad_io_soc_in[17]
  PIN gfpga_pad_io_soc_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.570 2711.000 1259.850 2715.000 ;
    END
  END gfpga_pad_io_soc_in[18]
  PIN gfpga_pad_io_soc_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 2711.000 1327.470 2715.000 ;
    END
  END gfpga_pad_io_soc_in[19]
  PIN gfpga_pad_io_soc_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 2711.000 87.770 2715.000 ;
    END
  END gfpga_pad_io_soc_in[1]
  PIN gfpga_pad_io_soc_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 2711.000 1395.090 2715.000 ;
    END
  END gfpga_pad_io_soc_in[20]
  PIN gfpga_pad_io_soc_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 2711.000 1462.710 2715.000 ;
    END
  END gfpga_pad_io_soc_in[21]
  PIN gfpga_pad_io_soc_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.050 2711.000 1530.330 2715.000 ;
    END
  END gfpga_pad_io_soc_in[22]
  PIN gfpga_pad_io_soc_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 2711.000 1597.950 2715.000 ;
    END
  END gfpga_pad_io_soc_in[23]
  PIN gfpga_pad_io_soc_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.290 2711.000 1665.570 2715.000 ;
    END
  END gfpga_pad_io_soc_in[24]
  PIN gfpga_pad_io_soc_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 2711.000 1733.190 2715.000 ;
    END
  END gfpga_pad_io_soc_in[25]
  PIN gfpga_pad_io_soc_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.530 2711.000 1800.810 2715.000 ;
    END
  END gfpga_pad_io_soc_in[26]
  PIN gfpga_pad_io_soc_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 2711.000 1868.430 2715.000 ;
    END
  END gfpga_pad_io_soc_in[27]
  PIN gfpga_pad_io_soc_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.770 2711.000 1936.050 2715.000 ;
    END
  END gfpga_pad_io_soc_in[28]
  PIN gfpga_pad_io_soc_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.390 2711.000 2003.670 2715.000 ;
    END
  END gfpga_pad_io_soc_in[29]
  PIN gfpga_pad_io_soc_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 2711.000 155.390 2715.000 ;
    END
  END gfpga_pad_io_soc_in[2]
  PIN gfpga_pad_io_soc_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.010 2711.000 2071.290 2715.000 ;
    END
  END gfpga_pad_io_soc_in[30]
  PIN gfpga_pad_io_soc_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.630 2711.000 2138.910 2715.000 ;
    END
  END gfpga_pad_io_soc_in[31]
  PIN gfpga_pad_io_soc_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.250 2711.000 2206.530 2715.000 ;
    END
  END gfpga_pad_io_soc_in[32]
  PIN gfpga_pad_io_soc_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.870 2711.000 2274.150 2715.000 ;
    END
  END gfpga_pad_io_soc_in[33]
  PIN gfpga_pad_io_soc_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.490 2711.000 2341.770 2715.000 ;
    END
  END gfpga_pad_io_soc_in[34]
  PIN gfpga_pad_io_soc_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2409.110 2711.000 2409.390 2715.000 ;
    END
  END gfpga_pad_io_soc_in[35]
  PIN gfpga_pad_io_soc_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2656.120 2475.000 2656.720 ;
    END
  END gfpga_pad_io_soc_in[36]
  PIN gfpga_pad_io_soc_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2576.560 2475.000 2577.160 ;
    END
  END gfpga_pad_io_soc_in[37]
  PIN gfpga_pad_io_soc_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2497.000 2475.000 2497.600 ;
    END
  END gfpga_pad_io_soc_in[38]
  PIN gfpga_pad_io_soc_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2417.440 2475.000 2418.040 ;
    END
  END gfpga_pad_io_soc_in[39]
  PIN gfpga_pad_io_soc_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 2711.000 223.010 2715.000 ;
    END
  END gfpga_pad_io_soc_in[3]
  PIN gfpga_pad_io_soc_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2337.880 2475.000 2338.480 ;
    END
  END gfpga_pad_io_soc_in[40]
  PIN gfpga_pad_io_soc_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2258.320 2475.000 2258.920 ;
    END
  END gfpga_pad_io_soc_in[41]
  PIN gfpga_pad_io_soc_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2178.760 2475.000 2179.360 ;
    END
  END gfpga_pad_io_soc_in[42]
  PIN gfpga_pad_io_soc_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2099.200 2475.000 2099.800 ;
    END
  END gfpga_pad_io_soc_in[43]
  PIN gfpga_pad_io_soc_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2019.640 2475.000 2020.240 ;
    END
  END gfpga_pad_io_soc_in[44]
  PIN gfpga_pad_io_soc_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1940.080 2475.000 1940.680 ;
    END
  END gfpga_pad_io_soc_in[45]
  PIN gfpga_pad_io_soc_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1860.520 2475.000 1861.120 ;
    END
  END gfpga_pad_io_soc_in[46]
  PIN gfpga_pad_io_soc_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1780.960 2475.000 1781.560 ;
    END
  END gfpga_pad_io_soc_in[47]
  PIN gfpga_pad_io_soc_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1701.400 2475.000 1702.000 ;
    END
  END gfpga_pad_io_soc_in[48]
  PIN gfpga_pad_io_soc_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1621.840 2475.000 1622.440 ;
    END
  END gfpga_pad_io_soc_in[49]
  PIN gfpga_pad_io_soc_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 2711.000 313.170 2715.000 ;
    END
  END gfpga_pad_io_soc_in[4]
  PIN gfpga_pad_io_soc_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1542.280 2475.000 1542.880 ;
    END
  END gfpga_pad_io_soc_in[50]
  PIN gfpga_pad_io_soc_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1462.720 2475.000 1463.320 ;
    END
  END gfpga_pad_io_soc_in[51]
  PIN gfpga_pad_io_soc_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1383.160 2475.000 1383.760 ;
    END
  END gfpga_pad_io_soc_in[52]
  PIN gfpga_pad_io_soc_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1303.600 2475.000 1304.200 ;
    END
  END gfpga_pad_io_soc_in[53]
  PIN gfpga_pad_io_soc_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1224.040 2475.000 1224.640 ;
    END
  END gfpga_pad_io_soc_in[54]
  PIN gfpga_pad_io_soc_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1144.480 2475.000 1145.080 ;
    END
  END gfpga_pad_io_soc_in[55]
  PIN gfpga_pad_io_soc_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1064.920 2475.000 1065.520 ;
    END
  END gfpga_pad_io_soc_in[56]
  PIN gfpga_pad_io_soc_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 985.360 2475.000 985.960 ;
    END
  END gfpga_pad_io_soc_in[57]
  PIN gfpga_pad_io_soc_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 905.800 2475.000 906.400 ;
    END
  END gfpga_pad_io_soc_in[58]
  PIN gfpga_pad_io_soc_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 826.240 2475.000 826.840 ;
    END
  END gfpga_pad_io_soc_in[59]
  PIN gfpga_pad_io_soc_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 2711.000 380.790 2715.000 ;
    END
  END gfpga_pad_io_soc_in[5]
  PIN gfpga_pad_io_soc_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 746.680 2475.000 747.280 ;
    END
  END gfpga_pad_io_soc_in[60]
  PIN gfpga_pad_io_soc_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 667.120 2475.000 667.720 ;
    END
  END gfpga_pad_io_soc_in[61]
  PIN gfpga_pad_io_soc_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 587.560 2475.000 588.160 ;
    END
  END gfpga_pad_io_soc_in[62]
  PIN gfpga_pad_io_soc_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 508.000 2475.000 508.600 ;
    END
  END gfpga_pad_io_soc_in[63]
  PIN gfpga_pad_io_soc_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 428.440 2475.000 429.040 ;
    END
  END gfpga_pad_io_soc_in[64]
  PIN gfpga_pad_io_soc_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 348.880 2475.000 349.480 ;
    END
  END gfpga_pad_io_soc_in[65]
  PIN gfpga_pad_io_soc_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 269.320 2475.000 269.920 ;
    END
  END gfpga_pad_io_soc_in[66]
  PIN gfpga_pad_io_soc_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 189.760 2475.000 190.360 ;
    END
  END gfpga_pad_io_soc_in[67]
  PIN gfpga_pad_io_soc_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.190 0.000 2454.470 4.000 ;
    END
  END gfpga_pad_io_soc_in[68]
  PIN gfpga_pad_io_soc_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.250 0.000 2367.530 4.000 ;
    END
  END gfpga_pad_io_soc_in[69]
  PIN gfpga_pad_io_soc_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 2711.000 448.410 2715.000 ;
    END
  END gfpga_pad_io_soc_in[6]
  PIN gfpga_pad_io_soc_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.310 0.000 2280.590 4.000 ;
    END
  END gfpga_pad_io_soc_in[70]
  PIN gfpga_pad_io_soc_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.370 0.000 2193.650 4.000 ;
    END
  END gfpga_pad_io_soc_in[71]
  PIN gfpga_pad_io_soc_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.430 0.000 2106.710 4.000 ;
    END
  END gfpga_pad_io_soc_in[72]
  PIN gfpga_pad_io_soc_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.490 0.000 2019.770 4.000 ;
    END
  END gfpga_pad_io_soc_in[73]
  PIN gfpga_pad_io_soc_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.550 0.000 1932.830 4.000 ;
    END
  END gfpga_pad_io_soc_in[74]
  PIN gfpga_pad_io_soc_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.610 0.000 1845.890 4.000 ;
    END
  END gfpga_pad_io_soc_in[75]
  PIN gfpga_pad_io_soc_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.670 0.000 1758.950 4.000 ;
    END
  END gfpga_pad_io_soc_in[76]
  PIN gfpga_pad_io_soc_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.730 0.000 1672.010 4.000 ;
    END
  END gfpga_pad_io_soc_in[77]
  PIN gfpga_pad_io_soc_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 0.000 1585.070 4.000 ;
    END
  END gfpga_pad_io_soc_in[78]
  PIN gfpga_pad_io_soc_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.850 0.000 1498.130 4.000 ;
    END
  END gfpga_pad_io_soc_in[79]
  PIN gfpga_pad_io_soc_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 2711.000 516.030 2715.000 ;
    END
  END gfpga_pad_io_soc_in[7]
  PIN gfpga_pad_io_soc_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 0.000 1411.190 4.000 ;
    END
  END gfpga_pad_io_soc_in[80]
  PIN gfpga_pad_io_soc_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 4.000 ;
    END
  END gfpga_pad_io_soc_in[81]
  PIN gfpga_pad_io_soc_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 0.000 1237.310 4.000 ;
    END
  END gfpga_pad_io_soc_in[82]
  PIN gfpga_pad_io_soc_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END gfpga_pad_io_soc_in[83]
  PIN gfpga_pad_io_soc_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 0.000 1063.430 4.000 ;
    END
  END gfpga_pad_io_soc_in[84]
  PIN gfpga_pad_io_soc_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END gfpga_pad_io_soc_in[85]
  PIN gfpga_pad_io_soc_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 0.000 889.550 4.000 ;
    END
  END gfpga_pad_io_soc_in[86]
  PIN gfpga_pad_io_soc_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END gfpga_pad_io_soc_in[87]
  PIN gfpga_pad_io_soc_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END gfpga_pad_io_soc_in[88]
  PIN gfpga_pad_io_soc_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END gfpga_pad_io_soc_in[89]
  PIN gfpga_pad_io_soc_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 2711.000 583.650 2715.000 ;
    END
  END gfpga_pad_io_soc_in[8]
  PIN gfpga_pad_io_soc_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END gfpga_pad_io_soc_in[90]
  PIN gfpga_pad_io_soc_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END gfpga_pad_io_soc_in[91]
  PIN gfpga_pad_io_soc_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END gfpga_pad_io_soc_in[92]
  PIN gfpga_pad_io_soc_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END gfpga_pad_io_soc_in[93]
  PIN gfpga_pad_io_soc_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END gfpga_pad_io_soc_in[94]
  PIN gfpga_pad_io_soc_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END gfpga_pad_io_soc_in[95]
  PIN gfpga_pad_io_soc_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END gfpga_pad_io_soc_in[96]
  PIN gfpga_pad_io_soc_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END gfpga_pad_io_soc_in[97]
  PIN gfpga_pad_io_soc_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END gfpga_pad_io_soc_in[98]
  PIN gfpga_pad_io_soc_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END gfpga_pad_io_soc_in[99]
  PIN gfpga_pad_io_soc_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 2711.000 651.270 2715.000 ;
    END
  END gfpga_pad_io_soc_in[9]
  PIN gfpga_pad_io_soc_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 2711.000 42.690 2715.000 ;
    END
  END gfpga_pad_io_soc_out[0]
  PIN gfpga_pad_io_soc_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END gfpga_pad_io_soc_out[100]
  PIN gfpga_pad_io_soc_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END gfpga_pad_io_soc_out[101]
  PIN gfpga_pad_io_soc_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END gfpga_pad_io_soc_out[102]
  PIN gfpga_pad_io_soc_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END gfpga_pad_io_soc_out[103]
  PIN gfpga_pad_io_soc_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END gfpga_pad_io_soc_out[104]
  PIN gfpga_pad_io_soc_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END gfpga_pad_io_soc_out[105]
  PIN gfpga_pad_io_soc_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END gfpga_pad_io_soc_out[106]
  PIN gfpga_pad_io_soc_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END gfpga_pad_io_soc_out[107]
  PIN gfpga_pad_io_soc_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END gfpga_pad_io_soc_out[108]
  PIN gfpga_pad_io_soc_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END gfpga_pad_io_soc_out[109]
  PIN gfpga_pad_io_soc_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 2711.000 741.430 2715.000 ;
    END
  END gfpga_pad_io_soc_out[10]
  PIN gfpga_pad_io_soc_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END gfpga_pad_io_soc_out[110]
  PIN gfpga_pad_io_soc_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END gfpga_pad_io_soc_out[111]
  PIN gfpga_pad_io_soc_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.240 4.000 1438.840 ;
    END
  END gfpga_pad_io_soc_out[112]
  PIN gfpga_pad_io_soc_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.840 4.000 1520.440 ;
    END
  END gfpga_pad_io_soc_out[113]
  PIN gfpga_pad_io_soc_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1601.440 4.000 1602.040 ;
    END
  END gfpga_pad_io_soc_out[114]
  PIN gfpga_pad_io_soc_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END gfpga_pad_io_soc_out[115]
  PIN gfpga_pad_io_soc_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1764.640 4.000 1765.240 ;
    END
  END gfpga_pad_io_soc_out[116]
  PIN gfpga_pad_io_soc_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1846.240 4.000 1846.840 ;
    END
  END gfpga_pad_io_soc_out[117]
  PIN gfpga_pad_io_soc_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END gfpga_pad_io_soc_out[118]
  PIN gfpga_pad_io_soc_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2009.440 4.000 2010.040 ;
    END
  END gfpga_pad_io_soc_out[119]
  PIN gfpga_pad_io_soc_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 2711.000 809.050 2715.000 ;
    END
  END gfpga_pad_io_soc_out[11]
  PIN gfpga_pad_io_soc_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2091.040 4.000 2091.640 ;
    END
  END gfpga_pad_io_soc_out[120]
  PIN gfpga_pad_io_soc_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2172.640 4.000 2173.240 ;
    END
  END gfpga_pad_io_soc_out[121]
  PIN gfpga_pad_io_soc_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2254.240 4.000 2254.840 ;
    END
  END gfpga_pad_io_soc_out[122]
  PIN gfpga_pad_io_soc_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2335.840 4.000 2336.440 ;
    END
  END gfpga_pad_io_soc_out[123]
  PIN gfpga_pad_io_soc_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2417.440 4.000 2418.040 ;
    END
  END gfpga_pad_io_soc_out[124]
  PIN gfpga_pad_io_soc_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2499.040 4.000 2499.640 ;
    END
  END gfpga_pad_io_soc_out[125]
  PIN gfpga_pad_io_soc_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2580.640 4.000 2581.240 ;
    END
  END gfpga_pad_io_soc_out[126]
  PIN gfpga_pad_io_soc_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2662.240 4.000 2662.840 ;
    END
  END gfpga_pad_io_soc_out[127]
  PIN gfpga_pad_io_soc_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 2711.000 876.670 2715.000 ;
    END
  END gfpga_pad_io_soc_out[12]
  PIN gfpga_pad_io_soc_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 2711.000 944.290 2715.000 ;
    END
  END gfpga_pad_io_soc_out[13]
  PIN gfpga_pad_io_soc_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 2711.000 1011.910 2715.000 ;
    END
  END gfpga_pad_io_soc_out[14]
  PIN gfpga_pad_io_soc_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 2711.000 1079.530 2715.000 ;
    END
  END gfpga_pad_io_soc_out[15]
  PIN gfpga_pad_io_soc_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 2711.000 1147.150 2715.000 ;
    END
  END gfpga_pad_io_soc_out[16]
  PIN gfpga_pad_io_soc_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 2711.000 1214.770 2715.000 ;
    END
  END gfpga_pad_io_soc_out[17]
  PIN gfpga_pad_io_soc_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 2711.000 1282.390 2715.000 ;
    END
  END gfpga_pad_io_soc_out[18]
  PIN gfpga_pad_io_soc_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 2711.000 1350.010 2715.000 ;
    END
  END gfpga_pad_io_soc_out[19]
  PIN gfpga_pad_io_soc_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 2711.000 110.310 2715.000 ;
    END
  END gfpga_pad_io_soc_out[1]
  PIN gfpga_pad_io_soc_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 2711.000 1417.630 2715.000 ;
    END
  END gfpga_pad_io_soc_out[20]
  PIN gfpga_pad_io_soc_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 2711.000 1485.250 2715.000 ;
    END
  END gfpga_pad_io_soc_out[21]
  PIN gfpga_pad_io_soc_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.590 2711.000 1552.870 2715.000 ;
    END
  END gfpga_pad_io_soc_out[22]
  PIN gfpga_pad_io_soc_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.210 2711.000 1620.490 2715.000 ;
    END
  END gfpga_pad_io_soc_out[23]
  PIN gfpga_pad_io_soc_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 2711.000 1688.110 2715.000 ;
    END
  END gfpga_pad_io_soc_out[24]
  PIN gfpga_pad_io_soc_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.450 2711.000 1755.730 2715.000 ;
    END
  END gfpga_pad_io_soc_out[25]
  PIN gfpga_pad_io_soc_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.070 2711.000 1823.350 2715.000 ;
    END
  END gfpga_pad_io_soc_out[26]
  PIN gfpga_pad_io_soc_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.690 2711.000 1890.970 2715.000 ;
    END
  END gfpga_pad_io_soc_out[27]
  PIN gfpga_pad_io_soc_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.310 2711.000 1958.590 2715.000 ;
    END
  END gfpga_pad_io_soc_out[28]
  PIN gfpga_pad_io_soc_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.930 2711.000 2026.210 2715.000 ;
    END
  END gfpga_pad_io_soc_out[29]
  PIN gfpga_pad_io_soc_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 2711.000 177.930 2715.000 ;
    END
  END gfpga_pad_io_soc_out[2]
  PIN gfpga_pad_io_soc_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.550 2711.000 2093.830 2715.000 ;
    END
  END gfpga_pad_io_soc_out[30]
  PIN gfpga_pad_io_soc_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.170 2711.000 2161.450 2715.000 ;
    END
  END gfpga_pad_io_soc_out[31]
  PIN gfpga_pad_io_soc_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.790 2711.000 2229.070 2715.000 ;
    END
  END gfpga_pad_io_soc_out[32]
  PIN gfpga_pad_io_soc_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2296.410 2711.000 2296.690 2715.000 ;
    END
  END gfpga_pad_io_soc_out[33]
  PIN gfpga_pad_io_soc_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.030 2711.000 2364.310 2715.000 ;
    END
  END gfpga_pad_io_soc_out[34]
  PIN gfpga_pad_io_soc_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.650 2711.000 2431.930 2715.000 ;
    END
  END gfpga_pad_io_soc_out[35]
  PIN gfpga_pad_io_soc_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2629.600 2475.000 2630.200 ;
    END
  END gfpga_pad_io_soc_out[36]
  PIN gfpga_pad_io_soc_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2550.040 2475.000 2550.640 ;
    END
  END gfpga_pad_io_soc_out[37]
  PIN gfpga_pad_io_soc_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2470.480 2475.000 2471.080 ;
    END
  END gfpga_pad_io_soc_out[38]
  PIN gfpga_pad_io_soc_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2390.920 2475.000 2391.520 ;
    END
  END gfpga_pad_io_soc_out[39]
  PIN gfpga_pad_io_soc_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 2711.000 245.550 2715.000 ;
    END
  END gfpga_pad_io_soc_out[3]
  PIN gfpga_pad_io_soc_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2311.360 2475.000 2311.960 ;
    END
  END gfpga_pad_io_soc_out[40]
  PIN gfpga_pad_io_soc_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2231.800 2475.000 2232.400 ;
    END
  END gfpga_pad_io_soc_out[41]
  PIN gfpga_pad_io_soc_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2152.240 2475.000 2152.840 ;
    END
  END gfpga_pad_io_soc_out[42]
  PIN gfpga_pad_io_soc_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2072.680 2475.000 2073.280 ;
    END
  END gfpga_pad_io_soc_out[43]
  PIN gfpga_pad_io_soc_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1993.120 2475.000 1993.720 ;
    END
  END gfpga_pad_io_soc_out[44]
  PIN gfpga_pad_io_soc_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1913.560 2475.000 1914.160 ;
    END
  END gfpga_pad_io_soc_out[45]
  PIN gfpga_pad_io_soc_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1834.000 2475.000 1834.600 ;
    END
  END gfpga_pad_io_soc_out[46]
  PIN gfpga_pad_io_soc_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1754.440 2475.000 1755.040 ;
    END
  END gfpga_pad_io_soc_out[47]
  PIN gfpga_pad_io_soc_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1674.880 2475.000 1675.480 ;
    END
  END gfpga_pad_io_soc_out[48]
  PIN gfpga_pad_io_soc_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1595.320 2475.000 1595.920 ;
    END
  END gfpga_pad_io_soc_out[49]
  PIN gfpga_pad_io_soc_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 2711.000 335.710 2715.000 ;
    END
  END gfpga_pad_io_soc_out[4]
  PIN gfpga_pad_io_soc_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1515.760 2475.000 1516.360 ;
    END
  END gfpga_pad_io_soc_out[50]
  PIN gfpga_pad_io_soc_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1436.200 2475.000 1436.800 ;
    END
  END gfpga_pad_io_soc_out[51]
  PIN gfpga_pad_io_soc_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1356.640 2475.000 1357.240 ;
    END
  END gfpga_pad_io_soc_out[52]
  PIN gfpga_pad_io_soc_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1277.080 2475.000 1277.680 ;
    END
  END gfpga_pad_io_soc_out[53]
  PIN gfpga_pad_io_soc_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1197.520 2475.000 1198.120 ;
    END
  END gfpga_pad_io_soc_out[54]
  PIN gfpga_pad_io_soc_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1117.960 2475.000 1118.560 ;
    END
  END gfpga_pad_io_soc_out[55]
  PIN gfpga_pad_io_soc_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1038.400 2475.000 1039.000 ;
    END
  END gfpga_pad_io_soc_out[56]
  PIN gfpga_pad_io_soc_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 958.840 2475.000 959.440 ;
    END
  END gfpga_pad_io_soc_out[57]
  PIN gfpga_pad_io_soc_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 879.280 2475.000 879.880 ;
    END
  END gfpga_pad_io_soc_out[58]
  PIN gfpga_pad_io_soc_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 799.720 2475.000 800.320 ;
    END
  END gfpga_pad_io_soc_out[59]
  PIN gfpga_pad_io_soc_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 2711.000 403.330 2715.000 ;
    END
  END gfpga_pad_io_soc_out[5]
  PIN gfpga_pad_io_soc_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 720.160 2475.000 720.760 ;
    END
  END gfpga_pad_io_soc_out[60]
  PIN gfpga_pad_io_soc_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 640.600 2475.000 641.200 ;
    END
  END gfpga_pad_io_soc_out[61]
  PIN gfpga_pad_io_soc_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 561.040 2475.000 561.640 ;
    END
  END gfpga_pad_io_soc_out[62]
  PIN gfpga_pad_io_soc_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 481.480 2475.000 482.080 ;
    END
  END gfpga_pad_io_soc_out[63]
  PIN gfpga_pad_io_soc_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 401.920 2475.000 402.520 ;
    END
  END gfpga_pad_io_soc_out[64]
  PIN gfpga_pad_io_soc_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 322.360 2475.000 322.960 ;
    END
  END gfpga_pad_io_soc_out[65]
  PIN gfpga_pad_io_soc_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 242.800 2475.000 243.400 ;
    END
  END gfpga_pad_io_soc_out[66]
  PIN gfpga_pad_io_soc_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 163.240 2475.000 163.840 ;
    END
  END gfpga_pad_io_soc_out[67]
  PIN gfpga_pad_io_soc_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.210 0.000 2425.490 4.000 ;
    END
  END gfpga_pad_io_soc_out[68]
  PIN gfpga_pad_io_soc_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.270 0.000 2338.550 4.000 ;
    END
  END gfpga_pad_io_soc_out[69]
  PIN gfpga_pad_io_soc_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 2711.000 470.950 2715.000 ;
    END
  END gfpga_pad_io_soc_out[6]
  PIN gfpga_pad_io_soc_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.330 0.000 2251.610 4.000 ;
    END
  END gfpga_pad_io_soc_out[70]
  PIN gfpga_pad_io_soc_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.390 0.000 2164.670 4.000 ;
    END
  END gfpga_pad_io_soc_out[71]
  PIN gfpga_pad_io_soc_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.450 0.000 2077.730 4.000 ;
    END
  END gfpga_pad_io_soc_out[72]
  PIN gfpga_pad_io_soc_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.510 0.000 1990.790 4.000 ;
    END
  END gfpga_pad_io_soc_out[73]
  PIN gfpga_pad_io_soc_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END gfpga_pad_io_soc_out[74]
  PIN gfpga_pad_io_soc_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.630 0.000 1816.910 4.000 ;
    END
  END gfpga_pad_io_soc_out[75]
  PIN gfpga_pad_io_soc_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.690 0.000 1729.970 4.000 ;
    END
  END gfpga_pad_io_soc_out[76]
  PIN gfpga_pad_io_soc_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.750 0.000 1643.030 4.000 ;
    END
  END gfpga_pad_io_soc_out[77]
  PIN gfpga_pad_io_soc_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.810 0.000 1556.090 4.000 ;
    END
  END gfpga_pad_io_soc_out[78]
  PIN gfpga_pad_io_soc_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.870 0.000 1469.150 4.000 ;
    END
  END gfpga_pad_io_soc_out[79]
  PIN gfpga_pad_io_soc_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 2711.000 538.570 2715.000 ;
    END
  END gfpga_pad_io_soc_out[7]
  PIN gfpga_pad_io_soc_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 0.000 1382.210 4.000 ;
    END
  END gfpga_pad_io_soc_out[80]
  PIN gfpga_pad_io_soc_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 0.000 1295.270 4.000 ;
    END
  END gfpga_pad_io_soc_out[81]
  PIN gfpga_pad_io_soc_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.050 0.000 1208.330 4.000 ;
    END
  END gfpga_pad_io_soc_out[82]
  PIN gfpga_pad_io_soc_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END gfpga_pad_io_soc_out[83]
  PIN gfpga_pad_io_soc_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 4.000 ;
    END
  END gfpga_pad_io_soc_out[84]
  PIN gfpga_pad_io_soc_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END gfpga_pad_io_soc_out[85]
  PIN gfpga_pad_io_soc_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END gfpga_pad_io_soc_out[86]
  PIN gfpga_pad_io_soc_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END gfpga_pad_io_soc_out[87]
  PIN gfpga_pad_io_soc_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END gfpga_pad_io_soc_out[88]
  PIN gfpga_pad_io_soc_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END gfpga_pad_io_soc_out[89]
  PIN gfpga_pad_io_soc_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 2711.000 606.190 2715.000 ;
    END
  END gfpga_pad_io_soc_out[8]
  PIN gfpga_pad_io_soc_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END gfpga_pad_io_soc_out[90]
  PIN gfpga_pad_io_soc_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END gfpga_pad_io_soc_out[91]
  PIN gfpga_pad_io_soc_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END gfpga_pad_io_soc_out[92]
  PIN gfpga_pad_io_soc_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END gfpga_pad_io_soc_out[93]
  PIN gfpga_pad_io_soc_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END gfpga_pad_io_soc_out[94]
  PIN gfpga_pad_io_soc_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END gfpga_pad_io_soc_out[95]
  PIN gfpga_pad_io_soc_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END gfpga_pad_io_soc_out[96]
  PIN gfpga_pad_io_soc_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END gfpga_pad_io_soc_out[97]
  PIN gfpga_pad_io_soc_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END gfpga_pad_io_soc_out[98]
  PIN gfpga_pad_io_soc_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END gfpga_pad_io_soc_out[99]
  PIN gfpga_pad_io_soc_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 2711.000 673.810 2715.000 ;
    END
  END gfpga_pad_io_soc_out[9]
  PIN isol_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 57.160 2475.000 57.760 ;
    END
  END isol_n
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END prog_clk
  PIN prog_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 83.680 2475.000 84.280 ;
    END
  END prog_reset
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 110.200 2475.000 110.800 ;
    END
  END reset
  PIN sc_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 2711.000 290.630 2715.000 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2682.640 2475.000 2683.240 ;
    END
  END sc_tail
  PIN test_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 30.640 2475.000 31.240 ;
    END
  END test_enable
  OBS
      LAYER li1 ;
        RECT 1.840 10.795 2472.960 2703.765 ;
      LAYER met1 ;
        RECT 1.840 9.900 2472.960 2703.920 ;
      LAYER met2 ;
        RECT 3.770 2710.720 19.590 2711.570 ;
        RECT 20.430 2710.720 42.130 2711.570 ;
        RECT 42.970 2710.720 64.670 2711.570 ;
        RECT 65.510 2710.720 87.210 2711.570 ;
        RECT 88.050 2710.720 109.750 2711.570 ;
        RECT 110.590 2710.720 132.290 2711.570 ;
        RECT 133.130 2710.720 154.830 2711.570 ;
        RECT 155.670 2710.720 177.370 2711.570 ;
        RECT 178.210 2710.720 199.910 2711.570 ;
        RECT 200.750 2710.720 222.450 2711.570 ;
        RECT 223.290 2710.720 244.990 2711.570 ;
        RECT 245.830 2710.720 267.530 2711.570 ;
        RECT 268.370 2710.720 290.070 2711.570 ;
        RECT 290.910 2710.720 312.610 2711.570 ;
        RECT 313.450 2710.720 335.150 2711.570 ;
        RECT 335.990 2710.720 357.690 2711.570 ;
        RECT 358.530 2710.720 380.230 2711.570 ;
        RECT 381.070 2710.720 402.770 2711.570 ;
        RECT 403.610 2710.720 425.310 2711.570 ;
        RECT 426.150 2710.720 447.850 2711.570 ;
        RECT 448.690 2710.720 470.390 2711.570 ;
        RECT 471.230 2710.720 492.930 2711.570 ;
        RECT 493.770 2710.720 515.470 2711.570 ;
        RECT 516.310 2710.720 538.010 2711.570 ;
        RECT 538.850 2710.720 560.550 2711.570 ;
        RECT 561.390 2710.720 583.090 2711.570 ;
        RECT 583.930 2710.720 605.630 2711.570 ;
        RECT 606.470 2710.720 628.170 2711.570 ;
        RECT 629.010 2710.720 650.710 2711.570 ;
        RECT 651.550 2710.720 673.250 2711.570 ;
        RECT 674.090 2710.720 695.790 2711.570 ;
        RECT 696.630 2710.720 718.330 2711.570 ;
        RECT 719.170 2710.720 740.870 2711.570 ;
        RECT 741.710 2710.720 763.410 2711.570 ;
        RECT 764.250 2710.720 785.950 2711.570 ;
        RECT 786.790 2710.720 808.490 2711.570 ;
        RECT 809.330 2710.720 831.030 2711.570 ;
        RECT 831.870 2710.720 853.570 2711.570 ;
        RECT 854.410 2710.720 876.110 2711.570 ;
        RECT 876.950 2710.720 898.650 2711.570 ;
        RECT 899.490 2710.720 921.190 2711.570 ;
        RECT 922.030 2710.720 943.730 2711.570 ;
        RECT 944.570 2710.720 966.270 2711.570 ;
        RECT 967.110 2710.720 988.810 2711.570 ;
        RECT 989.650 2710.720 1011.350 2711.570 ;
        RECT 1012.190 2710.720 1033.890 2711.570 ;
        RECT 1034.730 2710.720 1056.430 2711.570 ;
        RECT 1057.270 2710.720 1078.970 2711.570 ;
        RECT 1079.810 2710.720 1101.510 2711.570 ;
        RECT 1102.350 2710.720 1124.050 2711.570 ;
        RECT 1124.890 2710.720 1146.590 2711.570 ;
        RECT 1147.430 2710.720 1169.130 2711.570 ;
        RECT 1169.970 2710.720 1191.670 2711.570 ;
        RECT 1192.510 2710.720 1214.210 2711.570 ;
        RECT 1215.050 2710.720 1236.750 2711.570 ;
        RECT 1237.590 2710.720 1259.290 2711.570 ;
        RECT 1260.130 2710.720 1281.830 2711.570 ;
        RECT 1282.670 2710.720 1304.370 2711.570 ;
        RECT 1305.210 2710.720 1326.910 2711.570 ;
        RECT 1327.750 2710.720 1349.450 2711.570 ;
        RECT 1350.290 2710.720 1371.990 2711.570 ;
        RECT 1372.830 2710.720 1394.530 2711.570 ;
        RECT 1395.370 2710.720 1417.070 2711.570 ;
        RECT 1417.910 2710.720 1439.610 2711.570 ;
        RECT 1440.450 2710.720 1462.150 2711.570 ;
        RECT 1462.990 2710.720 1484.690 2711.570 ;
        RECT 1485.530 2710.720 1507.230 2711.570 ;
        RECT 1508.070 2710.720 1529.770 2711.570 ;
        RECT 1530.610 2710.720 1552.310 2711.570 ;
        RECT 1553.150 2710.720 1574.850 2711.570 ;
        RECT 1575.690 2710.720 1597.390 2711.570 ;
        RECT 1598.230 2710.720 1619.930 2711.570 ;
        RECT 1620.770 2710.720 1642.470 2711.570 ;
        RECT 1643.310 2710.720 1665.010 2711.570 ;
        RECT 1665.850 2710.720 1687.550 2711.570 ;
        RECT 1688.390 2710.720 1710.090 2711.570 ;
        RECT 1710.930 2710.720 1732.630 2711.570 ;
        RECT 1733.470 2710.720 1755.170 2711.570 ;
        RECT 1756.010 2710.720 1777.710 2711.570 ;
        RECT 1778.550 2710.720 1800.250 2711.570 ;
        RECT 1801.090 2710.720 1822.790 2711.570 ;
        RECT 1823.630 2710.720 1845.330 2711.570 ;
        RECT 1846.170 2710.720 1867.870 2711.570 ;
        RECT 1868.710 2710.720 1890.410 2711.570 ;
        RECT 1891.250 2710.720 1912.950 2711.570 ;
        RECT 1913.790 2710.720 1935.490 2711.570 ;
        RECT 1936.330 2710.720 1958.030 2711.570 ;
        RECT 1958.870 2710.720 1980.570 2711.570 ;
        RECT 1981.410 2710.720 2003.110 2711.570 ;
        RECT 2003.950 2710.720 2025.650 2711.570 ;
        RECT 2026.490 2710.720 2048.190 2711.570 ;
        RECT 2049.030 2710.720 2070.730 2711.570 ;
        RECT 2071.570 2710.720 2093.270 2711.570 ;
        RECT 2094.110 2710.720 2115.810 2711.570 ;
        RECT 2116.650 2710.720 2138.350 2711.570 ;
        RECT 2139.190 2710.720 2160.890 2711.570 ;
        RECT 2161.730 2710.720 2183.430 2711.570 ;
        RECT 2184.270 2710.720 2205.970 2711.570 ;
        RECT 2206.810 2710.720 2228.510 2711.570 ;
        RECT 2229.350 2710.720 2251.050 2711.570 ;
        RECT 2251.890 2710.720 2273.590 2711.570 ;
        RECT 2274.430 2710.720 2296.130 2711.570 ;
        RECT 2296.970 2710.720 2318.670 2711.570 ;
        RECT 2319.510 2710.720 2341.210 2711.570 ;
        RECT 2342.050 2710.720 2363.750 2711.570 ;
        RECT 2364.590 2710.720 2386.290 2711.570 ;
        RECT 2387.130 2710.720 2408.830 2711.570 ;
        RECT 2409.670 2710.720 2431.370 2711.570 ;
        RECT 2432.210 2710.720 2453.910 2711.570 ;
        RECT 2454.750 2710.720 2471.020 2711.570 ;
        RECT 3.770 4.280 2471.020 2710.720 ;
        RECT 3.770 3.670 19.590 4.280 ;
        RECT 20.430 3.670 48.570 4.280 ;
        RECT 49.410 3.670 77.550 4.280 ;
        RECT 78.390 3.670 106.530 4.280 ;
        RECT 107.370 3.670 135.510 4.280 ;
        RECT 136.350 3.670 164.490 4.280 ;
        RECT 165.330 3.670 193.470 4.280 ;
        RECT 194.310 3.670 222.450 4.280 ;
        RECT 223.290 3.670 251.430 4.280 ;
        RECT 252.270 3.670 280.410 4.280 ;
        RECT 281.250 3.670 309.390 4.280 ;
        RECT 310.230 3.670 338.370 4.280 ;
        RECT 339.210 3.670 367.350 4.280 ;
        RECT 368.190 3.670 396.330 4.280 ;
        RECT 397.170 3.670 425.310 4.280 ;
        RECT 426.150 3.670 454.290 4.280 ;
        RECT 455.130 3.670 483.270 4.280 ;
        RECT 484.110 3.670 512.250 4.280 ;
        RECT 513.090 3.670 541.230 4.280 ;
        RECT 542.070 3.670 570.210 4.280 ;
        RECT 571.050 3.670 599.190 4.280 ;
        RECT 600.030 3.670 628.170 4.280 ;
        RECT 629.010 3.670 657.150 4.280 ;
        RECT 657.990 3.670 686.130 4.280 ;
        RECT 686.970 3.670 715.110 4.280 ;
        RECT 715.950 3.670 744.090 4.280 ;
        RECT 744.930 3.670 773.070 4.280 ;
        RECT 773.910 3.670 802.050 4.280 ;
        RECT 802.890 3.670 831.030 4.280 ;
        RECT 831.870 3.670 860.010 4.280 ;
        RECT 860.850 3.670 888.990 4.280 ;
        RECT 889.830 3.670 917.970 4.280 ;
        RECT 918.810 3.670 946.950 4.280 ;
        RECT 947.790 3.670 975.930 4.280 ;
        RECT 976.770 3.670 1004.910 4.280 ;
        RECT 1005.750 3.670 1033.890 4.280 ;
        RECT 1034.730 3.670 1062.870 4.280 ;
        RECT 1063.710 3.670 1091.850 4.280 ;
        RECT 1092.690 3.670 1120.830 4.280 ;
        RECT 1121.670 3.670 1149.810 4.280 ;
        RECT 1150.650 3.670 1178.790 4.280 ;
        RECT 1179.630 3.670 1207.770 4.280 ;
        RECT 1208.610 3.670 1236.750 4.280 ;
        RECT 1237.590 3.670 1265.730 4.280 ;
        RECT 1266.570 3.670 1294.710 4.280 ;
        RECT 1295.550 3.670 1323.690 4.280 ;
        RECT 1324.530 3.670 1352.670 4.280 ;
        RECT 1353.510 3.670 1381.650 4.280 ;
        RECT 1382.490 3.670 1410.630 4.280 ;
        RECT 1411.470 3.670 1439.610 4.280 ;
        RECT 1440.450 3.670 1468.590 4.280 ;
        RECT 1469.430 3.670 1497.570 4.280 ;
        RECT 1498.410 3.670 1526.550 4.280 ;
        RECT 1527.390 3.670 1555.530 4.280 ;
        RECT 1556.370 3.670 1584.510 4.280 ;
        RECT 1585.350 3.670 1613.490 4.280 ;
        RECT 1614.330 3.670 1642.470 4.280 ;
        RECT 1643.310 3.670 1671.450 4.280 ;
        RECT 1672.290 3.670 1700.430 4.280 ;
        RECT 1701.270 3.670 1729.410 4.280 ;
        RECT 1730.250 3.670 1758.390 4.280 ;
        RECT 1759.230 3.670 1787.370 4.280 ;
        RECT 1788.210 3.670 1816.350 4.280 ;
        RECT 1817.190 3.670 1845.330 4.280 ;
        RECT 1846.170 3.670 1874.310 4.280 ;
        RECT 1875.150 3.670 1903.290 4.280 ;
        RECT 1904.130 3.670 1932.270 4.280 ;
        RECT 1933.110 3.670 1961.250 4.280 ;
        RECT 1962.090 3.670 1990.230 4.280 ;
        RECT 1991.070 3.670 2019.210 4.280 ;
        RECT 2020.050 3.670 2048.190 4.280 ;
        RECT 2049.030 3.670 2077.170 4.280 ;
        RECT 2078.010 3.670 2106.150 4.280 ;
        RECT 2106.990 3.670 2135.130 4.280 ;
        RECT 2135.970 3.670 2164.110 4.280 ;
        RECT 2164.950 3.670 2193.090 4.280 ;
        RECT 2193.930 3.670 2222.070 4.280 ;
        RECT 2222.910 3.670 2251.050 4.280 ;
        RECT 2251.890 3.670 2280.030 4.280 ;
        RECT 2280.870 3.670 2309.010 4.280 ;
        RECT 2309.850 3.670 2337.990 4.280 ;
        RECT 2338.830 3.670 2366.970 4.280 ;
        RECT 2367.810 3.670 2395.950 4.280 ;
        RECT 2396.790 3.670 2424.930 4.280 ;
        RECT 2425.770 3.670 2453.910 4.280 ;
        RECT 2454.750 3.670 2471.020 4.280 ;
      LAYER met3 ;
        RECT 3.745 2690.440 2471.000 2703.845 ;
        RECT 4.400 2689.040 2471.000 2690.440 ;
        RECT 3.745 2683.640 2471.000 2689.040 ;
        RECT 3.745 2682.240 2470.600 2683.640 ;
        RECT 3.745 2663.240 2471.000 2682.240 ;
        RECT 4.400 2661.840 2471.000 2663.240 ;
        RECT 3.745 2657.120 2471.000 2661.840 ;
        RECT 3.745 2655.720 2470.600 2657.120 ;
        RECT 3.745 2636.040 2471.000 2655.720 ;
        RECT 4.400 2634.640 2471.000 2636.040 ;
        RECT 3.745 2630.600 2471.000 2634.640 ;
        RECT 3.745 2629.200 2470.600 2630.600 ;
        RECT 3.745 2608.840 2471.000 2629.200 ;
        RECT 4.400 2607.440 2471.000 2608.840 ;
        RECT 3.745 2604.080 2471.000 2607.440 ;
        RECT 3.745 2602.680 2470.600 2604.080 ;
        RECT 3.745 2581.640 2471.000 2602.680 ;
        RECT 4.400 2580.240 2471.000 2581.640 ;
        RECT 3.745 2577.560 2471.000 2580.240 ;
        RECT 3.745 2576.160 2470.600 2577.560 ;
        RECT 3.745 2554.440 2471.000 2576.160 ;
        RECT 4.400 2553.040 2471.000 2554.440 ;
        RECT 3.745 2551.040 2471.000 2553.040 ;
        RECT 3.745 2549.640 2470.600 2551.040 ;
        RECT 3.745 2527.240 2471.000 2549.640 ;
        RECT 4.400 2525.840 2471.000 2527.240 ;
        RECT 3.745 2524.520 2471.000 2525.840 ;
        RECT 3.745 2523.120 2470.600 2524.520 ;
        RECT 3.745 2500.040 2471.000 2523.120 ;
        RECT 4.400 2498.640 2471.000 2500.040 ;
        RECT 3.745 2498.000 2471.000 2498.640 ;
        RECT 3.745 2496.600 2470.600 2498.000 ;
        RECT 3.745 2472.840 2471.000 2496.600 ;
        RECT 4.400 2471.480 2471.000 2472.840 ;
        RECT 4.400 2471.440 2470.600 2471.480 ;
        RECT 3.745 2470.080 2470.600 2471.440 ;
        RECT 3.745 2445.640 2471.000 2470.080 ;
        RECT 4.400 2444.960 2471.000 2445.640 ;
        RECT 4.400 2444.240 2470.600 2444.960 ;
        RECT 3.745 2443.560 2470.600 2444.240 ;
        RECT 3.745 2418.440 2471.000 2443.560 ;
        RECT 4.400 2417.040 2470.600 2418.440 ;
        RECT 3.745 2391.920 2471.000 2417.040 ;
        RECT 3.745 2391.240 2470.600 2391.920 ;
        RECT 4.400 2390.520 2470.600 2391.240 ;
        RECT 4.400 2389.840 2471.000 2390.520 ;
        RECT 3.745 2365.400 2471.000 2389.840 ;
        RECT 3.745 2364.040 2470.600 2365.400 ;
        RECT 4.400 2364.000 2470.600 2364.040 ;
        RECT 4.400 2362.640 2471.000 2364.000 ;
        RECT 3.745 2338.880 2471.000 2362.640 ;
        RECT 3.745 2337.480 2470.600 2338.880 ;
        RECT 3.745 2336.840 2471.000 2337.480 ;
        RECT 4.400 2335.440 2471.000 2336.840 ;
        RECT 3.745 2312.360 2471.000 2335.440 ;
        RECT 3.745 2310.960 2470.600 2312.360 ;
        RECT 3.745 2309.640 2471.000 2310.960 ;
        RECT 4.400 2308.240 2471.000 2309.640 ;
        RECT 3.745 2285.840 2471.000 2308.240 ;
        RECT 3.745 2284.440 2470.600 2285.840 ;
        RECT 3.745 2282.440 2471.000 2284.440 ;
        RECT 4.400 2281.040 2471.000 2282.440 ;
        RECT 3.745 2259.320 2471.000 2281.040 ;
        RECT 3.745 2257.920 2470.600 2259.320 ;
        RECT 3.745 2255.240 2471.000 2257.920 ;
        RECT 4.400 2253.840 2471.000 2255.240 ;
        RECT 3.745 2232.800 2471.000 2253.840 ;
        RECT 3.745 2231.400 2470.600 2232.800 ;
        RECT 3.745 2228.040 2471.000 2231.400 ;
        RECT 4.400 2226.640 2471.000 2228.040 ;
        RECT 3.745 2206.280 2471.000 2226.640 ;
        RECT 3.745 2204.880 2470.600 2206.280 ;
        RECT 3.745 2200.840 2471.000 2204.880 ;
        RECT 4.400 2199.440 2471.000 2200.840 ;
        RECT 3.745 2179.760 2471.000 2199.440 ;
        RECT 3.745 2178.360 2470.600 2179.760 ;
        RECT 3.745 2173.640 2471.000 2178.360 ;
        RECT 4.400 2172.240 2471.000 2173.640 ;
        RECT 3.745 2153.240 2471.000 2172.240 ;
        RECT 3.745 2151.840 2470.600 2153.240 ;
        RECT 3.745 2146.440 2471.000 2151.840 ;
        RECT 4.400 2145.040 2471.000 2146.440 ;
        RECT 3.745 2126.720 2471.000 2145.040 ;
        RECT 3.745 2125.320 2470.600 2126.720 ;
        RECT 3.745 2119.240 2471.000 2125.320 ;
        RECT 4.400 2117.840 2471.000 2119.240 ;
        RECT 3.745 2100.200 2471.000 2117.840 ;
        RECT 3.745 2098.800 2470.600 2100.200 ;
        RECT 3.745 2092.040 2471.000 2098.800 ;
        RECT 4.400 2090.640 2471.000 2092.040 ;
        RECT 3.745 2073.680 2471.000 2090.640 ;
        RECT 3.745 2072.280 2470.600 2073.680 ;
        RECT 3.745 2064.840 2471.000 2072.280 ;
        RECT 4.400 2063.440 2471.000 2064.840 ;
        RECT 3.745 2047.160 2471.000 2063.440 ;
        RECT 3.745 2045.760 2470.600 2047.160 ;
        RECT 3.745 2037.640 2471.000 2045.760 ;
        RECT 4.400 2036.240 2471.000 2037.640 ;
        RECT 3.745 2020.640 2471.000 2036.240 ;
        RECT 3.745 2019.240 2470.600 2020.640 ;
        RECT 3.745 2010.440 2471.000 2019.240 ;
        RECT 4.400 2009.040 2471.000 2010.440 ;
        RECT 3.745 1994.120 2471.000 2009.040 ;
        RECT 3.745 1992.720 2470.600 1994.120 ;
        RECT 3.745 1983.240 2471.000 1992.720 ;
        RECT 4.400 1981.840 2471.000 1983.240 ;
        RECT 3.745 1967.600 2471.000 1981.840 ;
        RECT 3.745 1966.200 2470.600 1967.600 ;
        RECT 3.745 1956.040 2471.000 1966.200 ;
        RECT 4.400 1954.640 2471.000 1956.040 ;
        RECT 3.745 1941.080 2471.000 1954.640 ;
        RECT 3.745 1939.680 2470.600 1941.080 ;
        RECT 3.745 1928.840 2471.000 1939.680 ;
        RECT 4.400 1927.440 2471.000 1928.840 ;
        RECT 3.745 1914.560 2471.000 1927.440 ;
        RECT 3.745 1913.160 2470.600 1914.560 ;
        RECT 3.745 1901.640 2471.000 1913.160 ;
        RECT 4.400 1900.240 2471.000 1901.640 ;
        RECT 3.745 1888.040 2471.000 1900.240 ;
        RECT 3.745 1886.640 2470.600 1888.040 ;
        RECT 3.745 1874.440 2471.000 1886.640 ;
        RECT 4.400 1873.040 2471.000 1874.440 ;
        RECT 3.745 1861.520 2471.000 1873.040 ;
        RECT 3.745 1860.120 2470.600 1861.520 ;
        RECT 3.745 1847.240 2471.000 1860.120 ;
        RECT 4.400 1845.840 2471.000 1847.240 ;
        RECT 3.745 1835.000 2471.000 1845.840 ;
        RECT 3.745 1833.600 2470.600 1835.000 ;
        RECT 3.745 1820.040 2471.000 1833.600 ;
        RECT 4.400 1818.640 2471.000 1820.040 ;
        RECT 3.745 1808.480 2471.000 1818.640 ;
        RECT 3.745 1807.080 2470.600 1808.480 ;
        RECT 3.745 1792.840 2471.000 1807.080 ;
        RECT 4.400 1791.440 2471.000 1792.840 ;
        RECT 3.745 1781.960 2471.000 1791.440 ;
        RECT 3.745 1780.560 2470.600 1781.960 ;
        RECT 3.745 1765.640 2471.000 1780.560 ;
        RECT 4.400 1764.240 2471.000 1765.640 ;
        RECT 3.745 1755.440 2471.000 1764.240 ;
        RECT 3.745 1754.040 2470.600 1755.440 ;
        RECT 3.745 1738.440 2471.000 1754.040 ;
        RECT 4.400 1737.040 2471.000 1738.440 ;
        RECT 3.745 1728.920 2471.000 1737.040 ;
        RECT 3.745 1727.520 2470.600 1728.920 ;
        RECT 3.745 1711.240 2471.000 1727.520 ;
        RECT 4.400 1709.840 2471.000 1711.240 ;
        RECT 3.745 1702.400 2471.000 1709.840 ;
        RECT 3.745 1701.000 2470.600 1702.400 ;
        RECT 3.745 1684.040 2471.000 1701.000 ;
        RECT 4.400 1682.640 2471.000 1684.040 ;
        RECT 3.745 1675.880 2471.000 1682.640 ;
        RECT 3.745 1674.480 2470.600 1675.880 ;
        RECT 3.745 1656.840 2471.000 1674.480 ;
        RECT 4.400 1655.440 2471.000 1656.840 ;
        RECT 3.745 1649.360 2471.000 1655.440 ;
        RECT 3.745 1647.960 2470.600 1649.360 ;
        RECT 3.745 1629.640 2471.000 1647.960 ;
        RECT 4.400 1628.240 2471.000 1629.640 ;
        RECT 3.745 1622.840 2471.000 1628.240 ;
        RECT 3.745 1621.440 2470.600 1622.840 ;
        RECT 3.745 1602.440 2471.000 1621.440 ;
        RECT 4.400 1601.040 2471.000 1602.440 ;
        RECT 3.745 1596.320 2471.000 1601.040 ;
        RECT 3.745 1594.920 2470.600 1596.320 ;
        RECT 3.745 1575.240 2471.000 1594.920 ;
        RECT 4.400 1573.840 2471.000 1575.240 ;
        RECT 3.745 1569.800 2471.000 1573.840 ;
        RECT 3.745 1568.400 2470.600 1569.800 ;
        RECT 3.745 1548.040 2471.000 1568.400 ;
        RECT 4.400 1546.640 2471.000 1548.040 ;
        RECT 3.745 1543.280 2471.000 1546.640 ;
        RECT 3.745 1541.880 2470.600 1543.280 ;
        RECT 3.745 1520.840 2471.000 1541.880 ;
        RECT 4.400 1519.440 2471.000 1520.840 ;
        RECT 3.745 1516.760 2471.000 1519.440 ;
        RECT 3.745 1515.360 2470.600 1516.760 ;
        RECT 3.745 1493.640 2471.000 1515.360 ;
        RECT 4.400 1492.240 2471.000 1493.640 ;
        RECT 3.745 1490.240 2471.000 1492.240 ;
        RECT 3.745 1488.840 2470.600 1490.240 ;
        RECT 3.745 1466.440 2471.000 1488.840 ;
        RECT 4.400 1465.040 2471.000 1466.440 ;
        RECT 3.745 1463.720 2471.000 1465.040 ;
        RECT 3.745 1462.320 2470.600 1463.720 ;
        RECT 3.745 1439.240 2471.000 1462.320 ;
        RECT 4.400 1437.840 2471.000 1439.240 ;
        RECT 3.745 1437.200 2471.000 1437.840 ;
        RECT 3.745 1435.800 2470.600 1437.200 ;
        RECT 3.745 1412.040 2471.000 1435.800 ;
        RECT 4.400 1410.680 2471.000 1412.040 ;
        RECT 4.400 1410.640 2470.600 1410.680 ;
        RECT 3.745 1409.280 2470.600 1410.640 ;
        RECT 3.745 1384.840 2471.000 1409.280 ;
        RECT 4.400 1384.160 2471.000 1384.840 ;
        RECT 4.400 1383.440 2470.600 1384.160 ;
        RECT 3.745 1382.760 2470.600 1383.440 ;
        RECT 3.745 1357.640 2471.000 1382.760 ;
        RECT 4.400 1356.240 2470.600 1357.640 ;
        RECT 3.745 1331.120 2471.000 1356.240 ;
        RECT 3.745 1330.440 2470.600 1331.120 ;
        RECT 4.400 1329.720 2470.600 1330.440 ;
        RECT 4.400 1329.040 2471.000 1329.720 ;
        RECT 3.745 1304.600 2471.000 1329.040 ;
        RECT 3.745 1303.240 2470.600 1304.600 ;
        RECT 4.400 1303.200 2470.600 1303.240 ;
        RECT 4.400 1301.840 2471.000 1303.200 ;
        RECT 3.745 1278.080 2471.000 1301.840 ;
        RECT 3.745 1276.680 2470.600 1278.080 ;
        RECT 3.745 1276.040 2471.000 1276.680 ;
        RECT 4.400 1274.640 2471.000 1276.040 ;
        RECT 3.745 1251.560 2471.000 1274.640 ;
        RECT 3.745 1250.160 2470.600 1251.560 ;
        RECT 3.745 1248.840 2471.000 1250.160 ;
        RECT 4.400 1247.440 2471.000 1248.840 ;
        RECT 3.745 1225.040 2471.000 1247.440 ;
        RECT 3.745 1223.640 2470.600 1225.040 ;
        RECT 3.745 1221.640 2471.000 1223.640 ;
        RECT 4.400 1220.240 2471.000 1221.640 ;
        RECT 3.745 1198.520 2471.000 1220.240 ;
        RECT 3.745 1197.120 2470.600 1198.520 ;
        RECT 3.745 1194.440 2471.000 1197.120 ;
        RECT 4.400 1193.040 2471.000 1194.440 ;
        RECT 3.745 1172.000 2471.000 1193.040 ;
        RECT 3.745 1170.600 2470.600 1172.000 ;
        RECT 3.745 1167.240 2471.000 1170.600 ;
        RECT 4.400 1165.840 2471.000 1167.240 ;
        RECT 3.745 1145.480 2471.000 1165.840 ;
        RECT 3.745 1144.080 2470.600 1145.480 ;
        RECT 3.745 1140.040 2471.000 1144.080 ;
        RECT 4.400 1138.640 2471.000 1140.040 ;
        RECT 3.745 1118.960 2471.000 1138.640 ;
        RECT 3.745 1117.560 2470.600 1118.960 ;
        RECT 3.745 1112.840 2471.000 1117.560 ;
        RECT 4.400 1111.440 2471.000 1112.840 ;
        RECT 3.745 1092.440 2471.000 1111.440 ;
        RECT 3.745 1091.040 2470.600 1092.440 ;
        RECT 3.745 1085.640 2471.000 1091.040 ;
        RECT 4.400 1084.240 2471.000 1085.640 ;
        RECT 3.745 1065.920 2471.000 1084.240 ;
        RECT 3.745 1064.520 2470.600 1065.920 ;
        RECT 3.745 1058.440 2471.000 1064.520 ;
        RECT 4.400 1057.040 2471.000 1058.440 ;
        RECT 3.745 1039.400 2471.000 1057.040 ;
        RECT 3.745 1038.000 2470.600 1039.400 ;
        RECT 3.745 1031.240 2471.000 1038.000 ;
        RECT 4.400 1029.840 2471.000 1031.240 ;
        RECT 3.745 1012.880 2471.000 1029.840 ;
        RECT 3.745 1011.480 2470.600 1012.880 ;
        RECT 3.745 1004.040 2471.000 1011.480 ;
        RECT 4.400 1002.640 2471.000 1004.040 ;
        RECT 3.745 986.360 2471.000 1002.640 ;
        RECT 3.745 984.960 2470.600 986.360 ;
        RECT 3.745 976.840 2471.000 984.960 ;
        RECT 4.400 975.440 2471.000 976.840 ;
        RECT 3.745 959.840 2471.000 975.440 ;
        RECT 3.745 958.440 2470.600 959.840 ;
        RECT 3.745 949.640 2471.000 958.440 ;
        RECT 4.400 948.240 2471.000 949.640 ;
        RECT 3.745 933.320 2471.000 948.240 ;
        RECT 3.745 931.920 2470.600 933.320 ;
        RECT 3.745 922.440 2471.000 931.920 ;
        RECT 4.400 921.040 2471.000 922.440 ;
        RECT 3.745 906.800 2471.000 921.040 ;
        RECT 3.745 905.400 2470.600 906.800 ;
        RECT 3.745 895.240 2471.000 905.400 ;
        RECT 4.400 893.840 2471.000 895.240 ;
        RECT 3.745 880.280 2471.000 893.840 ;
        RECT 3.745 878.880 2470.600 880.280 ;
        RECT 3.745 868.040 2471.000 878.880 ;
        RECT 4.400 866.640 2471.000 868.040 ;
        RECT 3.745 853.760 2471.000 866.640 ;
        RECT 3.745 852.360 2470.600 853.760 ;
        RECT 3.745 840.840 2471.000 852.360 ;
        RECT 4.400 839.440 2471.000 840.840 ;
        RECT 3.745 827.240 2471.000 839.440 ;
        RECT 3.745 825.840 2470.600 827.240 ;
        RECT 3.745 813.640 2471.000 825.840 ;
        RECT 4.400 812.240 2471.000 813.640 ;
        RECT 3.745 800.720 2471.000 812.240 ;
        RECT 3.745 799.320 2470.600 800.720 ;
        RECT 3.745 786.440 2471.000 799.320 ;
        RECT 4.400 785.040 2471.000 786.440 ;
        RECT 3.745 774.200 2471.000 785.040 ;
        RECT 3.745 772.800 2470.600 774.200 ;
        RECT 3.745 759.240 2471.000 772.800 ;
        RECT 4.400 757.840 2471.000 759.240 ;
        RECT 3.745 747.680 2471.000 757.840 ;
        RECT 3.745 746.280 2470.600 747.680 ;
        RECT 3.745 732.040 2471.000 746.280 ;
        RECT 4.400 730.640 2471.000 732.040 ;
        RECT 3.745 721.160 2471.000 730.640 ;
        RECT 3.745 719.760 2470.600 721.160 ;
        RECT 3.745 704.840 2471.000 719.760 ;
        RECT 4.400 703.440 2471.000 704.840 ;
        RECT 3.745 694.640 2471.000 703.440 ;
        RECT 3.745 693.240 2470.600 694.640 ;
        RECT 3.745 677.640 2471.000 693.240 ;
        RECT 4.400 676.240 2471.000 677.640 ;
        RECT 3.745 668.120 2471.000 676.240 ;
        RECT 3.745 666.720 2470.600 668.120 ;
        RECT 3.745 650.440 2471.000 666.720 ;
        RECT 4.400 649.040 2471.000 650.440 ;
        RECT 3.745 641.600 2471.000 649.040 ;
        RECT 3.745 640.200 2470.600 641.600 ;
        RECT 3.745 623.240 2471.000 640.200 ;
        RECT 4.400 621.840 2471.000 623.240 ;
        RECT 3.745 615.080 2471.000 621.840 ;
        RECT 3.745 613.680 2470.600 615.080 ;
        RECT 3.745 596.040 2471.000 613.680 ;
        RECT 4.400 594.640 2471.000 596.040 ;
        RECT 3.745 588.560 2471.000 594.640 ;
        RECT 3.745 587.160 2470.600 588.560 ;
        RECT 3.745 568.840 2471.000 587.160 ;
        RECT 4.400 567.440 2471.000 568.840 ;
        RECT 3.745 562.040 2471.000 567.440 ;
        RECT 3.745 560.640 2470.600 562.040 ;
        RECT 3.745 541.640 2471.000 560.640 ;
        RECT 4.400 540.240 2471.000 541.640 ;
        RECT 3.745 535.520 2471.000 540.240 ;
        RECT 3.745 534.120 2470.600 535.520 ;
        RECT 3.745 514.440 2471.000 534.120 ;
        RECT 4.400 513.040 2471.000 514.440 ;
        RECT 3.745 509.000 2471.000 513.040 ;
        RECT 3.745 507.600 2470.600 509.000 ;
        RECT 3.745 487.240 2471.000 507.600 ;
        RECT 4.400 485.840 2471.000 487.240 ;
        RECT 3.745 482.480 2471.000 485.840 ;
        RECT 3.745 481.080 2470.600 482.480 ;
        RECT 3.745 460.040 2471.000 481.080 ;
        RECT 4.400 458.640 2471.000 460.040 ;
        RECT 3.745 455.960 2471.000 458.640 ;
        RECT 3.745 454.560 2470.600 455.960 ;
        RECT 3.745 432.840 2471.000 454.560 ;
        RECT 4.400 431.440 2471.000 432.840 ;
        RECT 3.745 429.440 2471.000 431.440 ;
        RECT 3.745 428.040 2470.600 429.440 ;
        RECT 3.745 405.640 2471.000 428.040 ;
        RECT 4.400 404.240 2471.000 405.640 ;
        RECT 3.745 402.920 2471.000 404.240 ;
        RECT 3.745 401.520 2470.600 402.920 ;
        RECT 3.745 378.440 2471.000 401.520 ;
        RECT 4.400 377.040 2471.000 378.440 ;
        RECT 3.745 376.400 2471.000 377.040 ;
        RECT 3.745 375.000 2470.600 376.400 ;
        RECT 3.745 351.240 2471.000 375.000 ;
        RECT 4.400 349.880 2471.000 351.240 ;
        RECT 4.400 349.840 2470.600 349.880 ;
        RECT 3.745 348.480 2470.600 349.840 ;
        RECT 3.745 324.040 2471.000 348.480 ;
        RECT 4.400 323.360 2471.000 324.040 ;
        RECT 4.400 322.640 2470.600 323.360 ;
        RECT 3.745 321.960 2470.600 322.640 ;
        RECT 3.745 296.840 2471.000 321.960 ;
        RECT 4.400 295.440 2470.600 296.840 ;
        RECT 3.745 270.320 2471.000 295.440 ;
        RECT 3.745 269.640 2470.600 270.320 ;
        RECT 4.400 268.920 2470.600 269.640 ;
        RECT 4.400 268.240 2471.000 268.920 ;
        RECT 3.745 243.800 2471.000 268.240 ;
        RECT 3.745 242.440 2470.600 243.800 ;
        RECT 4.400 242.400 2470.600 242.440 ;
        RECT 4.400 241.040 2471.000 242.400 ;
        RECT 3.745 217.280 2471.000 241.040 ;
        RECT 3.745 215.880 2470.600 217.280 ;
        RECT 3.745 215.240 2471.000 215.880 ;
        RECT 4.400 213.840 2471.000 215.240 ;
        RECT 3.745 190.760 2471.000 213.840 ;
        RECT 3.745 189.360 2470.600 190.760 ;
        RECT 3.745 188.040 2471.000 189.360 ;
        RECT 4.400 186.640 2471.000 188.040 ;
        RECT 3.745 164.240 2471.000 186.640 ;
        RECT 3.745 162.840 2470.600 164.240 ;
        RECT 3.745 160.840 2471.000 162.840 ;
        RECT 4.400 159.440 2471.000 160.840 ;
        RECT 3.745 137.720 2471.000 159.440 ;
        RECT 3.745 136.320 2470.600 137.720 ;
        RECT 3.745 133.640 2471.000 136.320 ;
        RECT 4.400 132.240 2471.000 133.640 ;
        RECT 3.745 111.200 2471.000 132.240 ;
        RECT 3.745 109.800 2470.600 111.200 ;
        RECT 3.745 106.440 2471.000 109.800 ;
        RECT 4.400 105.040 2471.000 106.440 ;
        RECT 3.745 84.680 2471.000 105.040 ;
        RECT 3.745 83.280 2470.600 84.680 ;
        RECT 3.745 79.240 2471.000 83.280 ;
        RECT 4.400 77.840 2471.000 79.240 ;
        RECT 3.745 58.160 2471.000 77.840 ;
        RECT 3.745 56.760 2470.600 58.160 ;
        RECT 3.745 52.040 2471.000 56.760 ;
        RECT 4.400 50.640 2471.000 52.040 ;
        RECT 3.745 31.640 2471.000 50.640 ;
        RECT 3.745 30.240 2470.600 31.640 ;
        RECT 3.745 24.840 2471.000 30.240 ;
        RECT 4.400 23.440 2471.000 24.840 ;
        RECT 3.745 10.715 2471.000 23.440 ;
      LAYER met4 ;
        RECT 44.720 170.965 61.720 2672.240 ;
        RECT 65.720 2618.485 123.520 2672.240 ;
        RECT 127.520 2618.485 175.720 2672.240 ;
        RECT 65.720 2402.515 175.720 2618.485 ;
        RECT 65.720 2400.740 123.520 2402.515 ;
        RECT 65.720 2367.140 66.520 2400.740 ;
        RECT 70.520 2367.140 118.720 2400.740 ;
        RECT 122.720 2367.140 123.520 2400.740 ;
        RECT 65.720 2364.685 123.520 2367.140 ;
        RECT 127.520 2364.685 175.720 2402.515 ;
        RECT 65.720 2089.555 175.720 2364.685 ;
        RECT 65.720 2085.740 123.520 2089.555 ;
        RECT 65.720 2052.140 66.520 2085.740 ;
        RECT 70.520 2052.140 118.720 2085.740 ;
        RECT 122.720 2052.140 123.520 2085.740 ;
        RECT 65.720 2049.685 123.520 2052.140 ;
        RECT 127.520 2049.685 175.720 2089.555 ;
        RECT 65.720 1774.555 175.720 2049.685 ;
        RECT 65.720 1770.740 123.520 1774.555 ;
        RECT 65.720 1737.140 66.520 1770.740 ;
        RECT 70.520 1737.140 118.720 1770.740 ;
        RECT 122.720 1737.140 123.520 1770.740 ;
        RECT 65.720 1734.685 123.520 1737.140 ;
        RECT 127.520 1734.685 175.720 1774.555 ;
        RECT 65.720 1459.555 175.720 1734.685 ;
        RECT 65.720 1455.740 123.520 1459.555 ;
        RECT 65.720 1422.140 66.520 1455.740 ;
        RECT 70.520 1422.140 118.720 1455.740 ;
        RECT 122.720 1422.140 123.520 1455.740 ;
        RECT 65.720 1419.685 123.520 1422.140 ;
        RECT 127.520 1419.685 175.720 1459.555 ;
        RECT 65.720 1144.555 175.720 1419.685 ;
        RECT 65.720 1140.740 123.520 1144.555 ;
        RECT 65.720 1107.140 66.520 1140.740 ;
        RECT 70.520 1107.140 118.720 1140.740 ;
        RECT 122.720 1107.140 123.520 1140.740 ;
        RECT 65.720 1104.685 123.520 1107.140 ;
        RECT 127.520 1104.685 175.720 1144.555 ;
        RECT 65.720 829.555 175.720 1104.685 ;
        RECT 65.720 825.740 123.520 829.555 ;
        RECT 65.720 792.140 66.520 825.740 ;
        RECT 70.520 792.140 118.720 825.740 ;
        RECT 122.720 792.140 123.520 825.740 ;
        RECT 65.720 789.685 123.520 792.140 ;
        RECT 127.520 789.685 175.720 829.555 ;
        RECT 65.720 514.555 175.720 789.685 ;
        RECT 65.720 510.740 123.520 514.555 ;
        RECT 65.720 477.140 66.520 510.740 ;
        RECT 70.520 477.140 118.720 510.740 ;
        RECT 122.720 477.140 123.520 510.740 ;
        RECT 65.720 474.685 123.520 477.140 ;
        RECT 127.520 474.685 175.720 514.555 ;
        RECT 65.720 199.555 175.720 474.685 ;
        RECT 65.720 195.740 123.520 199.555 ;
        RECT 65.720 170.965 66.520 195.740 ;
        RECT 70.520 170.965 118.720 195.740 ;
        RECT 122.720 170.965 123.520 195.740 ;
        RECT 127.520 170.965 175.720 199.555 ;
        RECT 44.720 67.875 175.720 170.965 ;
        RECT 44.720 40.640 61.720 67.875 ;
        RECT 65.720 40.640 123.520 67.875 ;
        RECT 127.520 40.640 175.720 67.875 ;
        RECT 179.720 40.640 180.520 2672.240 ;
        RECT 184.520 2655.885 237.520 2672.240 ;
        RECT 241.520 2655.885 289.720 2672.240 ;
        RECT 293.720 2655.885 294.520 2672.240 ;
        RECT 298.520 2655.885 346.720 2672.240 ;
        RECT 350.720 2655.885 351.520 2672.240 ;
        RECT 355.520 2655.885 403.720 2672.240 ;
        RECT 407.720 2655.885 460.720 2672.240 ;
        RECT 184.520 2421.555 460.720 2655.885 ;
        RECT 184.520 2400.740 237.520 2421.555 ;
        RECT 184.520 2367.140 232.720 2400.740 ;
        RECT 236.720 2367.140 237.520 2400.740 ;
        RECT 184.520 2343.605 237.520 2367.140 ;
        RECT 241.520 2343.605 289.720 2421.555 ;
        RECT 293.720 2343.605 294.520 2421.555 ;
        RECT 298.520 2343.605 346.720 2421.555 ;
        RECT 350.720 2343.605 351.520 2421.555 ;
        RECT 355.520 2343.605 403.720 2421.555 ;
        RECT 407.720 2400.740 460.720 2421.555 ;
        RECT 407.720 2367.140 408.520 2400.740 ;
        RECT 412.520 2367.140 460.720 2400.740 ;
        RECT 407.720 2343.605 460.720 2367.140 ;
        RECT 184.520 2113.355 460.720 2343.605 ;
        RECT 184.520 2085.740 237.520 2113.355 ;
        RECT 184.520 2052.140 232.720 2085.740 ;
        RECT 236.720 2052.140 237.520 2085.740 ;
        RECT 184.520 2028.605 237.520 2052.140 ;
        RECT 241.520 2028.605 289.720 2113.355 ;
        RECT 293.720 2028.605 294.520 2113.355 ;
        RECT 298.520 2028.605 346.720 2113.355 ;
        RECT 350.720 2028.605 351.520 2113.355 ;
        RECT 355.520 2028.605 403.720 2113.355 ;
        RECT 407.720 2085.740 460.720 2113.355 ;
        RECT 407.720 2052.140 408.520 2085.740 ;
        RECT 412.520 2052.140 460.720 2085.740 ;
        RECT 407.720 2028.605 460.720 2052.140 ;
        RECT 184.520 1798.355 460.720 2028.605 ;
        RECT 184.520 1770.740 237.520 1798.355 ;
        RECT 184.520 1737.140 232.720 1770.740 ;
        RECT 236.720 1737.140 237.520 1770.740 ;
        RECT 184.520 1713.605 237.520 1737.140 ;
        RECT 241.520 1713.605 289.720 1798.355 ;
        RECT 293.720 1713.605 294.520 1798.355 ;
        RECT 298.520 1713.605 346.720 1798.355 ;
        RECT 350.720 1713.605 351.520 1798.355 ;
        RECT 355.520 1713.605 403.720 1798.355 ;
        RECT 407.720 1770.740 460.720 1798.355 ;
        RECT 407.720 1737.140 408.520 1770.740 ;
        RECT 412.520 1737.140 460.720 1770.740 ;
        RECT 407.720 1713.605 460.720 1737.140 ;
        RECT 184.520 1483.355 460.720 1713.605 ;
        RECT 184.520 1455.740 237.520 1483.355 ;
        RECT 184.520 1422.140 232.720 1455.740 ;
        RECT 236.720 1422.140 237.520 1455.740 ;
        RECT 184.520 1398.605 237.520 1422.140 ;
        RECT 241.520 1398.605 289.720 1483.355 ;
        RECT 293.720 1398.605 294.520 1483.355 ;
        RECT 298.520 1398.605 346.720 1483.355 ;
        RECT 350.720 1398.605 351.520 1483.355 ;
        RECT 355.520 1398.605 403.720 1483.355 ;
        RECT 407.720 1455.740 460.720 1483.355 ;
        RECT 407.720 1422.140 408.520 1455.740 ;
        RECT 412.520 1422.140 460.720 1455.740 ;
        RECT 407.720 1398.605 460.720 1422.140 ;
        RECT 184.520 1168.355 460.720 1398.605 ;
        RECT 184.520 1140.740 237.520 1168.355 ;
        RECT 184.520 1107.140 232.720 1140.740 ;
        RECT 236.720 1107.140 237.520 1140.740 ;
        RECT 184.520 1083.605 237.520 1107.140 ;
        RECT 241.520 1083.605 289.720 1168.355 ;
        RECT 293.720 1083.605 294.520 1168.355 ;
        RECT 298.520 1083.605 346.720 1168.355 ;
        RECT 350.720 1083.605 351.520 1168.355 ;
        RECT 355.520 1083.605 403.720 1168.355 ;
        RECT 407.720 1140.740 460.720 1168.355 ;
        RECT 407.720 1107.140 408.520 1140.740 ;
        RECT 412.520 1107.140 460.720 1140.740 ;
        RECT 407.720 1083.605 460.720 1107.140 ;
        RECT 184.520 853.355 460.720 1083.605 ;
        RECT 184.520 825.740 237.520 853.355 ;
        RECT 184.520 792.140 232.720 825.740 ;
        RECT 236.720 792.140 237.520 825.740 ;
        RECT 184.520 768.605 237.520 792.140 ;
        RECT 241.520 768.605 289.720 853.355 ;
        RECT 293.720 768.605 294.520 853.355 ;
        RECT 298.520 768.605 346.720 853.355 ;
        RECT 350.720 768.605 351.520 853.355 ;
        RECT 355.520 768.605 403.720 853.355 ;
        RECT 407.720 825.740 460.720 853.355 ;
        RECT 407.720 792.140 408.520 825.740 ;
        RECT 412.520 792.140 460.720 825.740 ;
        RECT 407.720 768.605 460.720 792.140 ;
        RECT 184.520 538.355 460.720 768.605 ;
        RECT 184.520 510.740 237.520 538.355 ;
        RECT 184.520 477.140 232.720 510.740 ;
        RECT 236.720 477.140 237.520 510.740 ;
        RECT 184.520 453.605 237.520 477.140 ;
        RECT 241.520 453.605 289.720 538.355 ;
        RECT 293.720 453.605 294.520 538.355 ;
        RECT 298.520 453.605 346.720 538.355 ;
        RECT 350.720 453.605 351.520 538.355 ;
        RECT 355.520 453.605 403.720 538.355 ;
        RECT 407.720 510.740 460.720 538.355 ;
        RECT 407.720 477.140 408.520 510.740 ;
        RECT 412.520 477.140 460.720 510.740 ;
        RECT 407.720 453.605 460.720 477.140 ;
        RECT 184.520 223.355 460.720 453.605 ;
        RECT 184.520 195.740 237.520 223.355 ;
        RECT 184.520 162.540 232.720 195.740 ;
        RECT 236.720 162.540 237.520 195.740 ;
        RECT 184.520 40.640 237.520 162.540 ;
        RECT 241.520 164.845 289.720 223.355 ;
        RECT 293.720 164.845 294.520 223.355 ;
        RECT 298.520 164.845 346.720 223.355 ;
        RECT 350.720 164.845 351.520 223.355 ;
        RECT 355.520 164.845 403.720 223.355 ;
        RECT 241.520 67.875 403.720 164.845 ;
        RECT 241.520 40.640 289.720 67.875 ;
        RECT 293.720 40.640 294.520 67.875 ;
        RECT 298.520 40.640 346.720 67.875 ;
        RECT 350.720 40.640 351.520 67.875 ;
        RECT 355.520 40.640 403.720 67.875 ;
        RECT 407.720 195.740 460.720 223.355 ;
        RECT 407.720 162.540 408.520 195.740 ;
        RECT 412.520 162.540 460.720 195.740 ;
        RECT 407.720 40.640 460.720 162.540 ;
        RECT 464.720 40.640 465.520 2672.240 ;
        RECT 469.520 2655.885 522.520 2672.240 ;
        RECT 526.520 2655.885 574.720 2672.240 ;
        RECT 578.720 2655.885 579.520 2672.240 ;
        RECT 583.520 2655.885 631.720 2672.240 ;
        RECT 635.720 2655.885 636.520 2672.240 ;
        RECT 640.520 2655.885 688.720 2672.240 ;
        RECT 692.720 2655.885 745.720 2672.240 ;
        RECT 469.520 2421.555 745.720 2655.885 ;
        RECT 469.520 2400.740 522.520 2421.555 ;
        RECT 469.520 2367.140 517.720 2400.740 ;
        RECT 521.720 2367.140 522.520 2400.740 ;
        RECT 469.520 2343.605 522.520 2367.140 ;
        RECT 526.520 2343.605 574.720 2421.555 ;
        RECT 578.720 2343.605 579.520 2421.555 ;
        RECT 583.520 2343.605 631.720 2421.555 ;
        RECT 635.720 2343.605 636.520 2421.555 ;
        RECT 640.520 2343.605 688.720 2421.555 ;
        RECT 692.720 2400.740 745.720 2421.555 ;
        RECT 692.720 2367.140 693.520 2400.740 ;
        RECT 697.520 2367.140 745.720 2400.740 ;
        RECT 692.720 2343.605 745.720 2367.140 ;
        RECT 469.520 2113.355 745.720 2343.605 ;
        RECT 469.520 2085.740 522.520 2113.355 ;
        RECT 469.520 2052.140 517.720 2085.740 ;
        RECT 521.720 2052.140 522.520 2085.740 ;
        RECT 469.520 2028.605 522.520 2052.140 ;
        RECT 526.520 2028.605 574.720 2113.355 ;
        RECT 578.720 2028.605 579.520 2113.355 ;
        RECT 583.520 2028.605 631.720 2113.355 ;
        RECT 635.720 2028.605 636.520 2113.355 ;
        RECT 640.520 2028.605 688.720 2113.355 ;
        RECT 692.720 2085.740 745.720 2113.355 ;
        RECT 692.720 2052.140 693.520 2085.740 ;
        RECT 697.520 2052.140 745.720 2085.740 ;
        RECT 692.720 2028.605 745.720 2052.140 ;
        RECT 469.520 1798.355 745.720 2028.605 ;
        RECT 469.520 1770.740 522.520 1798.355 ;
        RECT 469.520 1737.140 517.720 1770.740 ;
        RECT 521.720 1737.140 522.520 1770.740 ;
        RECT 469.520 1713.605 522.520 1737.140 ;
        RECT 526.520 1713.605 574.720 1798.355 ;
        RECT 578.720 1713.605 579.520 1798.355 ;
        RECT 583.520 1713.605 631.720 1798.355 ;
        RECT 635.720 1713.605 636.520 1798.355 ;
        RECT 640.520 1713.605 688.720 1798.355 ;
        RECT 692.720 1770.740 745.720 1798.355 ;
        RECT 692.720 1737.140 693.520 1770.740 ;
        RECT 697.520 1737.140 745.720 1770.740 ;
        RECT 692.720 1713.605 745.720 1737.140 ;
        RECT 469.520 1483.355 745.720 1713.605 ;
        RECT 469.520 1455.740 522.520 1483.355 ;
        RECT 469.520 1422.140 517.720 1455.740 ;
        RECT 521.720 1422.140 522.520 1455.740 ;
        RECT 469.520 1398.605 522.520 1422.140 ;
        RECT 526.520 1398.605 574.720 1483.355 ;
        RECT 578.720 1398.605 579.520 1483.355 ;
        RECT 583.520 1398.605 631.720 1483.355 ;
        RECT 635.720 1398.605 636.520 1483.355 ;
        RECT 640.520 1398.605 688.720 1483.355 ;
        RECT 692.720 1455.740 745.720 1483.355 ;
        RECT 692.720 1422.140 693.520 1455.740 ;
        RECT 697.520 1422.140 745.720 1455.740 ;
        RECT 692.720 1398.605 745.720 1422.140 ;
        RECT 469.520 1168.355 745.720 1398.605 ;
        RECT 469.520 1140.740 522.520 1168.355 ;
        RECT 469.520 1107.140 517.720 1140.740 ;
        RECT 521.720 1107.140 522.520 1140.740 ;
        RECT 469.520 1083.605 522.520 1107.140 ;
        RECT 526.520 1083.605 574.720 1168.355 ;
        RECT 578.720 1083.605 579.520 1168.355 ;
        RECT 583.520 1083.605 631.720 1168.355 ;
        RECT 635.720 1083.605 636.520 1168.355 ;
        RECT 640.520 1083.605 688.720 1168.355 ;
        RECT 692.720 1140.740 745.720 1168.355 ;
        RECT 692.720 1107.140 693.520 1140.740 ;
        RECT 697.520 1107.140 745.720 1140.740 ;
        RECT 692.720 1083.605 745.720 1107.140 ;
        RECT 469.520 853.355 745.720 1083.605 ;
        RECT 469.520 825.740 522.520 853.355 ;
        RECT 469.520 792.140 517.720 825.740 ;
        RECT 521.720 792.140 522.520 825.740 ;
        RECT 469.520 768.605 522.520 792.140 ;
        RECT 526.520 768.605 574.720 853.355 ;
        RECT 578.720 768.605 579.520 853.355 ;
        RECT 583.520 768.605 631.720 853.355 ;
        RECT 635.720 768.605 636.520 853.355 ;
        RECT 640.520 768.605 688.720 853.355 ;
        RECT 692.720 825.740 745.720 853.355 ;
        RECT 692.720 792.140 693.520 825.740 ;
        RECT 697.520 792.140 745.720 825.740 ;
        RECT 692.720 768.605 745.720 792.140 ;
        RECT 469.520 538.355 745.720 768.605 ;
        RECT 469.520 510.740 522.520 538.355 ;
        RECT 469.520 477.140 517.720 510.740 ;
        RECT 521.720 477.140 522.520 510.740 ;
        RECT 469.520 453.605 522.520 477.140 ;
        RECT 526.520 453.605 574.720 538.355 ;
        RECT 578.720 453.605 579.520 538.355 ;
        RECT 583.520 453.605 631.720 538.355 ;
        RECT 635.720 453.605 636.520 538.355 ;
        RECT 640.520 453.605 688.720 538.355 ;
        RECT 692.720 510.740 745.720 538.355 ;
        RECT 692.720 477.140 693.520 510.740 ;
        RECT 697.520 477.140 745.720 510.740 ;
        RECT 692.720 453.605 745.720 477.140 ;
        RECT 469.520 223.355 745.720 453.605 ;
        RECT 469.520 195.740 522.520 223.355 ;
        RECT 469.520 162.540 517.720 195.740 ;
        RECT 521.720 162.540 522.520 195.740 ;
        RECT 469.520 40.640 522.520 162.540 ;
        RECT 526.520 164.845 574.720 223.355 ;
        RECT 578.720 164.845 579.520 223.355 ;
        RECT 583.520 164.845 631.720 223.355 ;
        RECT 635.720 164.845 636.520 223.355 ;
        RECT 640.520 164.845 688.720 223.355 ;
        RECT 526.520 67.875 688.720 164.845 ;
        RECT 526.520 40.640 574.720 67.875 ;
        RECT 578.720 40.640 579.520 67.875 ;
        RECT 583.520 40.640 631.720 67.875 ;
        RECT 635.720 40.640 636.520 67.875 ;
        RECT 640.520 40.640 688.720 67.875 ;
        RECT 692.720 195.740 745.720 223.355 ;
        RECT 692.720 162.540 693.520 195.740 ;
        RECT 697.520 162.540 745.720 195.740 ;
        RECT 692.720 40.640 745.720 162.540 ;
        RECT 749.720 40.640 750.520 2672.240 ;
        RECT 754.520 2655.885 807.520 2672.240 ;
        RECT 811.520 2655.885 859.720 2672.240 ;
        RECT 863.720 2655.885 864.520 2672.240 ;
        RECT 868.520 2655.885 916.720 2672.240 ;
        RECT 920.720 2655.885 921.520 2672.240 ;
        RECT 925.520 2655.885 973.720 2672.240 ;
        RECT 977.720 2655.885 1030.720 2672.240 ;
        RECT 754.520 2421.555 1030.720 2655.885 ;
        RECT 754.520 2400.740 807.520 2421.555 ;
        RECT 754.520 2367.140 802.720 2400.740 ;
        RECT 806.720 2367.140 807.520 2400.740 ;
        RECT 754.520 2343.605 807.520 2367.140 ;
        RECT 811.520 2343.605 859.720 2421.555 ;
        RECT 863.720 2343.605 864.520 2421.555 ;
        RECT 868.520 2343.605 916.720 2421.555 ;
        RECT 920.720 2343.605 921.520 2421.555 ;
        RECT 925.520 2343.605 973.720 2421.555 ;
        RECT 977.720 2400.740 1030.720 2421.555 ;
        RECT 977.720 2367.140 978.520 2400.740 ;
        RECT 982.520 2367.140 1030.720 2400.740 ;
        RECT 977.720 2343.605 1030.720 2367.140 ;
        RECT 754.520 2113.355 1030.720 2343.605 ;
        RECT 754.520 2085.740 807.520 2113.355 ;
        RECT 754.520 2052.140 802.720 2085.740 ;
        RECT 806.720 2052.140 807.520 2085.740 ;
        RECT 754.520 2028.605 807.520 2052.140 ;
        RECT 811.520 2028.605 859.720 2113.355 ;
        RECT 863.720 2028.605 864.520 2113.355 ;
        RECT 868.520 2028.605 916.720 2113.355 ;
        RECT 920.720 2028.605 921.520 2113.355 ;
        RECT 925.520 2028.605 973.720 2113.355 ;
        RECT 977.720 2085.740 1030.720 2113.355 ;
        RECT 977.720 2052.140 978.520 2085.740 ;
        RECT 982.520 2052.140 1030.720 2085.740 ;
        RECT 977.720 2028.605 1030.720 2052.140 ;
        RECT 754.520 1798.355 1030.720 2028.605 ;
        RECT 754.520 1770.740 807.520 1798.355 ;
        RECT 754.520 1737.140 802.720 1770.740 ;
        RECT 806.720 1737.140 807.520 1770.740 ;
        RECT 754.520 1713.605 807.520 1737.140 ;
        RECT 811.520 1713.605 859.720 1798.355 ;
        RECT 863.720 1713.605 864.520 1798.355 ;
        RECT 868.520 1713.605 916.720 1798.355 ;
        RECT 920.720 1713.605 921.520 1798.355 ;
        RECT 925.520 1713.605 973.720 1798.355 ;
        RECT 977.720 1770.740 1030.720 1798.355 ;
        RECT 977.720 1737.140 978.520 1770.740 ;
        RECT 982.520 1737.140 1030.720 1770.740 ;
        RECT 977.720 1713.605 1030.720 1737.140 ;
        RECT 754.520 1483.355 1030.720 1713.605 ;
        RECT 754.520 1455.740 807.520 1483.355 ;
        RECT 754.520 1422.140 802.720 1455.740 ;
        RECT 806.720 1422.140 807.520 1455.740 ;
        RECT 754.520 1398.605 807.520 1422.140 ;
        RECT 811.520 1398.605 859.720 1483.355 ;
        RECT 863.720 1398.605 864.520 1483.355 ;
        RECT 868.520 1398.605 916.720 1483.355 ;
        RECT 920.720 1398.605 921.520 1483.355 ;
        RECT 925.520 1398.605 973.720 1483.355 ;
        RECT 977.720 1455.740 1030.720 1483.355 ;
        RECT 977.720 1422.140 978.520 1455.740 ;
        RECT 982.520 1422.140 1030.720 1455.740 ;
        RECT 977.720 1398.605 1030.720 1422.140 ;
        RECT 754.520 1168.355 1030.720 1398.605 ;
        RECT 754.520 1140.740 807.520 1168.355 ;
        RECT 754.520 1107.140 802.720 1140.740 ;
        RECT 806.720 1107.140 807.520 1140.740 ;
        RECT 754.520 1083.605 807.520 1107.140 ;
        RECT 811.520 1083.605 859.720 1168.355 ;
        RECT 863.720 1083.605 864.520 1168.355 ;
        RECT 868.520 1083.605 916.720 1168.355 ;
        RECT 920.720 1083.605 921.520 1168.355 ;
        RECT 925.520 1083.605 973.720 1168.355 ;
        RECT 977.720 1140.740 1030.720 1168.355 ;
        RECT 977.720 1107.140 978.520 1140.740 ;
        RECT 982.520 1107.140 1030.720 1140.740 ;
        RECT 977.720 1083.605 1030.720 1107.140 ;
        RECT 754.520 853.355 1030.720 1083.605 ;
        RECT 754.520 825.740 807.520 853.355 ;
        RECT 754.520 792.140 802.720 825.740 ;
        RECT 806.720 792.140 807.520 825.740 ;
        RECT 754.520 768.605 807.520 792.140 ;
        RECT 811.520 768.605 859.720 853.355 ;
        RECT 863.720 768.605 864.520 853.355 ;
        RECT 868.520 768.605 916.720 853.355 ;
        RECT 920.720 768.605 921.520 853.355 ;
        RECT 925.520 768.605 973.720 853.355 ;
        RECT 977.720 825.740 1030.720 853.355 ;
        RECT 977.720 792.140 978.520 825.740 ;
        RECT 982.520 792.140 1030.720 825.740 ;
        RECT 977.720 768.605 1030.720 792.140 ;
        RECT 754.520 538.355 1030.720 768.605 ;
        RECT 754.520 510.740 807.520 538.355 ;
        RECT 754.520 477.140 802.720 510.740 ;
        RECT 806.720 477.140 807.520 510.740 ;
        RECT 754.520 453.605 807.520 477.140 ;
        RECT 811.520 453.605 859.720 538.355 ;
        RECT 863.720 453.605 864.520 538.355 ;
        RECT 868.520 453.605 916.720 538.355 ;
        RECT 920.720 453.605 921.520 538.355 ;
        RECT 925.520 453.605 973.720 538.355 ;
        RECT 977.720 510.740 1030.720 538.355 ;
        RECT 977.720 477.140 978.520 510.740 ;
        RECT 982.520 477.140 1030.720 510.740 ;
        RECT 977.720 453.605 1030.720 477.140 ;
        RECT 754.520 223.355 1030.720 453.605 ;
        RECT 754.520 195.740 807.520 223.355 ;
        RECT 754.520 162.540 802.720 195.740 ;
        RECT 806.720 162.540 807.520 195.740 ;
        RECT 754.520 40.640 807.520 162.540 ;
        RECT 811.520 164.845 859.720 223.355 ;
        RECT 863.720 164.845 864.520 223.355 ;
        RECT 868.520 164.845 916.720 223.355 ;
        RECT 920.720 164.845 921.520 223.355 ;
        RECT 925.520 164.845 973.720 223.355 ;
        RECT 811.520 67.875 973.720 164.845 ;
        RECT 811.520 40.640 859.720 67.875 ;
        RECT 863.720 40.640 864.520 67.875 ;
        RECT 868.520 40.640 916.720 67.875 ;
        RECT 920.720 40.640 921.520 67.875 ;
        RECT 925.520 40.640 973.720 67.875 ;
        RECT 977.720 195.740 1030.720 223.355 ;
        RECT 977.720 162.540 978.520 195.740 ;
        RECT 982.520 162.540 1030.720 195.740 ;
        RECT 977.720 40.640 1030.720 162.540 ;
        RECT 1034.720 40.640 1035.520 2672.240 ;
        RECT 1039.520 2655.885 1092.520 2672.240 ;
        RECT 1096.520 2655.885 1144.720 2672.240 ;
        RECT 1148.720 2655.885 1149.520 2672.240 ;
        RECT 1153.520 2655.885 1201.720 2672.240 ;
        RECT 1205.720 2655.885 1206.520 2672.240 ;
        RECT 1210.520 2655.885 1258.720 2672.240 ;
        RECT 1262.720 2655.885 1315.720 2672.240 ;
        RECT 1039.520 2421.555 1315.720 2655.885 ;
        RECT 1039.520 2400.740 1092.520 2421.555 ;
        RECT 1039.520 2367.140 1087.720 2400.740 ;
        RECT 1091.720 2367.140 1092.520 2400.740 ;
        RECT 1039.520 2343.605 1092.520 2367.140 ;
        RECT 1096.520 2343.605 1144.720 2421.555 ;
        RECT 1148.720 2343.605 1149.520 2421.555 ;
        RECT 1153.520 2343.605 1201.720 2421.555 ;
        RECT 1205.720 2343.605 1206.520 2421.555 ;
        RECT 1210.520 2343.605 1258.720 2421.555 ;
        RECT 1262.720 2400.740 1315.720 2421.555 ;
        RECT 1262.720 2367.140 1263.520 2400.740 ;
        RECT 1267.520 2367.140 1315.720 2400.740 ;
        RECT 1262.720 2343.605 1315.720 2367.140 ;
        RECT 1039.520 2113.355 1315.720 2343.605 ;
        RECT 1039.520 2085.740 1092.520 2113.355 ;
        RECT 1039.520 2052.140 1087.720 2085.740 ;
        RECT 1091.720 2052.140 1092.520 2085.740 ;
        RECT 1039.520 2028.605 1092.520 2052.140 ;
        RECT 1096.520 2028.605 1144.720 2113.355 ;
        RECT 1148.720 2028.605 1149.520 2113.355 ;
        RECT 1153.520 2028.605 1201.720 2113.355 ;
        RECT 1205.720 2028.605 1206.520 2113.355 ;
        RECT 1210.520 2028.605 1258.720 2113.355 ;
        RECT 1262.720 2085.740 1315.720 2113.355 ;
        RECT 1262.720 2052.140 1263.520 2085.740 ;
        RECT 1267.520 2052.140 1315.720 2085.740 ;
        RECT 1262.720 2028.605 1315.720 2052.140 ;
        RECT 1039.520 1798.355 1315.720 2028.605 ;
        RECT 1039.520 1770.740 1092.520 1798.355 ;
        RECT 1039.520 1737.140 1087.720 1770.740 ;
        RECT 1091.720 1737.140 1092.520 1770.740 ;
        RECT 1039.520 1713.605 1092.520 1737.140 ;
        RECT 1096.520 1713.605 1144.720 1798.355 ;
        RECT 1148.720 1713.605 1149.520 1798.355 ;
        RECT 1153.520 1713.605 1201.720 1798.355 ;
        RECT 1205.720 1713.605 1206.520 1798.355 ;
        RECT 1210.520 1713.605 1258.720 1798.355 ;
        RECT 1262.720 1770.740 1315.720 1798.355 ;
        RECT 1262.720 1737.140 1263.520 1770.740 ;
        RECT 1267.520 1737.140 1315.720 1770.740 ;
        RECT 1262.720 1713.605 1315.720 1737.140 ;
        RECT 1039.520 1483.355 1315.720 1713.605 ;
        RECT 1039.520 1455.740 1092.520 1483.355 ;
        RECT 1039.520 1422.140 1087.720 1455.740 ;
        RECT 1091.720 1422.140 1092.520 1455.740 ;
        RECT 1039.520 1398.605 1092.520 1422.140 ;
        RECT 1096.520 1398.605 1144.720 1483.355 ;
        RECT 1148.720 1398.605 1149.520 1483.355 ;
        RECT 1153.520 1398.605 1201.720 1483.355 ;
        RECT 1205.720 1398.605 1206.520 1483.355 ;
        RECT 1210.520 1398.605 1258.720 1483.355 ;
        RECT 1262.720 1455.740 1315.720 1483.355 ;
        RECT 1262.720 1422.140 1263.520 1455.740 ;
        RECT 1267.520 1422.140 1315.720 1455.740 ;
        RECT 1262.720 1398.605 1315.720 1422.140 ;
        RECT 1039.520 1168.355 1315.720 1398.605 ;
        RECT 1039.520 1140.740 1092.520 1168.355 ;
        RECT 1039.520 1107.140 1087.720 1140.740 ;
        RECT 1091.720 1107.140 1092.520 1140.740 ;
        RECT 1039.520 1083.605 1092.520 1107.140 ;
        RECT 1096.520 1083.605 1144.720 1168.355 ;
        RECT 1148.720 1083.605 1149.520 1168.355 ;
        RECT 1153.520 1083.605 1201.720 1168.355 ;
        RECT 1205.720 1083.605 1206.520 1168.355 ;
        RECT 1210.520 1083.605 1258.720 1168.355 ;
        RECT 1262.720 1140.740 1315.720 1168.355 ;
        RECT 1262.720 1107.140 1263.520 1140.740 ;
        RECT 1267.520 1107.140 1315.720 1140.740 ;
        RECT 1262.720 1083.605 1315.720 1107.140 ;
        RECT 1039.520 853.355 1315.720 1083.605 ;
        RECT 1039.520 825.740 1092.520 853.355 ;
        RECT 1039.520 792.140 1087.720 825.740 ;
        RECT 1091.720 792.140 1092.520 825.740 ;
        RECT 1039.520 768.605 1092.520 792.140 ;
        RECT 1096.520 768.605 1144.720 853.355 ;
        RECT 1148.720 768.605 1149.520 853.355 ;
        RECT 1153.520 768.605 1201.720 853.355 ;
        RECT 1205.720 768.605 1206.520 853.355 ;
        RECT 1210.520 768.605 1258.720 853.355 ;
        RECT 1262.720 825.740 1315.720 853.355 ;
        RECT 1262.720 792.140 1263.520 825.740 ;
        RECT 1267.520 792.140 1315.720 825.740 ;
        RECT 1262.720 768.605 1315.720 792.140 ;
        RECT 1039.520 538.355 1315.720 768.605 ;
        RECT 1039.520 510.740 1092.520 538.355 ;
        RECT 1039.520 477.140 1087.720 510.740 ;
        RECT 1091.720 477.140 1092.520 510.740 ;
        RECT 1039.520 453.605 1092.520 477.140 ;
        RECT 1096.520 453.605 1144.720 538.355 ;
        RECT 1148.720 453.605 1149.520 538.355 ;
        RECT 1153.520 453.605 1201.720 538.355 ;
        RECT 1205.720 453.605 1206.520 538.355 ;
        RECT 1210.520 453.605 1258.720 538.355 ;
        RECT 1262.720 510.740 1315.720 538.355 ;
        RECT 1262.720 477.140 1263.520 510.740 ;
        RECT 1267.520 477.140 1315.720 510.740 ;
        RECT 1262.720 453.605 1315.720 477.140 ;
        RECT 1039.520 223.355 1315.720 453.605 ;
        RECT 1039.520 195.740 1092.520 223.355 ;
        RECT 1039.520 162.540 1087.720 195.740 ;
        RECT 1091.720 162.540 1092.520 195.740 ;
        RECT 1039.520 40.640 1092.520 162.540 ;
        RECT 1096.520 164.845 1144.720 223.355 ;
        RECT 1148.720 164.845 1149.520 223.355 ;
        RECT 1153.520 164.845 1201.720 223.355 ;
        RECT 1205.720 164.845 1206.520 223.355 ;
        RECT 1210.520 164.845 1258.720 223.355 ;
        RECT 1096.520 67.875 1258.720 164.845 ;
        RECT 1096.520 40.640 1144.720 67.875 ;
        RECT 1148.720 40.640 1149.520 67.875 ;
        RECT 1153.520 40.640 1201.720 67.875 ;
        RECT 1205.720 40.640 1206.520 67.875 ;
        RECT 1210.520 40.640 1258.720 67.875 ;
        RECT 1262.720 195.740 1315.720 223.355 ;
        RECT 1262.720 162.540 1263.520 195.740 ;
        RECT 1267.520 162.540 1315.720 195.740 ;
        RECT 1262.720 40.640 1315.720 162.540 ;
        RECT 1319.720 40.640 1320.520 2672.240 ;
        RECT 1324.520 2655.885 1377.520 2672.240 ;
        RECT 1381.520 2655.885 1429.720 2672.240 ;
        RECT 1433.720 2655.885 1434.520 2672.240 ;
        RECT 1438.520 2655.885 1486.720 2672.240 ;
        RECT 1490.720 2655.885 1491.520 2672.240 ;
        RECT 1495.520 2655.885 1543.720 2672.240 ;
        RECT 1547.720 2655.885 1600.720 2672.240 ;
        RECT 1324.520 2421.555 1600.720 2655.885 ;
        RECT 1324.520 2400.740 1377.520 2421.555 ;
        RECT 1324.520 2367.140 1372.720 2400.740 ;
        RECT 1376.720 2367.140 1377.520 2400.740 ;
        RECT 1324.520 2343.605 1377.520 2367.140 ;
        RECT 1381.520 2343.605 1429.720 2421.555 ;
        RECT 1433.720 2343.605 1434.520 2421.555 ;
        RECT 1438.520 2343.605 1486.720 2421.555 ;
        RECT 1490.720 2343.605 1491.520 2421.555 ;
        RECT 1495.520 2343.605 1543.720 2421.555 ;
        RECT 1547.720 2400.740 1600.720 2421.555 ;
        RECT 1547.720 2367.140 1548.520 2400.740 ;
        RECT 1552.520 2367.140 1600.720 2400.740 ;
        RECT 1547.720 2343.605 1600.720 2367.140 ;
        RECT 1324.520 2113.355 1600.720 2343.605 ;
        RECT 1324.520 2085.740 1377.520 2113.355 ;
        RECT 1324.520 2052.140 1372.720 2085.740 ;
        RECT 1376.720 2052.140 1377.520 2085.740 ;
        RECT 1324.520 2028.605 1377.520 2052.140 ;
        RECT 1381.520 2028.605 1429.720 2113.355 ;
        RECT 1433.720 2028.605 1434.520 2113.355 ;
        RECT 1438.520 2028.605 1486.720 2113.355 ;
        RECT 1490.720 2028.605 1491.520 2113.355 ;
        RECT 1495.520 2028.605 1543.720 2113.355 ;
        RECT 1547.720 2085.740 1600.720 2113.355 ;
        RECT 1547.720 2052.140 1548.520 2085.740 ;
        RECT 1552.520 2052.140 1600.720 2085.740 ;
        RECT 1547.720 2028.605 1600.720 2052.140 ;
        RECT 1324.520 1798.355 1600.720 2028.605 ;
        RECT 1324.520 1770.740 1377.520 1798.355 ;
        RECT 1324.520 1737.140 1372.720 1770.740 ;
        RECT 1376.720 1737.140 1377.520 1770.740 ;
        RECT 1324.520 1713.605 1377.520 1737.140 ;
        RECT 1381.520 1713.605 1429.720 1798.355 ;
        RECT 1433.720 1713.605 1434.520 1798.355 ;
        RECT 1438.520 1713.605 1486.720 1798.355 ;
        RECT 1490.720 1713.605 1491.520 1798.355 ;
        RECT 1495.520 1713.605 1543.720 1798.355 ;
        RECT 1547.720 1770.740 1600.720 1798.355 ;
        RECT 1547.720 1737.140 1548.520 1770.740 ;
        RECT 1552.520 1737.140 1600.720 1770.740 ;
        RECT 1547.720 1713.605 1600.720 1737.140 ;
        RECT 1324.520 1483.355 1600.720 1713.605 ;
        RECT 1324.520 1455.740 1377.520 1483.355 ;
        RECT 1324.520 1422.140 1372.720 1455.740 ;
        RECT 1376.720 1422.140 1377.520 1455.740 ;
        RECT 1324.520 1398.605 1377.520 1422.140 ;
        RECT 1381.520 1398.605 1429.720 1483.355 ;
        RECT 1433.720 1398.605 1434.520 1483.355 ;
        RECT 1438.520 1398.605 1486.720 1483.355 ;
        RECT 1490.720 1398.605 1491.520 1483.355 ;
        RECT 1495.520 1398.605 1543.720 1483.355 ;
        RECT 1547.720 1455.740 1600.720 1483.355 ;
        RECT 1547.720 1422.140 1548.520 1455.740 ;
        RECT 1552.520 1422.140 1600.720 1455.740 ;
        RECT 1547.720 1398.605 1600.720 1422.140 ;
        RECT 1324.520 1168.355 1600.720 1398.605 ;
        RECT 1324.520 1140.740 1377.520 1168.355 ;
        RECT 1324.520 1107.140 1372.720 1140.740 ;
        RECT 1376.720 1107.140 1377.520 1140.740 ;
        RECT 1324.520 1083.605 1377.520 1107.140 ;
        RECT 1381.520 1083.605 1429.720 1168.355 ;
        RECT 1433.720 1083.605 1434.520 1168.355 ;
        RECT 1438.520 1083.605 1486.720 1168.355 ;
        RECT 1490.720 1083.605 1491.520 1168.355 ;
        RECT 1495.520 1083.605 1543.720 1168.355 ;
        RECT 1547.720 1140.740 1600.720 1168.355 ;
        RECT 1547.720 1107.140 1548.520 1140.740 ;
        RECT 1552.520 1107.140 1600.720 1140.740 ;
        RECT 1547.720 1083.605 1600.720 1107.140 ;
        RECT 1324.520 853.355 1600.720 1083.605 ;
        RECT 1324.520 825.740 1377.520 853.355 ;
        RECT 1324.520 792.140 1372.720 825.740 ;
        RECT 1376.720 792.140 1377.520 825.740 ;
        RECT 1324.520 768.605 1377.520 792.140 ;
        RECT 1381.520 768.605 1429.720 853.355 ;
        RECT 1433.720 768.605 1434.520 853.355 ;
        RECT 1438.520 768.605 1486.720 853.355 ;
        RECT 1490.720 768.605 1491.520 853.355 ;
        RECT 1495.520 768.605 1543.720 853.355 ;
        RECT 1547.720 825.740 1600.720 853.355 ;
        RECT 1547.720 792.140 1548.520 825.740 ;
        RECT 1552.520 792.140 1600.720 825.740 ;
        RECT 1547.720 768.605 1600.720 792.140 ;
        RECT 1324.520 538.355 1600.720 768.605 ;
        RECT 1324.520 510.740 1377.520 538.355 ;
        RECT 1324.520 477.140 1372.720 510.740 ;
        RECT 1376.720 477.140 1377.520 510.740 ;
        RECT 1324.520 453.605 1377.520 477.140 ;
        RECT 1381.520 453.605 1429.720 538.355 ;
        RECT 1433.720 453.605 1434.520 538.355 ;
        RECT 1438.520 453.605 1486.720 538.355 ;
        RECT 1490.720 453.605 1491.520 538.355 ;
        RECT 1495.520 453.605 1543.720 538.355 ;
        RECT 1547.720 510.740 1600.720 538.355 ;
        RECT 1547.720 477.140 1548.520 510.740 ;
        RECT 1552.520 477.140 1600.720 510.740 ;
        RECT 1547.720 453.605 1600.720 477.140 ;
        RECT 1324.520 223.355 1600.720 453.605 ;
        RECT 1324.520 195.740 1377.520 223.355 ;
        RECT 1324.520 162.540 1372.720 195.740 ;
        RECT 1376.720 162.540 1377.520 195.740 ;
        RECT 1324.520 40.640 1377.520 162.540 ;
        RECT 1381.520 164.845 1429.720 223.355 ;
        RECT 1433.720 164.845 1434.520 223.355 ;
        RECT 1438.520 164.845 1486.720 223.355 ;
        RECT 1490.720 164.845 1491.520 223.355 ;
        RECT 1495.520 164.845 1543.720 223.355 ;
        RECT 1381.520 67.875 1543.720 164.845 ;
        RECT 1381.520 40.640 1429.720 67.875 ;
        RECT 1433.720 40.640 1434.520 67.875 ;
        RECT 1438.520 40.640 1486.720 67.875 ;
        RECT 1490.720 40.640 1491.520 67.875 ;
        RECT 1495.520 40.640 1543.720 67.875 ;
        RECT 1547.720 195.740 1600.720 223.355 ;
        RECT 1547.720 162.540 1548.520 195.740 ;
        RECT 1552.520 162.540 1600.720 195.740 ;
        RECT 1547.720 40.640 1600.720 162.540 ;
        RECT 1604.720 40.640 1605.520 2672.240 ;
        RECT 1609.520 2655.885 1662.520 2672.240 ;
        RECT 1666.520 2655.885 1714.720 2672.240 ;
        RECT 1718.720 2655.885 1719.520 2672.240 ;
        RECT 1723.520 2655.885 1771.720 2672.240 ;
        RECT 1775.720 2655.885 1776.520 2672.240 ;
        RECT 1780.520 2655.885 1828.720 2672.240 ;
        RECT 1832.720 2655.885 1885.720 2672.240 ;
        RECT 1609.520 2421.555 1885.720 2655.885 ;
        RECT 1609.520 2400.740 1662.520 2421.555 ;
        RECT 1609.520 2367.140 1657.720 2400.740 ;
        RECT 1661.720 2367.140 1662.520 2400.740 ;
        RECT 1609.520 2343.605 1662.520 2367.140 ;
        RECT 1666.520 2343.605 1714.720 2421.555 ;
        RECT 1718.720 2343.605 1719.520 2421.555 ;
        RECT 1723.520 2343.605 1771.720 2421.555 ;
        RECT 1775.720 2343.605 1776.520 2421.555 ;
        RECT 1780.520 2343.605 1828.720 2421.555 ;
        RECT 1832.720 2400.740 1885.720 2421.555 ;
        RECT 1832.720 2367.140 1833.520 2400.740 ;
        RECT 1837.520 2367.140 1885.720 2400.740 ;
        RECT 1832.720 2343.605 1885.720 2367.140 ;
        RECT 1609.520 2113.355 1885.720 2343.605 ;
        RECT 1609.520 2085.740 1662.520 2113.355 ;
        RECT 1609.520 2052.140 1657.720 2085.740 ;
        RECT 1661.720 2052.140 1662.520 2085.740 ;
        RECT 1609.520 2028.605 1662.520 2052.140 ;
        RECT 1666.520 2028.605 1714.720 2113.355 ;
        RECT 1718.720 2028.605 1719.520 2113.355 ;
        RECT 1723.520 2028.605 1771.720 2113.355 ;
        RECT 1775.720 2028.605 1776.520 2113.355 ;
        RECT 1780.520 2028.605 1828.720 2113.355 ;
        RECT 1832.720 2085.740 1885.720 2113.355 ;
        RECT 1832.720 2052.140 1833.520 2085.740 ;
        RECT 1837.520 2052.140 1885.720 2085.740 ;
        RECT 1832.720 2028.605 1885.720 2052.140 ;
        RECT 1609.520 1798.355 1885.720 2028.605 ;
        RECT 1609.520 1770.740 1662.520 1798.355 ;
        RECT 1609.520 1737.140 1657.720 1770.740 ;
        RECT 1661.720 1737.140 1662.520 1770.740 ;
        RECT 1609.520 1713.605 1662.520 1737.140 ;
        RECT 1666.520 1713.605 1714.720 1798.355 ;
        RECT 1718.720 1713.605 1719.520 1798.355 ;
        RECT 1723.520 1713.605 1771.720 1798.355 ;
        RECT 1775.720 1713.605 1776.520 1798.355 ;
        RECT 1780.520 1713.605 1828.720 1798.355 ;
        RECT 1832.720 1770.740 1885.720 1798.355 ;
        RECT 1832.720 1737.140 1833.520 1770.740 ;
        RECT 1837.520 1737.140 1885.720 1770.740 ;
        RECT 1832.720 1713.605 1885.720 1737.140 ;
        RECT 1609.520 1483.355 1885.720 1713.605 ;
        RECT 1609.520 1455.740 1662.520 1483.355 ;
        RECT 1609.520 1422.140 1657.720 1455.740 ;
        RECT 1661.720 1422.140 1662.520 1455.740 ;
        RECT 1609.520 1398.605 1662.520 1422.140 ;
        RECT 1666.520 1398.605 1714.720 1483.355 ;
        RECT 1718.720 1398.605 1719.520 1483.355 ;
        RECT 1723.520 1398.605 1771.720 1483.355 ;
        RECT 1775.720 1398.605 1776.520 1483.355 ;
        RECT 1780.520 1398.605 1828.720 1483.355 ;
        RECT 1832.720 1455.740 1885.720 1483.355 ;
        RECT 1832.720 1422.140 1833.520 1455.740 ;
        RECT 1837.520 1422.140 1885.720 1455.740 ;
        RECT 1832.720 1398.605 1885.720 1422.140 ;
        RECT 1609.520 1168.355 1885.720 1398.605 ;
        RECT 1609.520 1140.740 1662.520 1168.355 ;
        RECT 1609.520 1107.140 1657.720 1140.740 ;
        RECT 1661.720 1107.140 1662.520 1140.740 ;
        RECT 1609.520 1083.605 1662.520 1107.140 ;
        RECT 1666.520 1083.605 1714.720 1168.355 ;
        RECT 1718.720 1083.605 1719.520 1168.355 ;
        RECT 1723.520 1083.605 1771.720 1168.355 ;
        RECT 1775.720 1083.605 1776.520 1168.355 ;
        RECT 1780.520 1083.605 1828.720 1168.355 ;
        RECT 1832.720 1140.740 1885.720 1168.355 ;
        RECT 1832.720 1107.140 1833.520 1140.740 ;
        RECT 1837.520 1107.140 1885.720 1140.740 ;
        RECT 1832.720 1083.605 1885.720 1107.140 ;
        RECT 1609.520 853.355 1885.720 1083.605 ;
        RECT 1609.520 825.740 1662.520 853.355 ;
        RECT 1609.520 792.140 1657.720 825.740 ;
        RECT 1661.720 792.140 1662.520 825.740 ;
        RECT 1609.520 768.605 1662.520 792.140 ;
        RECT 1666.520 768.605 1714.720 853.355 ;
        RECT 1718.720 768.605 1719.520 853.355 ;
        RECT 1723.520 768.605 1771.720 853.355 ;
        RECT 1775.720 768.605 1776.520 853.355 ;
        RECT 1780.520 768.605 1828.720 853.355 ;
        RECT 1832.720 825.740 1885.720 853.355 ;
        RECT 1832.720 792.140 1833.520 825.740 ;
        RECT 1837.520 792.140 1885.720 825.740 ;
        RECT 1832.720 768.605 1885.720 792.140 ;
        RECT 1609.520 538.355 1885.720 768.605 ;
        RECT 1609.520 510.740 1662.520 538.355 ;
        RECT 1609.520 477.140 1657.720 510.740 ;
        RECT 1661.720 477.140 1662.520 510.740 ;
        RECT 1609.520 453.605 1662.520 477.140 ;
        RECT 1666.520 453.605 1714.720 538.355 ;
        RECT 1718.720 453.605 1719.520 538.355 ;
        RECT 1723.520 453.605 1771.720 538.355 ;
        RECT 1775.720 453.605 1776.520 538.355 ;
        RECT 1780.520 453.605 1828.720 538.355 ;
        RECT 1832.720 510.740 1885.720 538.355 ;
        RECT 1832.720 477.140 1833.520 510.740 ;
        RECT 1837.520 477.140 1885.720 510.740 ;
        RECT 1832.720 453.605 1885.720 477.140 ;
        RECT 1609.520 223.355 1885.720 453.605 ;
        RECT 1609.520 195.740 1662.520 223.355 ;
        RECT 1609.520 162.540 1657.720 195.740 ;
        RECT 1661.720 162.540 1662.520 195.740 ;
        RECT 1609.520 40.640 1662.520 162.540 ;
        RECT 1666.520 164.845 1714.720 223.355 ;
        RECT 1718.720 164.845 1719.520 223.355 ;
        RECT 1723.520 164.845 1771.720 223.355 ;
        RECT 1775.720 164.845 1776.520 223.355 ;
        RECT 1780.520 164.845 1828.720 223.355 ;
        RECT 1666.520 67.875 1828.720 164.845 ;
        RECT 1666.520 40.640 1714.720 67.875 ;
        RECT 1718.720 40.640 1719.520 67.875 ;
        RECT 1723.520 40.640 1771.720 67.875 ;
        RECT 1775.720 40.640 1776.520 67.875 ;
        RECT 1780.520 40.640 1828.720 67.875 ;
        RECT 1832.720 195.740 1885.720 223.355 ;
        RECT 1832.720 162.540 1833.520 195.740 ;
        RECT 1837.520 162.540 1885.720 195.740 ;
        RECT 1832.720 40.640 1885.720 162.540 ;
        RECT 1889.720 40.640 1890.520 2672.240 ;
        RECT 1894.520 2655.885 1947.520 2672.240 ;
        RECT 1951.520 2655.885 1999.720 2672.240 ;
        RECT 2003.720 2655.885 2004.520 2672.240 ;
        RECT 2008.520 2655.885 2056.720 2672.240 ;
        RECT 2060.720 2655.885 2061.520 2672.240 ;
        RECT 2065.520 2655.885 2113.720 2672.240 ;
        RECT 2117.720 2655.885 2170.720 2672.240 ;
        RECT 1894.520 2421.555 2170.720 2655.885 ;
        RECT 1894.520 2400.740 1947.520 2421.555 ;
        RECT 1894.520 2367.140 1942.720 2400.740 ;
        RECT 1946.720 2367.140 1947.520 2400.740 ;
        RECT 1894.520 2343.605 1947.520 2367.140 ;
        RECT 1951.520 2343.605 1999.720 2421.555 ;
        RECT 2003.720 2343.605 2004.520 2421.555 ;
        RECT 2008.520 2343.605 2056.720 2421.555 ;
        RECT 2060.720 2343.605 2061.520 2421.555 ;
        RECT 2065.520 2343.605 2113.720 2421.555 ;
        RECT 2117.720 2400.740 2170.720 2421.555 ;
        RECT 2117.720 2367.140 2118.520 2400.740 ;
        RECT 2122.520 2367.140 2170.720 2400.740 ;
        RECT 2117.720 2343.605 2170.720 2367.140 ;
        RECT 1894.520 2113.355 2170.720 2343.605 ;
        RECT 1894.520 2085.740 1947.520 2113.355 ;
        RECT 1894.520 2052.140 1942.720 2085.740 ;
        RECT 1946.720 2052.140 1947.520 2085.740 ;
        RECT 1894.520 2028.605 1947.520 2052.140 ;
        RECT 1951.520 2028.605 1999.720 2113.355 ;
        RECT 2003.720 2028.605 2004.520 2113.355 ;
        RECT 2008.520 2028.605 2056.720 2113.355 ;
        RECT 2060.720 2028.605 2061.520 2113.355 ;
        RECT 2065.520 2028.605 2113.720 2113.355 ;
        RECT 2117.720 2085.740 2170.720 2113.355 ;
        RECT 2117.720 2052.140 2118.520 2085.740 ;
        RECT 2122.520 2052.140 2170.720 2085.740 ;
        RECT 2117.720 2028.605 2170.720 2052.140 ;
        RECT 1894.520 1798.355 2170.720 2028.605 ;
        RECT 1894.520 1770.740 1947.520 1798.355 ;
        RECT 1894.520 1737.140 1942.720 1770.740 ;
        RECT 1946.720 1737.140 1947.520 1770.740 ;
        RECT 1894.520 1713.605 1947.520 1737.140 ;
        RECT 1951.520 1713.605 1999.720 1798.355 ;
        RECT 2003.720 1713.605 2004.520 1798.355 ;
        RECT 2008.520 1713.605 2056.720 1798.355 ;
        RECT 2060.720 1713.605 2061.520 1798.355 ;
        RECT 2065.520 1713.605 2113.720 1798.355 ;
        RECT 2117.720 1770.740 2170.720 1798.355 ;
        RECT 2117.720 1737.140 2118.520 1770.740 ;
        RECT 2122.520 1737.140 2170.720 1770.740 ;
        RECT 2117.720 1713.605 2170.720 1737.140 ;
        RECT 1894.520 1483.355 2170.720 1713.605 ;
        RECT 1894.520 1455.740 1947.520 1483.355 ;
        RECT 1894.520 1422.140 1942.720 1455.740 ;
        RECT 1946.720 1422.140 1947.520 1455.740 ;
        RECT 1894.520 1398.605 1947.520 1422.140 ;
        RECT 1951.520 1398.605 1999.720 1483.355 ;
        RECT 2003.720 1398.605 2004.520 1483.355 ;
        RECT 2008.520 1398.605 2056.720 1483.355 ;
        RECT 2060.720 1398.605 2061.520 1483.355 ;
        RECT 2065.520 1398.605 2113.720 1483.355 ;
        RECT 2117.720 1455.740 2170.720 1483.355 ;
        RECT 2117.720 1422.140 2118.520 1455.740 ;
        RECT 2122.520 1422.140 2170.720 1455.740 ;
        RECT 2117.720 1398.605 2170.720 1422.140 ;
        RECT 1894.520 1168.355 2170.720 1398.605 ;
        RECT 1894.520 1140.740 1947.520 1168.355 ;
        RECT 1894.520 1107.140 1942.720 1140.740 ;
        RECT 1946.720 1107.140 1947.520 1140.740 ;
        RECT 1894.520 1083.605 1947.520 1107.140 ;
        RECT 1951.520 1083.605 1999.720 1168.355 ;
        RECT 2003.720 1083.605 2004.520 1168.355 ;
        RECT 2008.520 1083.605 2056.720 1168.355 ;
        RECT 2060.720 1083.605 2061.520 1168.355 ;
        RECT 2065.520 1083.605 2113.720 1168.355 ;
        RECT 2117.720 1140.740 2170.720 1168.355 ;
        RECT 2117.720 1107.140 2118.520 1140.740 ;
        RECT 2122.520 1107.140 2170.720 1140.740 ;
        RECT 2117.720 1083.605 2170.720 1107.140 ;
        RECT 1894.520 853.355 2170.720 1083.605 ;
        RECT 1894.520 825.740 1947.520 853.355 ;
        RECT 1894.520 792.140 1942.720 825.740 ;
        RECT 1946.720 792.140 1947.520 825.740 ;
        RECT 1894.520 768.605 1947.520 792.140 ;
        RECT 1951.520 768.605 1999.720 853.355 ;
        RECT 2003.720 768.605 2004.520 853.355 ;
        RECT 2008.520 768.605 2056.720 853.355 ;
        RECT 2060.720 768.605 2061.520 853.355 ;
        RECT 2065.520 768.605 2113.720 853.355 ;
        RECT 2117.720 825.740 2170.720 853.355 ;
        RECT 2117.720 792.140 2118.520 825.740 ;
        RECT 2122.520 792.140 2170.720 825.740 ;
        RECT 2117.720 768.605 2170.720 792.140 ;
        RECT 1894.520 538.355 2170.720 768.605 ;
        RECT 1894.520 510.740 1947.520 538.355 ;
        RECT 1894.520 477.140 1942.720 510.740 ;
        RECT 1946.720 477.140 1947.520 510.740 ;
        RECT 1894.520 453.605 1947.520 477.140 ;
        RECT 1951.520 453.605 1999.720 538.355 ;
        RECT 2003.720 453.605 2004.520 538.355 ;
        RECT 2008.520 453.605 2056.720 538.355 ;
        RECT 2060.720 453.605 2061.520 538.355 ;
        RECT 2065.520 453.605 2113.720 538.355 ;
        RECT 2117.720 510.740 2170.720 538.355 ;
        RECT 2117.720 477.140 2118.520 510.740 ;
        RECT 2122.520 477.140 2170.720 510.740 ;
        RECT 2117.720 453.605 2170.720 477.140 ;
        RECT 1894.520 223.355 2170.720 453.605 ;
        RECT 1894.520 195.740 1947.520 223.355 ;
        RECT 1894.520 162.540 1942.720 195.740 ;
        RECT 1946.720 162.540 1947.520 195.740 ;
        RECT 1894.520 40.640 1947.520 162.540 ;
        RECT 1951.520 164.845 1999.720 223.355 ;
        RECT 2003.720 164.845 2004.520 223.355 ;
        RECT 2008.520 164.845 2056.720 223.355 ;
        RECT 2060.720 164.845 2061.520 223.355 ;
        RECT 2065.520 164.845 2113.720 223.355 ;
        RECT 1951.520 67.875 2113.720 164.845 ;
        RECT 1951.520 40.640 1999.720 67.875 ;
        RECT 2003.720 40.640 2004.520 67.875 ;
        RECT 2008.520 40.640 2056.720 67.875 ;
        RECT 2060.720 40.640 2061.520 67.875 ;
        RECT 2065.520 40.640 2113.720 67.875 ;
        RECT 2117.720 195.740 2170.720 223.355 ;
        RECT 2117.720 162.540 2118.520 195.740 ;
        RECT 2122.520 162.540 2170.720 195.740 ;
        RECT 2117.720 40.640 2170.720 162.540 ;
        RECT 2174.720 40.640 2175.520 2672.240 ;
        RECT 2179.520 2407.275 2431.320 2672.240 ;
        RECT 2179.520 2400.740 2232.520 2407.275 ;
        RECT 2179.520 2367.140 2227.720 2400.740 ;
        RECT 2231.720 2367.140 2232.520 2400.740 ;
        RECT 2179.520 2364.685 2232.520 2367.140 ;
        RECT 2236.520 2364.685 2284.720 2407.275 ;
        RECT 2288.720 2364.685 2289.520 2407.275 ;
        RECT 2293.520 2364.685 2341.720 2407.275 ;
        RECT 2345.720 2364.685 2346.520 2407.275 ;
        RECT 2350.520 2364.685 2398.720 2407.275 ;
        RECT 2402.720 2400.740 2431.320 2407.275 ;
        RECT 2402.720 2367.140 2403.520 2400.740 ;
        RECT 2407.520 2367.140 2431.320 2400.740 ;
        RECT 2402.720 2364.685 2431.320 2367.140 ;
        RECT 2179.520 2086.835 2431.320 2364.685 ;
        RECT 2179.520 2085.740 2232.520 2086.835 ;
        RECT 2179.520 2052.140 2227.720 2085.740 ;
        RECT 2231.720 2052.140 2232.520 2085.740 ;
        RECT 2179.520 2049.685 2232.520 2052.140 ;
        RECT 2236.520 2049.685 2284.720 2086.835 ;
        RECT 2288.720 2049.685 2289.520 2086.835 ;
        RECT 2293.520 2049.685 2341.720 2086.835 ;
        RECT 2345.720 2049.685 2346.520 2086.835 ;
        RECT 2350.520 2049.685 2398.720 2086.835 ;
        RECT 2402.720 2085.740 2431.320 2086.835 ;
        RECT 2402.720 2052.140 2403.520 2085.740 ;
        RECT 2407.520 2052.140 2431.320 2085.740 ;
        RECT 2402.720 2049.685 2431.320 2052.140 ;
        RECT 2179.520 1771.835 2431.320 2049.685 ;
        RECT 2179.520 1770.740 2232.520 1771.835 ;
        RECT 2179.520 1737.140 2227.720 1770.740 ;
        RECT 2231.720 1737.140 2232.520 1770.740 ;
        RECT 2179.520 1734.685 2232.520 1737.140 ;
        RECT 2236.520 1734.685 2284.720 1771.835 ;
        RECT 2288.720 1734.685 2289.520 1771.835 ;
        RECT 2293.520 1734.685 2341.720 1771.835 ;
        RECT 2345.720 1734.685 2346.520 1771.835 ;
        RECT 2350.520 1734.685 2398.720 1771.835 ;
        RECT 2402.720 1770.740 2431.320 1771.835 ;
        RECT 2402.720 1737.140 2403.520 1770.740 ;
        RECT 2407.520 1737.140 2431.320 1770.740 ;
        RECT 2402.720 1734.685 2431.320 1737.140 ;
        RECT 2179.520 1456.835 2431.320 1734.685 ;
        RECT 2179.520 1455.740 2232.520 1456.835 ;
        RECT 2179.520 1422.140 2227.720 1455.740 ;
        RECT 2231.720 1422.140 2232.520 1455.740 ;
        RECT 2179.520 1419.685 2232.520 1422.140 ;
        RECT 2236.520 1419.685 2284.720 1456.835 ;
        RECT 2288.720 1419.685 2289.520 1456.835 ;
        RECT 2293.520 1419.685 2341.720 1456.835 ;
        RECT 2345.720 1419.685 2346.520 1456.835 ;
        RECT 2350.520 1419.685 2398.720 1456.835 ;
        RECT 2402.720 1455.740 2431.320 1456.835 ;
        RECT 2402.720 1422.140 2403.520 1455.740 ;
        RECT 2407.520 1422.140 2431.320 1455.740 ;
        RECT 2402.720 1419.685 2431.320 1422.140 ;
        RECT 2179.520 1141.835 2431.320 1419.685 ;
        RECT 2179.520 1140.740 2232.520 1141.835 ;
        RECT 2179.520 1107.140 2227.720 1140.740 ;
        RECT 2231.720 1107.140 2232.520 1140.740 ;
        RECT 2179.520 1104.685 2232.520 1107.140 ;
        RECT 2236.520 1104.685 2284.720 1141.835 ;
        RECT 2288.720 1104.685 2289.520 1141.835 ;
        RECT 2293.520 1104.685 2341.720 1141.835 ;
        RECT 2345.720 1104.685 2346.520 1141.835 ;
        RECT 2350.520 1104.685 2398.720 1141.835 ;
        RECT 2402.720 1140.740 2431.320 1141.835 ;
        RECT 2402.720 1107.140 2403.520 1140.740 ;
        RECT 2407.520 1107.140 2431.320 1140.740 ;
        RECT 2402.720 1104.685 2431.320 1107.140 ;
        RECT 2179.520 826.835 2431.320 1104.685 ;
        RECT 2179.520 825.740 2232.520 826.835 ;
        RECT 2179.520 792.140 2227.720 825.740 ;
        RECT 2231.720 792.140 2232.520 825.740 ;
        RECT 2179.520 789.685 2232.520 792.140 ;
        RECT 2236.520 789.685 2284.720 826.835 ;
        RECT 2288.720 789.685 2289.520 826.835 ;
        RECT 2293.520 789.685 2341.720 826.835 ;
        RECT 2345.720 789.685 2346.520 826.835 ;
        RECT 2350.520 789.685 2398.720 826.835 ;
        RECT 2402.720 825.740 2431.320 826.835 ;
        RECT 2402.720 792.140 2403.520 825.740 ;
        RECT 2407.520 792.140 2431.320 825.740 ;
        RECT 2402.720 789.685 2431.320 792.140 ;
        RECT 2179.520 511.835 2431.320 789.685 ;
        RECT 2179.520 510.740 2232.520 511.835 ;
        RECT 2179.520 477.140 2227.720 510.740 ;
        RECT 2231.720 477.140 2232.520 510.740 ;
        RECT 2179.520 474.685 2232.520 477.140 ;
        RECT 2236.520 474.685 2284.720 511.835 ;
        RECT 2288.720 474.685 2289.520 511.835 ;
        RECT 2293.520 474.685 2341.720 511.835 ;
        RECT 2345.720 474.685 2346.520 511.835 ;
        RECT 2350.520 474.685 2398.720 511.835 ;
        RECT 2402.720 510.740 2431.320 511.835 ;
        RECT 2402.720 477.140 2403.520 510.740 ;
        RECT 2407.520 477.140 2431.320 510.740 ;
        RECT 2402.720 474.685 2431.320 477.140 ;
        RECT 2179.520 196.835 2431.320 474.685 ;
        RECT 2179.520 195.740 2232.520 196.835 ;
        RECT 2179.520 162.540 2227.720 195.740 ;
        RECT 2231.720 162.540 2232.520 195.740 ;
        RECT 2179.520 160.765 2232.520 162.540 ;
        RECT 2236.520 160.765 2284.720 196.835 ;
        RECT 2288.720 160.765 2289.520 196.835 ;
        RECT 2293.520 160.765 2341.720 196.835 ;
        RECT 2179.520 61.075 2341.720 160.765 ;
        RECT 2179.520 40.640 2232.520 61.075 ;
        RECT 2236.520 40.640 2284.720 61.075 ;
        RECT 2288.720 40.640 2289.520 61.075 ;
        RECT 2293.520 40.640 2341.720 61.075 ;
        RECT 2345.720 40.640 2346.520 196.835 ;
        RECT 2350.520 40.640 2398.720 196.835 ;
        RECT 2402.720 195.740 2431.320 196.835 ;
        RECT 2402.720 162.540 2403.520 195.740 ;
        RECT 2407.520 162.540 2431.320 195.740 ;
        RECT 2402.720 40.640 2431.320 162.540 ;
  END
END fpga_core
END LIBRARY

