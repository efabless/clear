magic
tech sky130A
magscale 1 2
timestamp 1679319064
<< obsli1 >>
rect 1104 2159 49864 54417
<< obsm1 >>
rect 934 1980 49864 54528
<< metal2 >>
rect 3330 56200 3386 57000
rect 3882 56200 3938 57000
rect 4434 56200 4490 57000
rect 4986 56200 5042 57000
rect 5538 56200 5594 57000
rect 6090 56200 6146 57000
rect 6642 56200 6698 57000
rect 7194 56200 7250 57000
rect 7746 56200 7802 57000
rect 8298 56200 8354 57000
rect 8850 56200 8906 57000
rect 9402 56200 9458 57000
rect 9954 56200 10010 57000
rect 10506 56200 10562 57000
rect 11058 56200 11114 57000
rect 11610 56200 11666 57000
rect 12162 56200 12218 57000
rect 12714 56200 12770 57000
rect 13266 56200 13322 57000
rect 13818 56200 13874 57000
rect 14370 56200 14426 57000
rect 14922 56200 14978 57000
rect 15474 56200 15530 57000
rect 16026 56200 16082 57000
rect 16578 56200 16634 57000
rect 17130 56200 17186 57000
rect 17682 56200 17738 57000
rect 18234 56200 18290 57000
rect 18786 56200 18842 57000
rect 19338 56200 19394 57000
rect 19890 56200 19946 57000
rect 20442 56200 20498 57000
rect 20994 56200 21050 57000
rect 21546 56200 21602 57000
rect 22098 56200 22154 57000
rect 22650 56200 22706 57000
rect 23202 56200 23258 57000
rect 23754 56200 23810 57000
rect 24306 56200 24362 57000
rect 24858 56200 24914 57000
rect 25410 56200 25466 57000
rect 25962 56200 26018 57000
rect 26514 56200 26570 57000
rect 27066 56200 27122 57000
rect 27618 56200 27674 57000
rect 28170 56200 28226 57000
rect 28722 56200 28778 57000
rect 29274 56200 29330 57000
rect 29826 56200 29882 57000
rect 30378 56200 30434 57000
rect 30930 56200 30986 57000
rect 31482 56200 31538 57000
rect 32034 56200 32090 57000
rect 32586 56200 32642 57000
rect 33138 56200 33194 57000
rect 33690 56200 33746 57000
rect 34242 56200 34298 57000
rect 34794 56200 34850 57000
rect 35346 56200 35402 57000
rect 35898 56200 35954 57000
rect 36450 56200 36506 57000
rect 38106 56200 38162 57000
rect 38658 56200 38714 57000
rect 39210 56200 39266 57000
rect 39762 56200 39818 57000
rect 40314 56200 40370 57000
rect 40866 56200 40922 57000
rect 41418 56200 41474 57000
rect 41970 56200 42026 57000
rect 42522 56200 42578 57000
rect 43074 56200 43130 57000
rect 43626 56200 43682 57000
rect 44178 56200 44234 57000
rect 44730 56200 44786 57000
rect 45282 56200 45338 57000
rect 45834 56200 45890 57000
rect 46386 56200 46442 57000
rect 46938 56200 46994 57000
rect 47490 56200 47546 57000
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4434 0 4490 800
rect 4986 0 5042 800
rect 5538 0 5594 800
rect 6090 0 6146 800
rect 6642 0 6698 800
rect 7194 0 7250 800
rect 7746 0 7802 800
rect 8298 0 8354 800
rect 8850 0 8906 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10506 0 10562 800
rect 11058 0 11114 800
rect 11610 0 11666 800
rect 12162 0 12218 800
rect 12714 0 12770 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19890 0 19946 800
rect 20442 0 20498 800
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
rect 23202 0 23258 800
rect 23754 0 23810 800
rect 24306 0 24362 800
rect 24858 0 24914 800
rect 25410 0 25466 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 27066 0 27122 800
rect 27618 0 27674 800
rect 28170 0 28226 800
rect 28722 0 28778 800
rect 29274 0 29330 800
rect 29826 0 29882 800
rect 30378 0 30434 800
rect 30930 0 30986 800
rect 31482 0 31538 800
rect 32034 0 32090 800
rect 32586 0 32642 800
rect 33138 0 33194 800
rect 33690 0 33746 800
rect 34242 0 34298 800
rect 34794 0 34850 800
rect 35346 0 35402 800
rect 35898 0 35954 800
rect 36450 0 36506 800
rect 37002 0 37058 800
rect 37554 0 37610 800
rect 38106 0 38162 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39762 0 39818 800
rect 40314 0 40370 800
rect 40866 0 40922 800
rect 41418 0 41474 800
rect 41970 0 42026 800
rect 42522 0 42578 800
rect 43074 0 43130 800
rect 43626 0 43682 800
rect 44178 0 44234 800
rect 44730 0 44786 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46386 0 46442 800
rect 46938 0 46994 800
<< obsm2 >>
rect 938 56144 3274 56250
rect 3442 56144 3826 56250
rect 3994 56144 4378 56250
rect 4546 56144 4930 56250
rect 5098 56144 5482 56250
rect 5650 56144 6034 56250
rect 6202 56144 6586 56250
rect 6754 56144 7138 56250
rect 7306 56144 7690 56250
rect 7858 56144 8242 56250
rect 8410 56144 8794 56250
rect 8962 56144 9346 56250
rect 9514 56144 9898 56250
rect 10066 56144 10450 56250
rect 10618 56144 11002 56250
rect 11170 56144 11554 56250
rect 11722 56144 12106 56250
rect 12274 56144 12658 56250
rect 12826 56144 13210 56250
rect 13378 56144 13762 56250
rect 13930 56144 14314 56250
rect 14482 56144 14866 56250
rect 15034 56144 15418 56250
rect 15586 56144 15970 56250
rect 16138 56144 16522 56250
rect 16690 56144 17074 56250
rect 17242 56144 17626 56250
rect 17794 56144 18178 56250
rect 18346 56144 18730 56250
rect 18898 56144 19282 56250
rect 19450 56144 19834 56250
rect 20002 56144 20386 56250
rect 20554 56144 20938 56250
rect 21106 56144 21490 56250
rect 21658 56144 22042 56250
rect 22210 56144 22594 56250
rect 22762 56144 23146 56250
rect 23314 56144 23698 56250
rect 23866 56144 24250 56250
rect 24418 56144 24802 56250
rect 24970 56144 25354 56250
rect 25522 56144 25906 56250
rect 26074 56144 26458 56250
rect 26626 56144 27010 56250
rect 27178 56144 27562 56250
rect 27730 56144 28114 56250
rect 28282 56144 28666 56250
rect 28834 56144 29218 56250
rect 29386 56144 29770 56250
rect 29938 56144 30322 56250
rect 30490 56144 30874 56250
rect 31042 56144 31426 56250
rect 31594 56144 31978 56250
rect 32146 56144 32530 56250
rect 32698 56144 33082 56250
rect 33250 56144 33634 56250
rect 33802 56144 34186 56250
rect 34354 56144 34738 56250
rect 34906 56144 35290 56250
rect 35458 56144 35842 56250
rect 36010 56144 36394 56250
rect 36562 56144 38050 56250
rect 38218 56144 38602 56250
rect 38770 56144 39154 56250
rect 39322 56144 39706 56250
rect 39874 56144 40258 56250
rect 40426 56144 40810 56250
rect 40978 56144 41362 56250
rect 41530 56144 41914 56250
rect 42082 56144 42466 56250
rect 42634 56144 43018 56250
rect 43186 56144 43570 56250
rect 43738 56144 44122 56250
rect 44290 56144 44674 56250
rect 44842 56144 45226 56250
rect 45394 56144 45778 56250
rect 45946 56144 46330 56250
rect 46498 56144 46882 56250
rect 47050 56144 47434 56250
rect 47602 56144 49386 56250
rect 938 856 49386 56144
rect 938 734 3274 856
rect 3442 734 3826 856
rect 3994 734 4378 856
rect 4546 734 4930 856
rect 5098 734 5482 856
rect 5650 734 6034 856
rect 6202 734 6586 856
rect 6754 734 7138 856
rect 7306 734 7690 856
rect 7858 734 8242 856
rect 8410 734 8794 856
rect 8962 734 9346 856
rect 9514 734 9898 856
rect 10066 734 10450 856
rect 10618 734 11002 856
rect 11170 734 11554 856
rect 11722 734 12106 856
rect 12274 734 12658 856
rect 12826 734 13210 856
rect 13378 734 13762 856
rect 13930 734 14314 856
rect 14482 734 14866 856
rect 15034 734 15418 856
rect 15586 734 15970 856
rect 16138 734 16522 856
rect 16690 734 17074 856
rect 17242 734 17626 856
rect 17794 734 18178 856
rect 18346 734 18730 856
rect 18898 734 19282 856
rect 19450 734 19834 856
rect 20002 734 20386 856
rect 20554 734 20938 856
rect 21106 734 21490 856
rect 21658 734 22042 856
rect 22210 734 22594 856
rect 22762 734 23146 856
rect 23314 734 23698 856
rect 23866 734 24250 856
rect 24418 734 24802 856
rect 24970 734 25354 856
rect 25522 734 25906 856
rect 26074 734 26458 856
rect 26626 734 27010 856
rect 27178 734 27562 856
rect 27730 734 28114 856
rect 28282 734 28666 856
rect 28834 734 29218 856
rect 29386 734 29770 856
rect 29938 734 30322 856
rect 30490 734 30874 856
rect 31042 734 31426 856
rect 31594 734 31978 856
rect 32146 734 32530 856
rect 32698 734 33082 856
rect 33250 734 33634 856
rect 33802 734 34186 856
rect 34354 734 34738 856
rect 34906 734 35290 856
rect 35458 734 35842 856
rect 36010 734 36394 856
rect 36562 734 36946 856
rect 37114 734 37498 856
rect 37666 734 38050 856
rect 38218 734 38602 856
rect 38770 734 39154 856
rect 39322 734 39706 856
rect 39874 734 40258 856
rect 40426 734 40810 856
rect 40978 734 41362 856
rect 41530 734 41914 856
rect 42082 734 42466 856
rect 42634 734 43018 856
rect 43186 734 43570 856
rect 43738 734 44122 856
rect 44290 734 44674 856
rect 44842 734 45226 856
rect 45394 734 45778 856
rect 45946 734 46330 856
rect 46498 734 46882 856
rect 47050 734 49386 856
<< metal3 >>
rect 50200 55632 51000 55752
rect 50200 53456 51000 53576
rect 0 52504 800 52624
rect 0 51824 800 51944
rect 0 51144 800 51264
rect 50200 51280 51000 51400
rect 0 50464 800 50584
rect 0 49784 800 49904
rect 0 49104 800 49224
rect 50200 49104 51000 49224
rect 0 48424 800 48544
rect 0 47744 800 47864
rect 0 47064 800 47184
rect 50200 46928 51000 47048
rect 0 46384 800 46504
rect 0 45704 800 45824
rect 0 45024 800 45144
rect 50200 44752 51000 44872
rect 0 44344 800 44464
rect 0 43664 800 43784
rect 0 42984 800 43104
rect 50200 42576 51000 42696
rect 0 42304 800 42424
rect 0 41624 800 41744
rect 0 40944 800 41064
rect 0 40264 800 40384
rect 50200 40400 51000 40520
rect 0 39584 800 39704
rect 0 38904 800 39024
rect 0 38224 800 38344
rect 50200 38224 51000 38344
rect 0 37544 800 37664
rect 0 36864 800 36984
rect 0 36184 800 36304
rect 50200 36048 51000 36168
rect 0 35504 800 35624
rect 0 34824 800 34944
rect 0 34144 800 34264
rect 50200 33872 51000 33992
rect 0 33464 800 33584
rect 0 32784 800 32904
rect 0 32104 800 32224
rect 50200 31696 51000 31816
rect 0 31424 800 31544
rect 0 30744 800 30864
rect 0 30064 800 30184
rect 0 29384 800 29504
rect 50200 29520 51000 29640
rect 0 28704 800 28824
rect 0 28024 800 28144
rect 0 27344 800 27464
rect 50200 27344 51000 27464
rect 0 26664 800 26784
rect 0 25984 800 26104
rect 0 25304 800 25424
rect 50200 25168 51000 25288
rect 0 24624 800 24744
rect 0 23944 800 24064
rect 0 23264 800 23384
rect 50200 22992 51000 23112
rect 0 22584 800 22704
rect 0 21904 800 22024
rect 0 21224 800 21344
rect 50200 20816 51000 20936
rect 0 20544 800 20664
rect 0 19864 800 19984
rect 0 19184 800 19304
rect 0 18504 800 18624
rect 50200 18640 51000 18760
rect 0 17824 800 17944
rect 0 17144 800 17264
rect 0 16464 800 16584
rect 50200 16464 51000 16584
rect 0 15784 800 15904
rect 0 15104 800 15224
rect 0 14424 800 14544
rect 50200 14288 51000 14408
rect 0 13744 800 13864
rect 0 13064 800 13184
rect 0 12384 800 12504
rect 50200 12112 51000 12232
rect 0 11704 800 11824
rect 0 11024 800 11144
rect 0 10344 800 10464
rect 50200 9936 51000 10056
rect 0 9664 800 9784
rect 0 8984 800 9104
rect 0 8304 800 8424
rect 0 7624 800 7744
rect 50200 7760 51000 7880
rect 0 6944 800 7064
rect 0 6264 800 6384
rect 0 5584 800 5704
rect 50200 5584 51000 5704
rect 0 4904 800 5024
rect 50200 3408 51000 3528
rect 50200 1232 51000 1352
<< obsm3 >>
rect 800 55552 50120 55725
rect 800 53656 50200 55552
rect 800 53376 50120 53656
rect 800 52704 50200 53376
rect 880 52424 50200 52704
rect 800 52024 50200 52424
rect 880 51744 50200 52024
rect 800 51480 50200 51744
rect 800 51344 50120 51480
rect 880 51200 50120 51344
rect 880 51064 50200 51200
rect 800 50664 50200 51064
rect 880 50384 50200 50664
rect 800 49984 50200 50384
rect 880 49704 50200 49984
rect 800 49304 50200 49704
rect 880 49024 50120 49304
rect 800 48624 50200 49024
rect 880 48344 50200 48624
rect 800 47944 50200 48344
rect 880 47664 50200 47944
rect 800 47264 50200 47664
rect 880 47128 50200 47264
rect 880 46984 50120 47128
rect 800 46848 50120 46984
rect 800 46584 50200 46848
rect 880 46304 50200 46584
rect 800 45904 50200 46304
rect 880 45624 50200 45904
rect 800 45224 50200 45624
rect 880 44952 50200 45224
rect 880 44944 50120 44952
rect 800 44672 50120 44944
rect 800 44544 50200 44672
rect 880 44264 50200 44544
rect 800 43864 50200 44264
rect 880 43584 50200 43864
rect 800 43184 50200 43584
rect 880 42904 50200 43184
rect 800 42776 50200 42904
rect 800 42504 50120 42776
rect 880 42496 50120 42504
rect 880 42224 50200 42496
rect 800 41824 50200 42224
rect 880 41544 50200 41824
rect 800 41144 50200 41544
rect 880 40864 50200 41144
rect 800 40600 50200 40864
rect 800 40464 50120 40600
rect 880 40320 50120 40464
rect 880 40184 50200 40320
rect 800 39784 50200 40184
rect 880 39504 50200 39784
rect 800 39104 50200 39504
rect 880 38824 50200 39104
rect 800 38424 50200 38824
rect 880 38144 50120 38424
rect 800 37744 50200 38144
rect 880 37464 50200 37744
rect 800 37064 50200 37464
rect 880 36784 50200 37064
rect 800 36384 50200 36784
rect 880 36248 50200 36384
rect 880 36104 50120 36248
rect 800 35968 50120 36104
rect 800 35704 50200 35968
rect 880 35424 50200 35704
rect 800 35024 50200 35424
rect 880 34744 50200 35024
rect 800 34344 50200 34744
rect 880 34072 50200 34344
rect 880 34064 50120 34072
rect 800 33792 50120 34064
rect 800 33664 50200 33792
rect 880 33384 50200 33664
rect 800 32984 50200 33384
rect 880 32704 50200 32984
rect 800 32304 50200 32704
rect 880 32024 50200 32304
rect 800 31896 50200 32024
rect 800 31624 50120 31896
rect 880 31616 50120 31624
rect 880 31344 50200 31616
rect 800 30944 50200 31344
rect 880 30664 50200 30944
rect 800 30264 50200 30664
rect 880 29984 50200 30264
rect 800 29720 50200 29984
rect 800 29584 50120 29720
rect 880 29440 50120 29584
rect 880 29304 50200 29440
rect 800 28904 50200 29304
rect 880 28624 50200 28904
rect 800 28224 50200 28624
rect 880 27944 50200 28224
rect 800 27544 50200 27944
rect 880 27264 50120 27544
rect 800 26864 50200 27264
rect 880 26584 50200 26864
rect 800 26184 50200 26584
rect 880 25904 50200 26184
rect 800 25504 50200 25904
rect 880 25368 50200 25504
rect 880 25224 50120 25368
rect 800 25088 50120 25224
rect 800 24824 50200 25088
rect 880 24544 50200 24824
rect 800 24144 50200 24544
rect 880 23864 50200 24144
rect 800 23464 50200 23864
rect 880 23192 50200 23464
rect 880 23184 50120 23192
rect 800 22912 50120 23184
rect 800 22784 50200 22912
rect 880 22504 50200 22784
rect 800 22104 50200 22504
rect 880 21824 50200 22104
rect 800 21424 50200 21824
rect 880 21144 50200 21424
rect 800 21016 50200 21144
rect 800 20744 50120 21016
rect 880 20736 50120 20744
rect 880 20464 50200 20736
rect 800 20064 50200 20464
rect 880 19784 50200 20064
rect 800 19384 50200 19784
rect 880 19104 50200 19384
rect 800 18840 50200 19104
rect 800 18704 50120 18840
rect 880 18560 50120 18704
rect 880 18424 50200 18560
rect 800 18024 50200 18424
rect 880 17744 50200 18024
rect 800 17344 50200 17744
rect 880 17064 50200 17344
rect 800 16664 50200 17064
rect 880 16384 50120 16664
rect 800 15984 50200 16384
rect 880 15704 50200 15984
rect 800 15304 50200 15704
rect 880 15024 50200 15304
rect 800 14624 50200 15024
rect 880 14488 50200 14624
rect 880 14344 50120 14488
rect 800 14208 50120 14344
rect 800 13944 50200 14208
rect 880 13664 50200 13944
rect 800 13264 50200 13664
rect 880 12984 50200 13264
rect 800 12584 50200 12984
rect 880 12312 50200 12584
rect 880 12304 50120 12312
rect 800 12032 50120 12304
rect 800 11904 50200 12032
rect 880 11624 50200 11904
rect 800 11224 50200 11624
rect 880 10944 50200 11224
rect 800 10544 50200 10944
rect 880 10264 50200 10544
rect 800 10136 50200 10264
rect 800 9864 50120 10136
rect 880 9856 50120 9864
rect 880 9584 50200 9856
rect 800 9184 50200 9584
rect 880 8904 50200 9184
rect 800 8504 50200 8904
rect 880 8224 50200 8504
rect 800 7960 50200 8224
rect 800 7824 50120 7960
rect 880 7680 50120 7824
rect 880 7544 50200 7680
rect 800 7144 50200 7544
rect 880 6864 50200 7144
rect 800 6464 50200 6864
rect 880 6184 50200 6464
rect 800 5784 50200 6184
rect 880 5504 50120 5784
rect 800 5104 50200 5504
rect 880 4824 50200 5104
rect 800 3608 50200 4824
rect 800 3328 50120 3608
rect 800 1432 50200 3328
rect 800 1259 50120 1432
<< metal4 >>
rect 2944 2128 3264 54448
rect 7944 2128 8264 54448
rect 12944 2128 13264 54448
rect 17944 2128 18264 54448
rect 22944 2128 23264 54448
rect 27944 2128 28264 54448
rect 32944 2128 33264 54448
rect 37944 2128 38264 54448
rect 42944 2128 43264 54448
rect 47944 2128 48264 54448
<< obsm4 >>
rect 3371 2347 7864 53957
rect 8344 2347 12864 53957
rect 13344 2347 17864 53957
rect 18344 2347 22864 53957
rect 23344 2347 27864 53957
rect 28344 2347 32864 53957
rect 33344 2347 37864 53957
rect 38344 2347 42864 53957
rect 43344 2347 46861 53957
<< labels >>
rlabel metal4 s 7944 2128 8264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27944 2128 28264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37944 2128 38264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47944 2128 48264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 32944 2128 33264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 42944 2128 43264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 45834 0 45890 800 6 bottom_width_0_height_0_subtile_0__pin_cout_0_
port 3 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 bottom_width_0_height_0_subtile_0__pin_reg_out_0_
port 4 nsew signal output
rlabel metal3 s 50200 1232 51000 1352 6 ccff_head_0_0
port 5 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 ccff_head_1
port 6 nsew signal input
rlabel metal2 s 47490 56200 47546 57000 6 ccff_head_2
port 7 nsew signal input
rlabel metal3 s 50200 55632 51000 55752 6 ccff_tail
port 8 nsew signal output
rlabel metal2 s 3330 56200 3386 57000 6 ccff_tail_0
port 9 nsew signal output
rlabel metal3 s 50200 53456 51000 53576 6 ccff_tail_1
port 10 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 chanx_left_in[0]
port 11 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[10]
port 12 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 chanx_left_in[11]
port 13 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[12]
port 14 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_in[13]
port 15 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 chanx_left_in[14]
port 16 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 chanx_left_in[15]
port 17 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 chanx_left_in[16]
port 18 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 chanx_left_in[17]
port 19 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 chanx_left_in[18]
port 20 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 chanx_left_in[19]
port 21 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[1]
port 22 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 chanx_left_in[20]
port 23 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 chanx_left_in[21]
port 24 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 chanx_left_in[22]
port 25 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 chanx_left_in[23]
port 26 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 chanx_left_in[24]
port 27 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 chanx_left_in[25]
port 28 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 chanx_left_in[26]
port 29 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 chanx_left_in[27]
port 30 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 chanx_left_in[28]
port 31 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 chanx_left_in[29]
port 32 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[2]
port 33 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[3]
port 34 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[4]
port 35 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[5]
port 36 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[6]
port 37 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[7]
port 38 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[8]
port 39 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[9]
port 40 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 chanx_left_out[0]
port 41 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 chanx_left_out[10]
port 42 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 chanx_left_out[11]
port 43 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 chanx_left_out[12]
port 44 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 chanx_left_out[13]
port 45 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 chanx_left_out[14]
port 46 nsew signal output
rlabel metal3 s 0 35504 800 35624 6 chanx_left_out[15]
port 47 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 chanx_left_out[16]
port 48 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 chanx_left_out[17]
port 49 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 chanx_left_out[18]
port 50 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 chanx_left_out[19]
port 51 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 chanx_left_out[1]
port 52 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 chanx_left_out[20]
port 53 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 chanx_left_out[21]
port 54 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 chanx_left_out[22]
port 55 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 chanx_left_out[23]
port 56 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 chanx_left_out[24]
port 57 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 chanx_left_out[25]
port 58 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 chanx_left_out[26]
port 59 nsew signal output
rlabel metal3 s 0 43664 800 43784 6 chanx_left_out[27]
port 60 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 chanx_left_out[28]
port 61 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 chanx_left_out[29]
port 62 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 chanx_left_out[2]
port 63 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 chanx_left_out[3]
port 64 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 chanx_left_out[4]
port 65 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 chanx_left_out[5]
port 66 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 chanx_left_out[6]
port 67 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 chanx_left_out[7]
port 68 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 chanx_left_out[8]
port 69 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 chanx_left_out[9]
port 70 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[0]
port 71 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[10]
port 72 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[11]
port 73 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[12]
port 74 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[13]
port 75 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_in[14]
port 76 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[15]
port 77 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_in[16]
port 78 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_in[17]
port 79 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_in[18]
port 80 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_in[19]
port 81 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_in[1]
port 82 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_in[20]
port 83 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_in[21]
port 84 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_in[22]
port 85 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_in[23]
port 86 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 chany_bottom_in[24]
port 87 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_in[25]
port 88 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_in[26]
port 89 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_in[27]
port 90 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_in[28]
port 91 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_in[29]
port 92 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[2]
port 93 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[3]
port 94 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 chany_bottom_in[4]
port 95 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[5]
port 96 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[6]
port 97 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[7]
port 98 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[8]
port 99 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in[9]
port 100 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[0]
port 101 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 chany_bottom_out[10]
port 102 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 chany_bottom_out[11]
port 103 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 chany_bottom_out[12]
port 104 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 chany_bottom_out[13]
port 105 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 chany_bottom_out[14]
port 106 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 chany_bottom_out[15]
port 107 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 chany_bottom_out[16]
port 108 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 chany_bottom_out[17]
port 109 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 chany_bottom_out[18]
port 110 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 chany_bottom_out[19]
port 111 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[1]
port 112 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 chany_bottom_out[20]
port 113 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 chany_bottom_out[21]
port 114 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 chany_bottom_out[22]
port 115 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 chany_bottom_out[23]
port 116 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 chany_bottom_out[24]
port 117 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 chany_bottom_out[25]
port 118 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 chany_bottom_out[26]
port 119 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 chany_bottom_out[27]
port 120 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 chany_bottom_out[28]
port 121 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 chany_bottom_out[29]
port 122 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[2]
port 123 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[3]
port 124 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 chany_bottom_out[4]
port 125 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 chany_bottom_out[5]
port 126 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 chany_bottom_out[6]
port 127 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 chany_bottom_out[7]
port 128 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 chany_bottom_out[8]
port 129 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 chany_bottom_out[9]
port 130 nsew signal output
rlabel metal2 s 20442 56200 20498 57000 6 chany_top_in_0[0]
port 131 nsew signal input
rlabel metal2 s 25962 56200 26018 57000 6 chany_top_in_0[10]
port 132 nsew signal input
rlabel metal2 s 26514 56200 26570 57000 6 chany_top_in_0[11]
port 133 nsew signal input
rlabel metal2 s 27066 56200 27122 57000 6 chany_top_in_0[12]
port 134 nsew signal input
rlabel metal2 s 27618 56200 27674 57000 6 chany_top_in_0[13]
port 135 nsew signal input
rlabel metal2 s 28170 56200 28226 57000 6 chany_top_in_0[14]
port 136 nsew signal input
rlabel metal2 s 28722 56200 28778 57000 6 chany_top_in_0[15]
port 137 nsew signal input
rlabel metal2 s 29274 56200 29330 57000 6 chany_top_in_0[16]
port 138 nsew signal input
rlabel metal2 s 29826 56200 29882 57000 6 chany_top_in_0[17]
port 139 nsew signal input
rlabel metal2 s 30378 56200 30434 57000 6 chany_top_in_0[18]
port 140 nsew signal input
rlabel metal2 s 30930 56200 30986 57000 6 chany_top_in_0[19]
port 141 nsew signal input
rlabel metal2 s 20994 56200 21050 57000 6 chany_top_in_0[1]
port 142 nsew signal input
rlabel metal2 s 31482 56200 31538 57000 6 chany_top_in_0[20]
port 143 nsew signal input
rlabel metal2 s 32034 56200 32090 57000 6 chany_top_in_0[21]
port 144 nsew signal input
rlabel metal2 s 32586 56200 32642 57000 6 chany_top_in_0[22]
port 145 nsew signal input
rlabel metal2 s 33138 56200 33194 57000 6 chany_top_in_0[23]
port 146 nsew signal input
rlabel metal2 s 33690 56200 33746 57000 6 chany_top_in_0[24]
port 147 nsew signal input
rlabel metal2 s 34242 56200 34298 57000 6 chany_top_in_0[25]
port 148 nsew signal input
rlabel metal2 s 34794 56200 34850 57000 6 chany_top_in_0[26]
port 149 nsew signal input
rlabel metal2 s 35346 56200 35402 57000 6 chany_top_in_0[27]
port 150 nsew signal input
rlabel metal2 s 35898 56200 35954 57000 6 chany_top_in_0[28]
port 151 nsew signal input
rlabel metal2 s 36450 56200 36506 57000 6 chany_top_in_0[29]
port 152 nsew signal input
rlabel metal2 s 21546 56200 21602 57000 6 chany_top_in_0[2]
port 153 nsew signal input
rlabel metal2 s 22098 56200 22154 57000 6 chany_top_in_0[3]
port 154 nsew signal input
rlabel metal2 s 22650 56200 22706 57000 6 chany_top_in_0[4]
port 155 nsew signal input
rlabel metal2 s 23202 56200 23258 57000 6 chany_top_in_0[5]
port 156 nsew signal input
rlabel metal2 s 23754 56200 23810 57000 6 chany_top_in_0[6]
port 157 nsew signal input
rlabel metal2 s 24306 56200 24362 57000 6 chany_top_in_0[7]
port 158 nsew signal input
rlabel metal2 s 24858 56200 24914 57000 6 chany_top_in_0[8]
port 159 nsew signal input
rlabel metal2 s 25410 56200 25466 57000 6 chany_top_in_0[9]
port 160 nsew signal input
rlabel metal2 s 3882 56200 3938 57000 6 chany_top_out_0[0]
port 161 nsew signal output
rlabel metal2 s 9402 56200 9458 57000 6 chany_top_out_0[10]
port 162 nsew signal output
rlabel metal2 s 9954 56200 10010 57000 6 chany_top_out_0[11]
port 163 nsew signal output
rlabel metal2 s 10506 56200 10562 57000 6 chany_top_out_0[12]
port 164 nsew signal output
rlabel metal2 s 11058 56200 11114 57000 6 chany_top_out_0[13]
port 165 nsew signal output
rlabel metal2 s 11610 56200 11666 57000 6 chany_top_out_0[14]
port 166 nsew signal output
rlabel metal2 s 12162 56200 12218 57000 6 chany_top_out_0[15]
port 167 nsew signal output
rlabel metal2 s 12714 56200 12770 57000 6 chany_top_out_0[16]
port 168 nsew signal output
rlabel metal2 s 13266 56200 13322 57000 6 chany_top_out_0[17]
port 169 nsew signal output
rlabel metal2 s 13818 56200 13874 57000 6 chany_top_out_0[18]
port 170 nsew signal output
rlabel metal2 s 14370 56200 14426 57000 6 chany_top_out_0[19]
port 171 nsew signal output
rlabel metal2 s 4434 56200 4490 57000 6 chany_top_out_0[1]
port 172 nsew signal output
rlabel metal2 s 14922 56200 14978 57000 6 chany_top_out_0[20]
port 173 nsew signal output
rlabel metal2 s 15474 56200 15530 57000 6 chany_top_out_0[21]
port 174 nsew signal output
rlabel metal2 s 16026 56200 16082 57000 6 chany_top_out_0[22]
port 175 nsew signal output
rlabel metal2 s 16578 56200 16634 57000 6 chany_top_out_0[23]
port 176 nsew signal output
rlabel metal2 s 17130 56200 17186 57000 6 chany_top_out_0[24]
port 177 nsew signal output
rlabel metal2 s 17682 56200 17738 57000 6 chany_top_out_0[25]
port 178 nsew signal output
rlabel metal2 s 18234 56200 18290 57000 6 chany_top_out_0[26]
port 179 nsew signal output
rlabel metal2 s 18786 56200 18842 57000 6 chany_top_out_0[27]
port 180 nsew signal output
rlabel metal2 s 19338 56200 19394 57000 6 chany_top_out_0[28]
port 181 nsew signal output
rlabel metal2 s 19890 56200 19946 57000 6 chany_top_out_0[29]
port 182 nsew signal output
rlabel metal2 s 4986 56200 5042 57000 6 chany_top_out_0[2]
port 183 nsew signal output
rlabel metal2 s 5538 56200 5594 57000 6 chany_top_out_0[3]
port 184 nsew signal output
rlabel metal2 s 6090 56200 6146 57000 6 chany_top_out_0[4]
port 185 nsew signal output
rlabel metal2 s 6642 56200 6698 57000 6 chany_top_out_0[5]
port 186 nsew signal output
rlabel metal2 s 7194 56200 7250 57000 6 chany_top_out_0[6]
port 187 nsew signal output
rlabel metal2 s 7746 56200 7802 57000 6 chany_top_out_0[7]
port 188 nsew signal output
rlabel metal2 s 8298 56200 8354 57000 6 chany_top_out_0[8]
port 189 nsew signal output
rlabel metal2 s 8850 56200 8906 57000 6 chany_top_out_0[9]
port 190 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 clk0
port 191 nsew signal input
rlabel metal3 s 50200 12112 51000 12232 6 gfpga_pad_io_soc_dir[0]
port 192 nsew signal output
rlabel metal3 s 50200 14288 51000 14408 6 gfpga_pad_io_soc_dir[1]
port 193 nsew signal output
rlabel metal3 s 50200 16464 51000 16584 6 gfpga_pad_io_soc_dir[2]
port 194 nsew signal output
rlabel metal3 s 50200 18640 51000 18760 6 gfpga_pad_io_soc_dir[3]
port 195 nsew signal output
rlabel metal3 s 50200 29520 51000 29640 6 gfpga_pad_io_soc_in[0]
port 196 nsew signal input
rlabel metal3 s 50200 31696 51000 31816 6 gfpga_pad_io_soc_in[1]
port 197 nsew signal input
rlabel metal3 s 50200 33872 51000 33992 6 gfpga_pad_io_soc_in[2]
port 198 nsew signal input
rlabel metal3 s 50200 36048 51000 36168 6 gfpga_pad_io_soc_in[3]
port 199 nsew signal input
rlabel metal3 s 50200 20816 51000 20936 6 gfpga_pad_io_soc_out[0]
port 200 nsew signal output
rlabel metal3 s 50200 22992 51000 23112 6 gfpga_pad_io_soc_out[1]
port 201 nsew signal output
rlabel metal3 s 50200 25168 51000 25288 6 gfpga_pad_io_soc_out[2]
port 202 nsew signal output
rlabel metal3 s 50200 27344 51000 27464 6 gfpga_pad_io_soc_out[3]
port 203 nsew signal output
rlabel metal3 s 50200 38224 51000 38344 6 isol_n
port 204 nsew signal input
rlabel metal3 s 50200 3408 51000 3528 6 left_width_0_height_0_subtile_0__pin_inpad_0_
port 205 nsew signal output
rlabel metal3 s 50200 5584 51000 5704 6 left_width_0_height_0_subtile_1__pin_inpad_0_
port 206 nsew signal output
rlabel metal3 s 50200 7760 51000 7880 6 left_width_0_height_0_subtile_2__pin_inpad_0_
port 207 nsew signal output
rlabel metal3 s 50200 9936 51000 10056 6 left_width_0_height_0_subtile_3__pin_inpad_0_
port 208 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 prog_clk
port 209 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 prog_reset_bottom_in
port 210 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 prog_reset_bottom_out
port 211 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 prog_reset_left_in
port 212 nsew signal input
rlabel metal2 s 38658 56200 38714 57000 6 prog_reset_top_in
port 213 nsew signal input
rlabel metal2 s 38106 56200 38162 57000 6 prog_reset_top_out
port 214 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 reset_bottom_in
port 215 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 reset_bottom_out
port 216 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 reset_left_out
port 217 nsew signal output
rlabel metal3 s 50200 42576 51000 42696 6 reset_right_in
port 218 nsew signal input
rlabel metal2 s 39762 56200 39818 57000 6 reset_top_in
port 219 nsew signal input
rlabel metal2 s 39210 56200 39266 57000 6 reset_top_out
port 220 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 right_width_0_height_0_subtile_0__pin_O_10_
port 221 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 right_width_0_height_0_subtile_0__pin_O_11_
port 222 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 right_width_0_height_0_subtile_0__pin_O_12_
port 223 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 right_width_0_height_0_subtile_0__pin_O_13_
port 224 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 right_width_0_height_0_subtile_0__pin_O_14_
port 225 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 right_width_0_height_0_subtile_0__pin_O_15_
port 226 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 right_width_0_height_0_subtile_0__pin_O_8_
port 227 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 right_width_0_height_0_subtile_0__pin_O_9_
port 228 nsew signal output
rlabel metal2 s 46938 56200 46994 57000 6 sc_in
port 229 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 sc_out
port 230 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 test_enable_bottom_in
port 231 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 test_enable_bottom_out
port 232 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 test_enable_left_out
port 233 nsew signal output
rlabel metal3 s 50200 40400 51000 40520 6 test_enable_right_in
port 234 nsew signal input
rlabel metal2 s 40866 56200 40922 57000 6 test_enable_top_in
port 235 nsew signal input
rlabel metal2 s 40314 56200 40370 57000 6 test_enable_top_out
port 236 nsew signal output
rlabel metal2 s 42522 56200 42578 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 237 nsew signal input
rlabel metal2 s 43074 56200 43130 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 238 nsew signal input
rlabel metal2 s 43626 56200 43682 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 239 nsew signal input
rlabel metal2 s 44178 56200 44234 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 240 nsew signal input
rlabel metal2 s 44730 56200 44786 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 241 nsew signal input
rlabel metal2 s 45282 56200 45338 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 242 nsew signal input
rlabel metal2 s 41418 56200 41474 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 243 nsew signal input
rlabel metal2 s 41970 56200 42026 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 244 nsew signal input
rlabel metal3 s 50200 44752 51000 44872 6 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 245 nsew signal input
rlabel metal3 s 50200 46928 51000 47048 6 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 246 nsew signal input
rlabel metal3 s 50200 49104 51000 49224 6 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 247 nsew signal input
rlabel metal3 s 50200 51280 51000 51400 6 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 248 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 top_width_0_height_0_subtile_0__pin_O_0_
port 249 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 top_width_0_height_0_subtile_0__pin_O_1_
port 250 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 top_width_0_height_0_subtile_0__pin_O_2_
port 251 nsew signal output
rlabel metal3 s 0 49104 800 49224 6 top_width_0_height_0_subtile_0__pin_O_3_
port 252 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 top_width_0_height_0_subtile_0__pin_O_4_
port 253 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 top_width_0_height_0_subtile_0__pin_O_5_
port 254 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 top_width_0_height_0_subtile_0__pin_O_6_
port 255 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 top_width_0_height_0_subtile_0__pin_O_7_
port 256 nsew signal output
rlabel metal2 s 45834 56200 45890 57000 6 top_width_0_height_0_subtile_0__pin_cin_0_
port 257 nsew signal input
rlabel metal2 s 46386 56200 46442 57000 6 top_width_0_height_0_subtile_0__pin_reg_in_0_
port 258 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 51000 57000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6792272
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/right_tile/runs/23_03_20_06_27/results/signoff/right_tile.magic.gds
string GDS_START 250542
<< end >>

