magic
tech sky130A
magscale 1 2
timestamp 1656943349
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 382 1912 22618 21072
<< metal2 >>
rect 386 22200 442 23000
rect 938 22200 994 23000
rect 1490 22200 1546 23000
rect 2042 22200 2098 23000
rect 2594 22200 2650 23000
rect 3146 22200 3202 23000
rect 3698 22200 3754 23000
rect 4250 22200 4306 23000
rect 4802 22200 4858 23000
rect 5354 22200 5410 23000
rect 5906 22200 5962 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 11978 22200 12034 23000
rect 12530 22200 12586 23000
rect 13082 22200 13138 23000
rect 13634 22200 13690 23000
rect 14186 22200 14242 23000
rect 14738 22200 14794 23000
rect 15290 22200 15346 23000
rect 15842 22200 15898 23000
rect 16394 22200 16450 23000
rect 16946 22200 17002 23000
rect 17498 22200 17554 23000
rect 18050 22200 18106 23000
rect 18602 22200 18658 23000
rect 19154 22200 19210 23000
rect 19706 22200 19762 23000
rect 20258 22200 20314 23000
rect 20810 22200 20866 23000
rect 21362 22200 21418 23000
rect 21914 22200 21970 23000
rect 22466 22200 22522 23000
rect 386 0 442 800
rect 938 0 994 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
<< obsm2 >>
rect 498 22144 882 22250
rect 1050 22144 1434 22250
rect 1602 22144 1986 22250
rect 2154 22144 2538 22250
rect 2706 22144 3090 22250
rect 3258 22144 3642 22250
rect 3810 22144 4194 22250
rect 4362 22144 4746 22250
rect 4914 22144 5298 22250
rect 5466 22144 5850 22250
rect 6018 22144 6402 22250
rect 6570 22144 6954 22250
rect 7122 22144 7506 22250
rect 7674 22144 8058 22250
rect 8226 22144 8610 22250
rect 8778 22144 9162 22250
rect 9330 22144 9714 22250
rect 9882 22144 10266 22250
rect 10434 22144 10818 22250
rect 10986 22144 11370 22250
rect 11538 22144 11922 22250
rect 12090 22144 12474 22250
rect 12642 22144 13026 22250
rect 13194 22144 13578 22250
rect 13746 22144 14130 22250
rect 14298 22144 14682 22250
rect 14850 22144 15234 22250
rect 15402 22144 15786 22250
rect 15954 22144 16338 22250
rect 16506 22144 16890 22250
rect 17058 22144 17442 22250
rect 17610 22144 17994 22250
rect 18162 22144 18546 22250
rect 18714 22144 19098 22250
rect 19266 22144 19650 22250
rect 19818 22144 20202 22250
rect 20370 22144 20754 22250
rect 20922 22144 21306 22250
rect 21474 22144 21858 22250
rect 22026 22144 22410 22250
rect 22578 22144 22612 22250
rect 386 856 22612 22144
rect 498 734 882 856
rect 1050 734 1434 856
rect 1602 734 1986 856
rect 2154 734 2538 856
rect 2706 734 3090 856
rect 3258 734 3642 856
rect 3810 734 4194 856
rect 4362 734 4746 856
rect 4914 734 5298 856
rect 5466 734 5850 856
rect 6018 734 6402 856
rect 6570 734 6954 856
rect 7122 734 7506 856
rect 7674 734 8058 856
rect 8226 734 8610 856
rect 8778 734 9162 856
rect 9330 734 9714 856
rect 9882 734 10266 856
rect 10434 734 10818 856
rect 10986 734 11370 856
rect 11538 734 11922 856
rect 12090 734 12474 856
rect 12642 734 13026 856
rect 13194 734 13578 856
rect 13746 734 14130 856
rect 14298 734 14682 856
rect 14850 734 15234 856
rect 15402 734 15786 856
rect 15954 734 16338 856
rect 16506 734 16890 856
rect 17058 734 17442 856
rect 17610 734 17994 856
rect 18162 734 18546 856
rect 18714 734 19098 856
rect 19266 734 19650 856
rect 19818 734 20202 856
rect 20370 734 20754 856
rect 20922 734 21306 856
rect 21474 734 21858 856
rect 22026 734 22410 856
rect 22578 734 22612 856
<< metal3 >>
rect 22200 21224 23000 21344
rect 22200 20816 23000 20936
rect 22200 20408 23000 20528
rect 22200 20000 23000 20120
rect 22200 19592 23000 19712
rect 22200 19184 23000 19304
rect 22200 18776 23000 18896
rect 22200 18368 23000 18488
rect 22200 17960 23000 18080
rect 22200 17552 23000 17672
rect 0 17144 800 17264
rect 22200 17144 23000 17264
rect 22200 16736 23000 16856
rect 22200 16328 23000 16448
rect 22200 15920 23000 16040
rect 22200 15512 23000 15632
rect 22200 15104 23000 15224
rect 22200 14696 23000 14816
rect 22200 14288 23000 14408
rect 22200 13880 23000 14000
rect 22200 13472 23000 13592
rect 22200 13064 23000 13184
rect 22200 12656 23000 12776
rect 22200 12248 23000 12368
rect 22200 11840 23000 11960
rect 22200 11432 23000 11552
rect 22200 11024 23000 11144
rect 22200 10616 23000 10736
rect 22200 10208 23000 10328
rect 22200 9800 23000 9920
rect 22200 9392 23000 9512
rect 22200 8984 23000 9104
rect 22200 8576 23000 8696
rect 22200 8168 23000 8288
rect 22200 7760 23000 7880
rect 22200 7352 23000 7472
rect 22200 6944 23000 7064
rect 22200 6536 23000 6656
rect 22200 6128 23000 6248
rect 0 5720 800 5840
rect 22200 5720 23000 5840
rect 22200 5312 23000 5432
rect 22200 4904 23000 5024
rect 22200 4496 23000 4616
rect 22200 4088 23000 4208
rect 22200 3680 23000 3800
rect 22200 3272 23000 3392
rect 22200 2864 23000 2984
rect 22200 2456 23000 2576
rect 22200 2048 23000 2168
rect 22200 1640 23000 1760
<< obsm3 >>
rect 381 21144 22120 21317
rect 381 21016 22202 21144
rect 381 20736 22120 21016
rect 381 20608 22202 20736
rect 381 20328 22120 20608
rect 381 20200 22202 20328
rect 381 19920 22120 20200
rect 381 19792 22202 19920
rect 381 19512 22120 19792
rect 381 19384 22202 19512
rect 381 19104 22120 19384
rect 381 18976 22202 19104
rect 381 18696 22120 18976
rect 381 18568 22202 18696
rect 381 18288 22120 18568
rect 381 18160 22202 18288
rect 381 17880 22120 18160
rect 381 17752 22202 17880
rect 381 17472 22120 17752
rect 381 17344 22202 17472
rect 880 17064 22120 17344
rect 381 16936 22202 17064
rect 381 16656 22120 16936
rect 381 16528 22202 16656
rect 381 16248 22120 16528
rect 381 16120 22202 16248
rect 381 15840 22120 16120
rect 381 15712 22202 15840
rect 381 15432 22120 15712
rect 381 15304 22202 15432
rect 381 15024 22120 15304
rect 381 14896 22202 15024
rect 381 14616 22120 14896
rect 381 14488 22202 14616
rect 381 14208 22120 14488
rect 381 14080 22202 14208
rect 381 13800 22120 14080
rect 381 13672 22202 13800
rect 381 13392 22120 13672
rect 381 13264 22202 13392
rect 381 12984 22120 13264
rect 381 12856 22202 12984
rect 381 12576 22120 12856
rect 381 12448 22202 12576
rect 381 12168 22120 12448
rect 381 12040 22202 12168
rect 381 11760 22120 12040
rect 381 11632 22202 11760
rect 381 11352 22120 11632
rect 381 11224 22202 11352
rect 381 10944 22120 11224
rect 381 10816 22202 10944
rect 381 10536 22120 10816
rect 381 10408 22202 10536
rect 381 10128 22120 10408
rect 381 10000 22202 10128
rect 381 9720 22120 10000
rect 381 9592 22202 9720
rect 381 9312 22120 9592
rect 381 9184 22202 9312
rect 381 8904 22120 9184
rect 381 8776 22202 8904
rect 381 8496 22120 8776
rect 381 8368 22202 8496
rect 381 8088 22120 8368
rect 381 7960 22202 8088
rect 381 7680 22120 7960
rect 381 7552 22202 7680
rect 381 7272 22120 7552
rect 381 7144 22202 7272
rect 381 6864 22120 7144
rect 381 6736 22202 6864
rect 381 6456 22120 6736
rect 381 6328 22202 6456
rect 381 6048 22120 6328
rect 381 5920 22202 6048
rect 880 5640 22120 5920
rect 381 5512 22202 5640
rect 381 5232 22120 5512
rect 381 5104 22202 5232
rect 381 4824 22120 5104
rect 381 4696 22202 4824
rect 381 4416 22120 4696
rect 381 4288 22202 4416
rect 381 4008 22120 4288
rect 381 3880 22202 4008
rect 381 3600 22120 3880
rect 381 3472 22202 3600
rect 381 3192 22120 3472
rect 381 3064 22202 3192
rect 381 2784 22120 3064
rect 381 2656 22202 2784
rect 381 2376 22120 2656
rect 381 2248 22202 2376
rect 381 1968 22120 2248
rect 381 1840 22202 1968
rect 381 1667 22120 1840
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 5947 3027 6062 20229
rect 6542 3027 8661 20229
rect 9141 3027 11260 20229
rect 11740 3027 13859 20229
rect 14339 3027 16458 20229
rect 16938 3027 19057 20229
rect 19537 3027 20365 20229
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 386 0 442 800 6 bottom_left_grid_pin_1_
port 3 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 4 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 5 nsew signal output
rlabel metal3 s 22200 4904 23000 5024 6 chanx_right_in[0]
port 6 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[10]
port 7 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[11]
port 8 nsew signal input
rlabel metal3 s 22200 9800 23000 9920 6 chanx_right_in[12]
port 9 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[13]
port 10 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[14]
port 11 nsew signal input
rlabel metal3 s 22200 11024 23000 11144 6 chanx_right_in[15]
port 12 nsew signal input
rlabel metal3 s 22200 11432 23000 11552 6 chanx_right_in[16]
port 13 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 14 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 15 nsew signal input
rlabel metal3 s 22200 12656 23000 12776 6 chanx_right_in[19]
port 16 nsew signal input
rlabel metal3 s 22200 5312 23000 5432 6 chanx_right_in[1]
port 17 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[2]
port 18 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[3]
port 19 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[4]
port 20 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[5]
port 21 nsew signal input
rlabel metal3 s 22200 7352 23000 7472 6 chanx_right_in[6]
port 22 nsew signal input
rlabel metal3 s 22200 7760 23000 7880 6 chanx_right_in[7]
port 23 nsew signal input
rlabel metal3 s 22200 8168 23000 8288 6 chanx_right_in[8]
port 24 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[9]
port 25 nsew signal input
rlabel metal3 s 22200 13064 23000 13184 6 chanx_right_out[0]
port 26 nsew signal output
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[10]
port 27 nsew signal output
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[11]
port 28 nsew signal output
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[12]
port 29 nsew signal output
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[13]
port 30 nsew signal output
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[14]
port 31 nsew signal output
rlabel metal3 s 22200 19184 23000 19304 6 chanx_right_out[15]
port 32 nsew signal output
rlabel metal3 s 22200 19592 23000 19712 6 chanx_right_out[16]
port 33 nsew signal output
rlabel metal3 s 22200 20000 23000 20120 6 chanx_right_out[17]
port 34 nsew signal output
rlabel metal3 s 22200 20408 23000 20528 6 chanx_right_out[18]
port 35 nsew signal output
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[19]
port 36 nsew signal output
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[1]
port 37 nsew signal output
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[2]
port 38 nsew signal output
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[3]
port 39 nsew signal output
rlabel metal3 s 22200 14696 23000 14816 6 chanx_right_out[4]
port 40 nsew signal output
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[5]
port 41 nsew signal output
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[6]
port 42 nsew signal output
rlabel metal3 s 22200 15920 23000 16040 6 chanx_right_out[7]
port 43 nsew signal output
rlabel metal3 s 22200 16328 23000 16448 6 chanx_right_out[8]
port 44 nsew signal output
rlabel metal3 s 22200 16736 23000 16856 6 chanx_right_out[9]
port 45 nsew signal output
rlabel metal2 s 938 0 994 800 6 chany_bottom_in[0]
port 46 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[10]
port 47 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_in[11]
port 48 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[12]
port 49 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[13]
port 50 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[14]
port 51 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[15]
port 52 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[16]
port 53 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[17]
port 54 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[18]
port 55 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[19]
port 56 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 chany_bottom_in[1]
port 57 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 chany_bottom_in[2]
port 58 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 chany_bottom_in[3]
port 59 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_in[4]
port 60 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[5]
port 61 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[6]
port 62 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_in[7]
port 63 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[8]
port 64 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[9]
port 65 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 chany_bottom_out[0]
port 66 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[10]
port 67 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 chany_bottom_out[11]
port 68 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[12]
port 69 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[13]
port 70 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 chany_bottom_out[14]
port 71 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[15]
port 72 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[16]
port 73 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[17]
port 74 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 chany_bottom_out[18]
port 75 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 chany_bottom_out[19]
port 76 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[1]
port 77 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[2]
port 78 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 chany_bottom_out[3]
port 79 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 chany_bottom_out[4]
port 80 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[5]
port 81 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 chany_bottom_out[6]
port 82 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[7]
port 83 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[8]
port 84 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[9]
port 85 nsew signal output
rlabel metal2 s 938 22200 994 23000 6 chany_top_in[0]
port 86 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 87 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 88 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 89 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 90 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 91 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 92 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 93 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 94 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 95 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 96 nsew signal input
rlabel metal2 s 1490 22200 1546 23000 6 chany_top_in[1]
port 97 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 chany_top_in[2]
port 98 nsew signal input
rlabel metal2 s 2594 22200 2650 23000 6 chany_top_in[3]
port 99 nsew signal input
rlabel metal2 s 3146 22200 3202 23000 6 chany_top_in[4]
port 100 nsew signal input
rlabel metal2 s 3698 22200 3754 23000 6 chany_top_in[5]
port 101 nsew signal input
rlabel metal2 s 4250 22200 4306 23000 6 chany_top_in[6]
port 102 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[7]
port 103 nsew signal input
rlabel metal2 s 5354 22200 5410 23000 6 chany_top_in[8]
port 104 nsew signal input
rlabel metal2 s 5906 22200 5962 23000 6 chany_top_in[9]
port 105 nsew signal input
rlabel metal2 s 11978 22200 12034 23000 6 chany_top_out[0]
port 106 nsew signal output
rlabel metal2 s 17498 22200 17554 23000 6 chany_top_out[10]
port 107 nsew signal output
rlabel metal2 s 18050 22200 18106 23000 6 chany_top_out[11]
port 108 nsew signal output
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 109 nsew signal output
rlabel metal2 s 19154 22200 19210 23000 6 chany_top_out[13]
port 110 nsew signal output
rlabel metal2 s 19706 22200 19762 23000 6 chany_top_out[14]
port 111 nsew signal output
rlabel metal2 s 20258 22200 20314 23000 6 chany_top_out[15]
port 112 nsew signal output
rlabel metal2 s 20810 22200 20866 23000 6 chany_top_out[16]
port 113 nsew signal output
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[17]
port 114 nsew signal output
rlabel metal2 s 21914 22200 21970 23000 6 chany_top_out[18]
port 115 nsew signal output
rlabel metal2 s 22466 22200 22522 23000 6 chany_top_out[19]
port 116 nsew signal output
rlabel metal2 s 12530 22200 12586 23000 6 chany_top_out[1]
port 117 nsew signal output
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[2]
port 118 nsew signal output
rlabel metal2 s 13634 22200 13690 23000 6 chany_top_out[3]
port 119 nsew signal output
rlabel metal2 s 14186 22200 14242 23000 6 chany_top_out[4]
port 120 nsew signal output
rlabel metal2 s 14738 22200 14794 23000 6 chany_top_out[5]
port 121 nsew signal output
rlabel metal2 s 15290 22200 15346 23000 6 chany_top_out[6]
port 122 nsew signal output
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[7]
port 123 nsew signal output
rlabel metal2 s 16394 22200 16450 23000 6 chany_top_out[8]
port 124 nsew signal output
rlabel metal2 s 16946 22200 17002 23000 6 chany_top_out[9]
port 125 nsew signal output
rlabel metal3 s 22200 21224 23000 21344 6 prog_clk_0_E_in
port 126 nsew signal input
rlabel metal3 s 22200 1640 23000 1760 6 right_bottom_grid_pin_34_
port 127 nsew signal input
rlabel metal3 s 22200 2048 23000 2168 6 right_bottom_grid_pin_35_
port 128 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_36_
port 129 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_37_
port 130 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_38_
port 131 nsew signal input
rlabel metal3 s 22200 3680 23000 3800 6 right_bottom_grid_pin_39_
port 132 nsew signal input
rlabel metal3 s 22200 4088 23000 4208 6 right_bottom_grid_pin_40_
port 133 nsew signal input
rlabel metal3 s 22200 4496 23000 4616 6 right_bottom_grid_pin_41_
port 134 nsew signal input
rlabel metal2 s 386 22200 442 23000 6 top_left_grid_pin_1_
port 135 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1390320
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_0__1_/runs/sb_0__1_/results/signoff/sb_0__1_.magic.gds
string GDS_START 65026
<< end >>

