magic
tech sky130A
magscale 1 2
timestamp 1625785457
<< obsli1 >>
rect 1104 2159 10856 11441
<< obsm1 >>
rect 750 2128 11210 11472
<< metal2 >>
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
<< obsm2 >>
rect 756 856 11204 11472
rect 866 800 2170 856
rect 2338 800 3642 856
rect 3810 800 5114 856
rect 5282 800 6678 856
rect 6846 800 8150 856
rect 8318 800 9622 856
rect 9790 800 11094 856
<< obsm3 >>
rect 2576 2143 9424 11457
<< metal4 >>
rect 2576 2128 2896 11472
rect 4208 2128 4528 11472
rect 5840 2128 6160 11472
rect 7472 2128 7792 11472
rect 9104 2128 9424 11472
<< labels >>
rlabel metal2 s 754 0 810 800 6 x[0]
port 1 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 x[1]
port 2 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 x[2]
port 3 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 x[3]
port 4 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 x[4]
port 5 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 x[5]
port 6 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 x[6]
port 7 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 x[7]
port 8 nsew signal output
rlabel metal4 s 9104 2128 9424 11472 6 VPWR
port 9 nsew power bidirectional
rlabel metal4 s 5840 2128 6160 11472 6 VPWR
port 10 nsew power bidirectional
rlabel metal4 s 2576 2128 2896 11472 6 VPWR
port 11 nsew power bidirectional
rlabel metal4 s 7472 2128 7792 11472 6 VGND
port 12 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 11472 6 VGND
port 13 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 12000 14000
string LEFview TRUE
string GDS_FILE /project/openlane/tie_array/runs/tie_array/results/magic/tie_array.gds
string GDS_END 105894
string GDS_START 28708
<< end >>

