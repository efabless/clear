magic
tech sky130A
magscale 1 2
timestamp 1681685601
<< viali >>
rect 1593 24361 1627 24395
rect 14381 24361 14415 24395
rect 16957 24361 16991 24395
rect 21833 24361 21867 24395
rect 11713 24293 11747 24327
rect 15577 24293 15611 24327
rect 18153 24293 18187 24327
rect 3249 24225 3283 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 12817 24225 12851 24259
rect 15025 24225 15059 24259
rect 16221 24225 16255 24259
rect 17417 24225 17451 24259
rect 17509 24225 17543 24259
rect 18705 24225 18739 24259
rect 25237 24225 25271 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7205 24157 7239 24191
rect 9781 24157 9815 24191
rect 11897 24157 11931 24191
rect 12449 24157 12483 24191
rect 18521 24157 18555 24191
rect 18613 24157 18647 24191
rect 20177 24157 20211 24191
rect 20545 24157 20579 24191
rect 21465 24157 21499 24191
rect 22293 24157 22327 24191
rect 24961 24157 24995 24191
rect 1685 24089 1719 24123
rect 5825 24089 5859 24123
rect 16037 24089 16071 24123
rect 22569 24089 22603 24123
rect 3985 24021 4019 24055
rect 6561 24021 6595 24055
rect 9137 24021 9171 24055
rect 14749 24021 14783 24055
rect 14841 24021 14875 24055
rect 15945 24021 15979 24055
rect 17325 24021 17359 24055
rect 19441 24021 19475 24055
rect 21281 24021 21315 24055
rect 24041 24021 24075 24055
rect 24593 24021 24627 24055
rect 25053 24021 25087 24055
rect 16681 23817 16715 23851
rect 16865 23817 16899 23851
rect 3985 23749 4019 23783
rect 5825 23749 5859 23783
rect 9137 23749 9171 23783
rect 10885 23749 10919 23783
rect 15945 23749 15979 23783
rect 16037 23749 16071 23783
rect 17325 23749 17359 23783
rect 20085 23749 20119 23783
rect 21833 23749 21867 23783
rect 24593 23749 24627 23783
rect 25145 23749 25179 23783
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6837 23681 6871 23715
rect 7941 23681 7975 23715
rect 9781 23681 9815 23715
rect 12081 23681 12115 23715
rect 13921 23681 13955 23715
rect 14473 23681 14507 23715
rect 14565 23681 14599 23715
rect 17233 23681 17267 23715
rect 20637 23681 20671 23715
rect 11713 23613 11747 23647
rect 12541 23613 12575 23647
rect 14749 23613 14783 23647
rect 16221 23613 16255 23647
rect 17509 23613 17543 23647
rect 18061 23613 18095 23647
rect 18337 23613 18371 23647
rect 20913 23613 20947 23647
rect 22293 23613 22327 23647
rect 22569 23613 22603 23647
rect 24041 23613 24075 23647
rect 7481 23545 7515 23579
rect 14105 23545 14139 23579
rect 20361 23545 20395 23579
rect 25329 23545 25363 23579
rect 2329 23477 2363 23511
rect 6561 23477 6595 23511
rect 11621 23477 11655 23511
rect 13829 23477 13863 23511
rect 15209 23477 15243 23511
rect 15577 23477 15611 23511
rect 19809 23477 19843 23511
rect 24409 23477 24443 23511
rect 1777 23273 1811 23307
rect 9321 23273 9355 23307
rect 21189 23273 21223 23307
rect 23397 23273 23431 23307
rect 24409 23273 24443 23307
rect 13553 23205 13587 23239
rect 24593 23205 24627 23239
rect 1593 23137 1627 23171
rect 4261 23137 4295 23171
rect 10517 23137 10551 23171
rect 12173 23137 12207 23171
rect 15301 23137 15335 23171
rect 17785 23137 17819 23171
rect 19717 23137 19751 23171
rect 21649 23137 21683 23171
rect 25053 23137 25087 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 3985 23069 4019 23103
rect 5457 23069 5491 23103
rect 7205 23069 7239 23103
rect 8217 23069 8251 23103
rect 9873 23069 9907 23103
rect 11713 23069 11747 23103
rect 13737 23069 13771 23103
rect 15025 23069 15059 23103
rect 17601 23069 17635 23103
rect 19441 23069 19475 23103
rect 24041 23069 24075 23103
rect 3249 23001 3283 23035
rect 6561 23001 6595 23035
rect 9229 23001 9263 23035
rect 14381 23001 14415 23035
rect 18521 23001 18555 23035
rect 21925 23001 21959 23035
rect 24961 23001 24995 23035
rect 14473 22933 14507 22967
rect 16773 22933 16807 22967
rect 17233 22933 17267 22967
rect 17693 22933 17727 22967
rect 18613 22933 18647 22967
rect 19073 22933 19107 22967
rect 23857 22933 23891 22967
rect 15393 22729 15427 22763
rect 19257 22729 19291 22763
rect 21097 22729 21131 22763
rect 25053 22729 25087 22763
rect 3985 22661 4019 22695
rect 5733 22661 5767 22695
rect 6929 22661 6963 22695
rect 8769 22661 8803 22695
rect 12081 22661 12115 22695
rect 17141 22661 17175 22695
rect 19165 22661 19199 22695
rect 23581 22661 23615 22695
rect 1685 22593 1719 22627
rect 2789 22593 2823 22627
rect 4813 22593 4847 22627
rect 7573 22593 7607 22627
rect 13001 22593 13035 22627
rect 13645 22593 13679 22627
rect 15945 22593 15979 22627
rect 16865 22593 16899 22627
rect 20177 22593 20211 22627
rect 20729 22593 20763 22627
rect 7113 22525 7147 22559
rect 9413 22525 9447 22559
rect 9689 22525 9723 22559
rect 12173 22525 12207 22559
rect 12265 22525 12299 22559
rect 13921 22525 13955 22559
rect 18613 22525 18647 22559
rect 21281 22525 21315 22559
rect 22017 22525 22051 22559
rect 22293 22525 22327 22559
rect 23305 22525 23339 22559
rect 11713 22457 11747 22491
rect 16129 22457 16163 22491
rect 16497 22457 16531 22491
rect 25329 22457 25363 22491
rect 2329 22389 2363 22423
rect 6469 22389 6503 22423
rect 11161 22389 11195 22423
rect 13093 22389 13127 22423
rect 19625 22389 19659 22423
rect 21465 22389 21499 22423
rect 10964 22185 10998 22219
rect 14552 22185 14586 22219
rect 16497 22185 16531 22219
rect 18705 22185 18739 22219
rect 20618 22185 20652 22219
rect 2881 22049 2915 22083
rect 3985 22049 4019 22083
rect 6101 22049 6135 22083
rect 8309 22049 8343 22083
rect 10701 22049 10735 22083
rect 12449 22049 12483 22083
rect 17141 22049 17175 22083
rect 18245 22049 18279 22083
rect 19993 22049 20027 22083
rect 25053 22049 25087 22083
rect 25145 22049 25179 22083
rect 2237 21981 2271 22015
rect 4261 21981 4295 22015
rect 5549 21981 5583 22015
rect 7389 21981 7423 22015
rect 9137 21981 9171 22015
rect 9608 21981 9642 22015
rect 13093 21981 13127 22015
rect 14289 21981 14323 22015
rect 20361 21981 20395 22015
rect 22661 21981 22695 22015
rect 24961 21981 24995 22015
rect 1777 21913 1811 21947
rect 13737 21913 13771 21947
rect 16957 21913 16991 21947
rect 19533 21913 19567 21947
rect 19717 21913 19751 21947
rect 23581 21913 23615 21947
rect 1593 21845 1627 21879
rect 4905 21845 4939 21879
rect 9321 21845 9355 21879
rect 10241 21845 10275 21879
rect 12817 21845 12851 21879
rect 16037 21845 16071 21879
rect 16865 21845 16899 21879
rect 17693 21845 17727 21879
rect 18061 21845 18095 21879
rect 18153 21845 18187 21879
rect 18889 21845 18923 21879
rect 22109 21845 22143 21879
rect 24593 21845 24627 21879
rect 1777 21641 1811 21675
rect 12633 21641 12667 21675
rect 12725 21641 12759 21675
rect 13829 21641 13863 21675
rect 20453 21641 20487 21675
rect 22017 21641 22051 21675
rect 22385 21641 22419 21675
rect 1685 21573 1719 21607
rect 6561 21573 6595 21607
rect 11161 21573 11195 21607
rect 11989 21573 12023 21607
rect 14289 21573 14323 21607
rect 20821 21573 20855 21607
rect 20913 21573 20947 21607
rect 2973 21505 3007 21539
rect 4813 21505 4847 21539
rect 7389 21505 7423 21539
rect 9045 21505 9079 21539
rect 14197 21505 14231 21539
rect 15393 21505 15427 21539
rect 15485 21505 15519 21539
rect 16129 21505 16163 21539
rect 17417 21505 17451 21539
rect 17509 21505 17543 21539
rect 18245 21505 18279 21539
rect 23397 21505 23431 21539
rect 3525 21437 3559 21471
rect 5089 21437 5123 21471
rect 7665 21437 7699 21471
rect 9321 21437 9355 21471
rect 11621 21437 11655 21471
rect 12817 21437 12851 21471
rect 14381 21437 14415 21471
rect 15669 21437 15703 21471
rect 17601 21437 17635 21471
rect 20269 21437 20303 21471
rect 21005 21437 21039 21471
rect 22477 21437 22511 21471
rect 22569 21437 22603 21471
rect 23673 21437 23707 21471
rect 2329 21369 2363 21403
rect 13369 21369 13403 21403
rect 16313 21369 16347 21403
rect 16773 21369 16807 21403
rect 21557 21369 21591 21403
rect 2513 21301 2547 21335
rect 10793 21301 10827 21335
rect 11345 21301 11379 21335
rect 11805 21301 11839 21335
rect 12265 21301 12299 21335
rect 13553 21301 13587 21335
rect 15025 21301 15059 21335
rect 16405 21301 16439 21335
rect 17049 21301 17083 21335
rect 19533 21301 19567 21335
rect 23029 21301 23063 21335
rect 25145 21301 25179 21335
rect 25421 21301 25455 21335
rect 1593 21097 1627 21131
rect 9321 21097 9355 21131
rect 12909 21097 12943 21131
rect 13645 21097 13679 21131
rect 16681 21097 16715 21131
rect 17877 21097 17911 21131
rect 18981 21097 19015 21131
rect 21189 21097 21223 21131
rect 9965 21029 9999 21063
rect 15485 21029 15519 21063
rect 24593 21029 24627 21063
rect 2881 20961 2915 20995
rect 4445 20961 4479 20995
rect 7389 20961 7423 20995
rect 8769 20961 8803 20995
rect 10425 20961 10459 20995
rect 10517 20961 10551 20995
rect 11161 20961 11195 20995
rect 11437 20961 11471 20995
rect 16037 20961 16071 20995
rect 17233 20961 17267 20995
rect 18521 20961 18555 20995
rect 19717 20961 19751 20995
rect 22201 20961 22235 20995
rect 22753 20961 22787 20995
rect 23029 20961 23063 20995
rect 25053 20961 25087 20995
rect 25145 20961 25179 20995
rect 2237 20893 2271 20927
rect 4169 20893 4203 20927
rect 5825 20893 5859 20927
rect 7113 20893 7147 20927
rect 14381 20893 14415 20927
rect 18245 20893 18279 20927
rect 19441 20893 19475 20927
rect 23857 20893 23891 20927
rect 9229 20825 9263 20859
rect 13553 20825 13587 20859
rect 15945 20825 15979 20859
rect 17049 20825 17083 20859
rect 18337 20825 18371 20859
rect 22109 20825 22143 20859
rect 22845 20825 22879 20859
rect 23213 20825 23247 20859
rect 24501 20825 24535 20859
rect 24961 20825 24995 20859
rect 1777 20757 1811 20791
rect 6469 20757 6503 20791
rect 10333 20757 10367 20791
rect 15025 20757 15059 20791
rect 15853 20757 15887 20791
rect 17141 20757 17175 20791
rect 21649 20757 21683 20791
rect 22017 20757 22051 20791
rect 23489 20757 23523 20791
rect 23949 20757 23983 20791
rect 2237 20553 2271 20587
rect 6561 20553 6595 20587
rect 11529 20553 11563 20587
rect 11713 20553 11747 20587
rect 12449 20553 12483 20587
rect 13185 20553 13219 20587
rect 18705 20553 18739 20587
rect 21005 20553 21039 20587
rect 21281 20553 21315 20587
rect 21465 20553 21499 20587
rect 22477 20553 22511 20587
rect 1685 20485 1719 20519
rect 4813 20485 4847 20519
rect 8585 20485 8619 20519
rect 11161 20485 11195 20519
rect 13816 20485 13850 20519
rect 15577 20485 15611 20519
rect 23765 20485 23799 20519
rect 3065 20417 3099 20451
rect 6193 20417 6227 20451
rect 6837 20417 6871 20451
rect 7941 20417 7975 20451
rect 9045 20417 9079 20451
rect 11253 20417 11287 20451
rect 13553 20417 13587 20451
rect 16129 20417 16163 20451
rect 16957 20417 16991 20451
rect 23489 20417 23523 20451
rect 2605 20349 2639 20383
rect 3433 20349 3467 20383
rect 5549 20349 5583 20383
rect 9321 20349 9355 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 15301 20349 15335 20383
rect 17233 20349 17267 20383
rect 19257 20349 19291 20383
rect 19533 20349 19567 20383
rect 22569 20349 22603 20383
rect 22661 20349 22695 20383
rect 1869 20281 1903 20315
rect 23121 20281 23155 20315
rect 2421 20213 2455 20247
rect 4905 20213 4939 20247
rect 7481 20213 7515 20247
rect 10793 20213 10827 20247
rect 12081 20213 12115 20247
rect 16221 20213 16255 20247
rect 22109 20213 22143 20247
rect 25237 20213 25271 20247
rect 1501 20009 1535 20043
rect 1685 20009 1719 20043
rect 5273 20009 5307 20043
rect 6653 20009 6687 20043
rect 7297 20009 7331 20043
rect 9045 20009 9079 20043
rect 14933 20009 14967 20043
rect 17693 20009 17727 20043
rect 20545 20009 20579 20043
rect 21360 20009 21394 20043
rect 24593 20009 24627 20043
rect 13369 19941 13403 19975
rect 13921 19941 13955 19975
rect 3985 19873 4019 19907
rect 10977 19873 11011 19907
rect 15485 19873 15519 19907
rect 17141 19873 17175 19907
rect 18153 19873 18187 19907
rect 18337 19873 18371 19907
rect 19901 19873 19935 19907
rect 19993 19873 20027 19907
rect 20637 19873 20671 19907
rect 21097 19873 21131 19907
rect 23949 19873 23983 19907
rect 25053 19873 25087 19907
rect 25145 19873 25179 19907
rect 2237 19805 2271 19839
rect 4261 19805 4295 19839
rect 5457 19805 5491 19839
rect 6837 19805 6871 19839
rect 7481 19805 7515 19839
rect 7941 19805 7975 19839
rect 9321 19805 9355 19839
rect 10793 19805 10827 19839
rect 11621 19805 11655 19839
rect 13737 19805 13771 19839
rect 15393 19805 15427 19839
rect 16129 19805 16163 19839
rect 16773 19805 16807 19839
rect 18981 19805 19015 19839
rect 23765 19805 23799 19839
rect 2973 19737 3007 19771
rect 6009 19737 6043 19771
rect 10885 19737 10919 19771
rect 11897 19737 11931 19771
rect 8585 19669 8619 19703
rect 9965 19669 9999 19703
rect 10425 19669 10459 19703
rect 14289 19669 14323 19703
rect 15301 19669 15335 19703
rect 17417 19669 17451 19703
rect 18061 19669 18095 19703
rect 18797 19669 18831 19703
rect 19349 19669 19383 19703
rect 19441 19669 19475 19703
rect 19809 19669 19843 19703
rect 22845 19669 22879 19703
rect 23305 19669 23339 19703
rect 23673 19669 23707 19703
rect 24961 19669 24995 19703
rect 4537 19465 4571 19499
rect 6561 19465 6595 19499
rect 8585 19465 8619 19499
rect 10793 19465 10827 19499
rect 14473 19465 14507 19499
rect 14933 19465 14967 19499
rect 15301 19465 15335 19499
rect 18797 19465 18831 19499
rect 19257 19465 19291 19499
rect 19625 19465 19659 19499
rect 20453 19465 20487 19499
rect 20913 19465 20947 19499
rect 22017 19465 22051 19499
rect 25053 19465 25087 19499
rect 9321 19397 9355 19431
rect 15393 19397 15427 19431
rect 1961 19329 1995 19363
rect 4077 19329 4111 19363
rect 4721 19329 4755 19363
rect 5457 19329 5491 19363
rect 6745 19329 6779 19363
rect 7297 19329 7331 19363
rect 7941 19329 7975 19363
rect 9045 19329 9079 19363
rect 11161 19329 11195 19363
rect 11621 19329 11655 19363
rect 12265 19329 12299 19363
rect 12725 19329 12759 19363
rect 16129 19329 16163 19363
rect 17049 19329 17083 19363
rect 19717 19329 19751 19363
rect 20821 19329 20855 19363
rect 22385 19329 22419 19363
rect 23305 19329 23339 19363
rect 1501 19261 1535 19295
rect 2237 19261 2271 19295
rect 3525 19261 3559 19295
rect 5181 19261 5215 19295
rect 13001 19261 13035 19295
rect 15577 19261 15611 19295
rect 17325 19261 17359 19295
rect 19901 19261 19935 19295
rect 21005 19261 21039 19295
rect 21557 19261 21591 19295
rect 22477 19261 22511 19295
rect 22569 19261 22603 19295
rect 23581 19261 23615 19295
rect 3893 19193 3927 19227
rect 11345 19125 11379 19159
rect 11713 19125 11747 19159
rect 12081 19125 12115 19159
rect 16681 19125 16715 19159
rect 20269 19125 20303 19159
rect 21925 19125 21959 19159
rect 25329 19125 25363 19159
rect 1777 18921 1811 18955
rect 4077 18921 4111 18955
rect 14289 18921 14323 18955
rect 19625 18921 19659 18955
rect 4261 18853 4295 18887
rect 13001 18853 13035 18887
rect 17233 18853 17267 18887
rect 17601 18853 17635 18887
rect 18061 18853 18095 18887
rect 2881 18785 2915 18819
rect 3893 18785 3927 18819
rect 4813 18785 4847 18819
rect 6469 18785 6503 18819
rect 6745 18785 6779 18819
rect 9781 18785 9815 18819
rect 13645 18785 13679 18819
rect 14841 18785 14875 18819
rect 18521 18785 18555 18819
rect 18613 18785 18647 18819
rect 19993 18785 20027 18819
rect 20637 18785 20671 18819
rect 23121 18785 23155 18819
rect 24041 18785 24075 18819
rect 25237 18785 25271 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2605 18717 2639 18751
rect 4537 18717 4571 18751
rect 6009 18717 6043 18751
rect 7941 18717 7975 18751
rect 10425 18717 10459 18751
rect 12541 18717 12575 18751
rect 15485 18717 15519 18751
rect 20361 18717 20395 18751
rect 9597 18649 9631 18683
rect 9689 18649 9723 18683
rect 13369 18649 13403 18683
rect 14749 18649 14783 18683
rect 15761 18649 15795 18683
rect 19533 18649 19567 18683
rect 23029 18649 23063 18683
rect 23857 18649 23891 18683
rect 25053 18649 25087 18683
rect 5825 18581 5859 18615
rect 7757 18581 7791 18615
rect 8401 18581 8435 18615
rect 9229 18581 9263 18615
rect 11713 18581 11747 18615
rect 12633 18581 12667 18615
rect 13461 18581 13495 18615
rect 14657 18581 14691 18615
rect 17693 18581 17727 18615
rect 18429 18581 18463 18615
rect 22109 18581 22143 18615
rect 22569 18581 22603 18615
rect 22937 18581 22971 18615
rect 24409 18581 24443 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 1961 18377 1995 18411
rect 2605 18377 2639 18411
rect 3893 18377 3927 18411
rect 6377 18377 6411 18411
rect 6745 18377 6779 18411
rect 8309 18377 8343 18411
rect 12173 18377 12207 18411
rect 14289 18377 14323 18411
rect 15209 18377 15243 18411
rect 21557 18377 21591 18411
rect 23305 18377 23339 18411
rect 24961 18377 24995 18411
rect 9229 18309 9263 18343
rect 18521 18309 18555 18343
rect 22017 18309 22051 18343
rect 25053 18309 25087 18343
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 2789 18241 2823 18275
rect 3433 18241 3467 18275
rect 4077 18241 4111 18275
rect 6009 18241 6043 18275
rect 7205 18241 7239 18275
rect 7849 18241 7883 18275
rect 8493 18241 8527 18275
rect 8953 18241 8987 18275
rect 11069 18241 11103 18275
rect 13001 18241 13035 18275
rect 15577 18241 15611 18275
rect 15669 18241 15703 18275
rect 16405 18241 16439 18275
rect 17233 18241 17267 18275
rect 17325 18241 17359 18275
rect 18429 18241 18463 18275
rect 19625 18241 19659 18275
rect 20821 18241 20855 18275
rect 4537 18173 4571 18207
rect 4813 18173 4847 18207
rect 11253 18173 11287 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 15761 18173 15795 18207
rect 17417 18173 17451 18207
rect 18613 18173 18647 18207
rect 19717 18173 19751 18207
rect 19901 18173 19935 18207
rect 20913 18173 20947 18207
rect 21097 18173 21131 18207
rect 25237 18173 25271 18207
rect 7665 18105 7699 18139
rect 11805 18105 11839 18139
rect 16221 18105 16255 18139
rect 24593 18105 24627 18139
rect 3249 18037 3283 18071
rect 5825 18037 5859 18071
rect 7021 18037 7055 18071
rect 10701 18037 10735 18071
rect 16865 18037 16899 18071
rect 18061 18037 18095 18071
rect 19257 18037 19291 18071
rect 20453 18037 20487 18071
rect 24041 18037 24075 18071
rect 24225 18037 24259 18071
rect 3893 17833 3927 17867
rect 4261 17833 4295 17867
rect 6469 17833 6503 17867
rect 7757 17833 7791 17867
rect 17141 17833 17175 17867
rect 20992 17833 21026 17867
rect 22477 17833 22511 17867
rect 23305 17833 23339 17867
rect 24593 17833 24627 17867
rect 9137 17765 9171 17799
rect 18705 17765 18739 17799
rect 1961 17697 1995 17731
rect 5457 17697 5491 17731
rect 9781 17697 9815 17731
rect 11989 17697 12023 17731
rect 12265 17697 12299 17731
rect 14933 17697 14967 17731
rect 15209 17697 15243 17731
rect 17693 17697 17727 17731
rect 20085 17697 20119 17731
rect 20729 17697 20763 17731
rect 23029 17697 23063 17731
rect 23857 17697 23891 17731
rect 25237 17697 25271 17731
rect 2789 17629 2823 17663
rect 3433 17629 3467 17663
rect 4077 17629 4111 17663
rect 4721 17629 4755 17663
rect 5181 17629 5215 17663
rect 6653 17629 6687 17663
rect 7297 17629 7331 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9321 17629 9355 17663
rect 14473 17629 14507 17663
rect 19901 17629 19935 17663
rect 23673 17629 23707 17663
rect 23765 17629 23799 17663
rect 10057 17561 10091 17595
rect 17509 17561 17543 17595
rect 18521 17561 18555 17595
rect 18981 17561 19015 17595
rect 19809 17561 19843 17595
rect 25053 17561 25087 17595
rect 2605 17493 2639 17527
rect 3249 17493 3283 17527
rect 4537 17493 4571 17527
rect 7113 17493 7147 17527
rect 8401 17493 8435 17527
rect 11529 17493 11563 17527
rect 13737 17493 13771 17527
rect 14289 17493 14323 17527
rect 16681 17493 16715 17527
rect 17601 17493 17635 17527
rect 19441 17493 19475 17527
rect 22845 17493 22879 17527
rect 24409 17493 24443 17527
rect 24961 17493 24995 17527
rect 1593 17289 1627 17323
rect 2605 17289 2639 17323
rect 7205 17289 7239 17323
rect 7849 17289 7883 17323
rect 15853 17289 15887 17323
rect 17877 17289 17911 17323
rect 20085 17289 20119 17323
rect 22293 17289 22327 17323
rect 2329 17221 2363 17255
rect 9505 17221 9539 17255
rect 24869 17221 24903 17255
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2789 17153 2823 17187
rect 3249 17153 3283 17187
rect 3525 17153 3559 17187
rect 4813 17153 4847 17187
rect 6009 17153 6043 17187
rect 6745 17153 6779 17187
rect 7389 17153 7423 17187
rect 8033 17153 8067 17187
rect 8769 17153 8803 17187
rect 9229 17153 9263 17187
rect 11253 17153 11287 17187
rect 11713 17153 11747 17187
rect 14381 17153 14415 17187
rect 17233 17153 17267 17187
rect 17325 17153 17359 17187
rect 18337 17153 18371 17187
rect 20545 17153 20579 17187
rect 22569 17153 22603 17187
rect 25329 17153 25363 17187
rect 4537 17085 4571 17119
rect 10977 17085 11011 17119
rect 11989 17085 12023 17119
rect 13461 17085 13495 17119
rect 15945 17085 15979 17119
rect 16037 17085 16071 17119
rect 17417 17085 17451 17119
rect 18613 17085 18647 17119
rect 21189 17085 21223 17119
rect 21557 17085 21591 17119
rect 21925 17085 21959 17119
rect 22109 17085 22143 17119
rect 24317 17085 24351 17119
rect 5825 17017 5859 17051
rect 8585 17017 8619 17051
rect 15025 17017 15059 17051
rect 25053 17017 25087 17051
rect 6561 16949 6595 16983
rect 13737 16949 13771 16983
rect 14105 16949 14139 16983
rect 15485 16949 15519 16983
rect 16865 16949 16899 16983
rect 22832 16949 22866 16983
rect 5825 16745 5859 16779
rect 7297 16745 7331 16779
rect 7757 16745 7791 16779
rect 9045 16745 9079 16779
rect 9229 16745 9263 16779
rect 16037 16745 16071 16779
rect 19704 16745 19738 16779
rect 6561 16677 6595 16711
rect 8401 16677 8435 16711
rect 9505 16677 9539 16711
rect 10793 16677 10827 16711
rect 2513 16609 2547 16643
rect 3893 16609 3927 16643
rect 4537 16609 4571 16643
rect 4813 16609 4847 16643
rect 7113 16609 7147 16643
rect 10149 16609 10183 16643
rect 11253 16609 11287 16643
rect 11437 16609 11471 16643
rect 14289 16609 14323 16643
rect 17417 16609 17451 16643
rect 19441 16609 19475 16643
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 2789 16541 2823 16575
rect 3433 16541 3467 16575
rect 6009 16541 6043 16575
rect 6745 16541 6779 16575
rect 7481 16541 7515 16575
rect 7941 16541 7975 16575
rect 8585 16541 8619 16575
rect 9689 16541 9723 16575
rect 11161 16541 11195 16575
rect 11989 16541 12023 16575
rect 17141 16541 17175 16575
rect 21833 16541 21867 16575
rect 24593 16541 24627 16575
rect 25237 16541 25271 16575
rect 12265 16473 12299 16507
rect 14565 16473 14599 16507
rect 1961 16405 1995 16439
rect 2605 16405 2639 16439
rect 3249 16405 3283 16439
rect 13737 16405 13771 16439
rect 16497 16405 16531 16439
rect 18889 16405 18923 16439
rect 21189 16405 21223 16439
rect 21649 16405 21683 16439
rect 24041 16405 24075 16439
rect 3249 16201 3283 16235
rect 3893 16201 3927 16235
rect 4537 16201 4571 16235
rect 10793 16201 10827 16235
rect 10885 16201 10919 16235
rect 14381 16201 14415 16235
rect 19349 16201 19383 16235
rect 20913 16201 20947 16235
rect 22477 16201 22511 16235
rect 23397 16201 23431 16235
rect 23857 16201 23891 16235
rect 19717 16133 19751 16167
rect 19809 16133 19843 16167
rect 21557 16133 21591 16167
rect 2145 16065 2179 16099
rect 2789 16065 2823 16099
rect 4077 16065 4111 16099
rect 5457 16065 5491 16099
rect 8033 16065 8067 16099
rect 8677 16065 8711 16099
rect 9321 16065 9355 16099
rect 9965 16065 9999 16099
rect 14289 16065 14323 16099
rect 15025 16065 15059 16099
rect 15853 16065 15887 16099
rect 17141 16065 17175 16099
rect 22385 16065 22419 16099
rect 23121 16065 23155 16099
rect 23765 16065 23799 16099
rect 24593 16065 24627 16099
rect 5181 15997 5215 16031
rect 6561 15997 6595 16031
rect 6837 15997 6871 16031
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 14565 15997 14599 16031
rect 15945 15997 15979 16031
rect 16037 15997 16071 16031
rect 18889 15997 18923 16031
rect 19993 15997 20027 16031
rect 21005 15997 21039 16031
rect 21189 15997 21223 16031
rect 22569 15997 22603 16031
rect 23949 15997 23983 16031
rect 1961 15929 1995 15963
rect 7849 15929 7883 15963
rect 9781 15929 9815 15963
rect 13921 15929 13955 15963
rect 15485 15929 15519 15963
rect 20545 15929 20579 15963
rect 2605 15861 2639 15895
rect 8493 15861 8527 15895
rect 9137 15861 9171 15895
rect 10425 15861 10459 15895
rect 13461 15861 13495 15895
rect 15209 15861 15243 15895
rect 16681 15861 16715 15895
rect 22017 15861 22051 15895
rect 23305 15861 23339 15895
rect 25237 15861 25271 15895
rect 2237 15657 2271 15691
rect 3985 15657 4019 15691
rect 6561 15657 6595 15691
rect 7757 15657 7791 15691
rect 8033 15657 8067 15691
rect 8309 15657 8343 15691
rect 9229 15657 9263 15691
rect 18705 15657 18739 15691
rect 23949 15657 23983 15691
rect 7849 15589 7883 15623
rect 12725 15589 12759 15623
rect 16037 15589 16071 15623
rect 16405 15589 16439 15623
rect 16589 15589 16623 15623
rect 20729 15589 20763 15623
rect 24133 15589 24167 15623
rect 5365 15521 5399 15555
rect 8401 15521 8435 15555
rect 13185 15521 13219 15555
rect 13369 15521 13403 15555
rect 14289 15521 14323 15555
rect 16957 15521 16991 15555
rect 17233 15521 17267 15555
rect 20085 15521 20119 15555
rect 21189 15521 21223 15555
rect 21373 15521 21407 15555
rect 4169 15453 4203 15487
rect 4905 15453 4939 15487
rect 6745 15453 6779 15487
rect 7389 15453 7423 15487
rect 9413 15453 9447 15487
rect 10057 15453 10091 15487
rect 10517 15453 10551 15487
rect 13093 15453 13127 15487
rect 19993 15453 20027 15487
rect 21925 15453 21959 15487
rect 23029 15453 23063 15487
rect 24685 15453 24719 15487
rect 10793 15385 10827 15419
rect 14565 15385 14599 15419
rect 18981 15385 19015 15419
rect 4721 15317 4755 15351
rect 5917 15317 5951 15351
rect 7205 15317 7239 15351
rect 9873 15317 9907 15351
rect 12265 15317 12299 15351
rect 13921 15317 13955 15351
rect 19533 15317 19567 15351
rect 19901 15317 19935 15351
rect 21097 15317 21131 15351
rect 22569 15317 22603 15351
rect 23673 15317 23707 15351
rect 25329 15317 25363 15351
rect 4261 15113 4295 15147
rect 9413 15113 9447 15147
rect 10333 15113 10367 15147
rect 10977 15113 11011 15147
rect 21557 15113 21591 15147
rect 24593 15113 24627 15147
rect 6929 15045 6963 15079
rect 9689 15045 9723 15079
rect 11989 15045 12023 15079
rect 17141 15045 17175 15079
rect 22109 15045 22143 15079
rect 23121 15045 23155 15079
rect 25145 15045 25179 15079
rect 10517 14977 10551 15011
rect 11161 14977 11195 15011
rect 14105 14977 14139 15011
rect 15669 14977 15703 15011
rect 11713 14909 11747 14943
rect 13461 14909 13495 14943
rect 14657 14909 14691 14943
rect 15209 14909 15243 14943
rect 16865 14909 16899 14943
rect 18889 14909 18923 14943
rect 19349 14909 19383 14943
rect 19625 14909 19659 14943
rect 21097 14909 21131 14943
rect 22845 14909 22879 14943
rect 9597 14841 9631 14875
rect 16313 14841 16347 14875
rect 25329 14841 25363 14875
rect 13921 14773 13955 14807
rect 18613 14773 18647 14807
rect 21373 14773 21407 14807
rect 22201 14773 22235 14807
rect 10057 14569 10091 14603
rect 19441 14569 19475 14603
rect 20453 14569 20487 14603
rect 22293 14569 22327 14603
rect 18245 14501 18279 14535
rect 10977 14433 11011 14467
rect 12449 14433 12483 14467
rect 13553 14433 13587 14467
rect 14289 14433 14323 14467
rect 14565 14433 14599 14467
rect 16773 14433 16807 14467
rect 19993 14433 20027 14467
rect 23765 14433 23799 14467
rect 23949 14433 23983 14467
rect 10241 14365 10275 14399
rect 10701 14365 10735 14399
rect 16497 14365 16531 14399
rect 19809 14365 19843 14399
rect 20821 14365 20855 14399
rect 24593 14365 24627 14399
rect 22937 14297 22971 14331
rect 12909 14229 12943 14263
rect 16037 14229 16071 14263
rect 18705 14229 18739 14263
rect 19901 14229 19935 14263
rect 23305 14229 23339 14263
rect 23673 14229 23707 14263
rect 25237 14229 25271 14263
rect 10609 14025 10643 14059
rect 10977 14025 11011 14059
rect 11621 14025 11655 14059
rect 12265 14025 12299 14059
rect 12909 14025 12943 14059
rect 17049 14025 17083 14059
rect 17509 14025 17543 14059
rect 19533 14025 19567 14059
rect 20361 14025 20395 14059
rect 21833 14025 21867 14059
rect 22201 14025 22235 14059
rect 16129 13957 16163 13991
rect 18245 13957 18279 13991
rect 21189 13957 21223 13991
rect 22109 13957 22143 13991
rect 23121 13957 23155 13991
rect 11161 13889 11195 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 12449 13889 12483 13923
rect 13093 13889 13127 13923
rect 13737 13889 13771 13923
rect 16681 13889 16715 13923
rect 17417 13889 17451 13923
rect 21097 13889 21131 13923
rect 22845 13889 22879 13923
rect 25145 13889 25179 13923
rect 10425 13821 10459 13855
rect 15485 13821 15519 13855
rect 16313 13821 16347 13855
rect 17693 13821 17727 13855
rect 21281 13821 21315 13855
rect 24593 13821 24627 13855
rect 25329 13821 25363 13855
rect 13461 13753 13495 13787
rect 14000 13685 14034 13719
rect 20729 13685 20763 13719
rect 13921 13481 13955 13515
rect 16037 13481 16071 13515
rect 19980 13481 20014 13515
rect 21465 13481 21499 13515
rect 23673 13481 23707 13515
rect 14289 13345 14323 13379
rect 16497 13345 16531 13379
rect 16773 13345 16807 13379
rect 19717 13345 19751 13379
rect 25053 13345 25087 13379
rect 25145 13345 25179 13379
rect 11805 13277 11839 13311
rect 18705 13277 18739 13311
rect 21925 13277 21959 13311
rect 9597 13209 9631 13243
rect 12081 13209 12115 13243
rect 14565 13209 14599 13243
rect 19349 13209 19383 13243
rect 22201 13209 22235 13243
rect 24961 13209 24995 13243
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 18245 13141 18279 13175
rect 23949 13141 23983 13175
rect 24133 13141 24167 13175
rect 24593 13141 24627 13175
rect 11345 12937 11379 12971
rect 12725 12937 12759 12971
rect 14289 12937 14323 12971
rect 19533 12937 19567 12971
rect 20729 12937 20763 12971
rect 23765 12937 23799 12971
rect 25329 12937 25363 12971
rect 13001 12869 13035 12903
rect 15025 12869 15059 12903
rect 19441 12869 19475 12903
rect 22293 12869 22327 12903
rect 11989 12801 12023 12835
rect 12357 12801 12391 12835
rect 15485 12801 15519 12835
rect 16313 12801 16347 12835
rect 16865 12801 16899 12835
rect 20637 12801 20671 12835
rect 22017 12801 22051 12835
rect 24225 12801 24259 12835
rect 17141 12733 17175 12767
rect 19625 12733 19659 12767
rect 20821 12733 20855 12767
rect 16129 12665 16163 12699
rect 18613 12665 18647 12699
rect 24869 12665 24903 12699
rect 11805 12597 11839 12631
rect 19073 12597 19107 12631
rect 20269 12597 20303 12631
rect 21281 12597 21315 12631
rect 21465 12597 21499 12631
rect 25145 12597 25179 12631
rect 14197 12393 14231 12427
rect 17509 12393 17543 12427
rect 24041 12393 24075 12427
rect 17969 12325 18003 12359
rect 14749 12257 14783 12291
rect 15761 12257 15795 12291
rect 22293 12257 22327 12291
rect 22569 12257 22603 12291
rect 12909 12189 12943 12223
rect 13185 12189 13219 12223
rect 14473 12189 14507 12223
rect 18153 12189 18187 12223
rect 19441 12189 19475 12223
rect 21649 12189 21683 12223
rect 24593 12189 24627 12223
rect 16037 12121 16071 12155
rect 18705 12121 18739 12155
rect 18889 12121 18923 12155
rect 19717 12121 19751 12155
rect 21189 12053 21223 12087
rect 25237 12053 25271 12087
rect 14565 11849 14599 11883
rect 15117 11849 15151 11883
rect 15577 11849 15611 11883
rect 16681 11849 16715 11883
rect 13093 11781 13127 11815
rect 15853 11781 15887 11815
rect 19717 11781 19751 11815
rect 23305 11781 23339 11815
rect 25145 11781 25179 11815
rect 12817 11713 12851 11747
rect 15301 11713 15335 11747
rect 16313 11713 16347 11747
rect 17141 11713 17175 11747
rect 19441 11713 19475 11747
rect 22293 11713 22327 11747
rect 23949 11713 23983 11747
rect 17417 11645 17451 11679
rect 16129 11577 16163 11611
rect 18889 11509 18923 11543
rect 21189 11509 21223 11543
rect 21557 11509 21591 11543
rect 15485 11305 15519 11339
rect 16129 11305 16163 11339
rect 16773 11305 16807 11339
rect 17417 11305 17451 11339
rect 18705 11305 18739 11339
rect 22109 11237 22143 11271
rect 14841 11169 14875 11203
rect 18061 11169 18095 11203
rect 19901 11169 19935 11203
rect 23857 11169 23891 11203
rect 13553 11101 13587 11135
rect 15669 11101 15703 11135
rect 16313 11101 16347 11135
rect 16957 11101 16991 11135
rect 17601 11101 17635 11135
rect 18889 11101 18923 11135
rect 20177 11101 20211 11135
rect 20361 11101 20395 11135
rect 21465 11101 21499 11135
rect 22661 11101 22695 11135
rect 24593 11101 24627 11135
rect 19717 11033 19751 11067
rect 25237 11033 25271 11067
rect 19349 10965 19383 10999
rect 21005 10965 21039 10999
rect 15761 10761 15795 10795
rect 16681 10761 16715 10795
rect 16957 10761 16991 10795
rect 17325 10761 17359 10795
rect 17417 10761 17451 10795
rect 18705 10761 18739 10795
rect 19809 10761 19843 10795
rect 20085 10761 20119 10795
rect 20177 10761 20211 10795
rect 20545 10761 20579 10795
rect 23305 10693 23339 10727
rect 16313 10625 16347 10659
rect 17049 10625 17083 10659
rect 18889 10625 18923 10659
rect 19533 10625 19567 10659
rect 21281 10625 21315 10659
rect 22109 10625 22143 10659
rect 23949 10625 23983 10659
rect 18061 10557 18095 10591
rect 24777 10557 24811 10591
rect 16129 10489 16163 10523
rect 19349 10489 19383 10523
rect 21465 10489 21499 10523
rect 16773 10217 16807 10251
rect 16497 10149 16531 10183
rect 18061 10149 18095 10183
rect 24593 10149 24627 10183
rect 20729 10081 20763 10115
rect 21373 10081 21407 10115
rect 25145 10081 25179 10115
rect 16957 10013 16991 10047
rect 17601 10013 17635 10047
rect 18245 10013 18279 10047
rect 18889 10013 18923 10047
rect 19625 10013 19659 10047
rect 20269 10013 20303 10047
rect 25053 10013 25087 10047
rect 21649 9945 21683 9979
rect 23857 9945 23891 9979
rect 24041 9945 24075 9979
rect 17417 9877 17451 9911
rect 18705 9877 18739 9911
rect 19441 9877 19475 9911
rect 20085 9877 20119 9911
rect 23121 9877 23155 9911
rect 24961 9877 24995 9911
rect 23305 9605 23339 9639
rect 17049 9537 17083 9571
rect 17601 9537 17635 9571
rect 18245 9537 18279 9571
rect 18889 9537 18923 9571
rect 19625 9537 19659 9571
rect 20269 9537 20303 9571
rect 20637 9537 20671 9571
rect 20821 9537 20855 9571
rect 21005 9537 21039 9571
rect 21465 9537 21499 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 24685 9469 24719 9503
rect 17417 9401 17451 9435
rect 18705 9401 18739 9435
rect 19441 9401 19475 9435
rect 20085 9401 20119 9435
rect 18061 9333 18095 9367
rect 21281 9333 21315 9367
rect 11805 9129 11839 9163
rect 17693 9129 17727 9163
rect 19441 9129 19475 9163
rect 20913 9129 20947 9163
rect 21097 9129 21131 9163
rect 24593 9129 24627 9163
rect 25053 9129 25087 9163
rect 10057 8993 10091 9027
rect 18061 8993 18095 9027
rect 20085 8993 20119 9027
rect 21649 8993 21683 9027
rect 23857 8993 23891 9027
rect 18337 8925 18371 8959
rect 19625 8925 19659 8959
rect 20729 8925 20763 8959
rect 21373 8925 21407 8959
rect 22661 8925 22695 8959
rect 10333 8857 10367 8891
rect 12173 8857 12207 8891
rect 24501 8789 24535 8823
rect 24869 8789 24903 8823
rect 25237 8789 25271 8823
rect 25421 8789 25455 8823
rect 19441 8585 19475 8619
rect 19993 8517 20027 8551
rect 20177 8517 20211 8551
rect 21281 8517 21315 8551
rect 23305 8517 23339 8551
rect 18981 8449 19015 8483
rect 19625 8449 19659 8483
rect 20821 8449 20855 8483
rect 22109 8449 22143 8483
rect 23949 8449 23983 8483
rect 20361 8381 20395 8415
rect 24777 8381 24811 8415
rect 18797 8313 18831 8347
rect 20637 8313 20671 8347
rect 18705 8041 18739 8075
rect 19993 8041 20027 8075
rect 24685 8041 24719 8075
rect 19717 7973 19751 8007
rect 24501 7973 24535 8007
rect 23857 7905 23891 7939
rect 18889 7837 18923 7871
rect 20177 7837 20211 7871
rect 20913 7837 20947 7871
rect 21557 7837 21591 7871
rect 22201 7837 22235 7871
rect 22661 7837 22695 7871
rect 25145 7837 25179 7871
rect 25329 7769 25363 7803
rect 20729 7701 20763 7735
rect 21373 7701 21407 7735
rect 22017 7701 22051 7735
rect 19993 7497 20027 7531
rect 23305 7429 23339 7463
rect 25145 7429 25179 7463
rect 20177 7361 20211 7395
rect 20821 7361 20855 7395
rect 21465 7361 21499 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 20637 7225 20671 7259
rect 21281 7157 21315 7191
rect 20637 6953 20671 6987
rect 21281 6817 21315 6851
rect 21557 6817 21591 6851
rect 23857 6817 23891 6851
rect 25237 6817 25271 6851
rect 20177 6749 20211 6783
rect 20821 6749 20855 6783
rect 22661 6749 22695 6783
rect 24869 6749 24903 6783
rect 25421 6681 25455 6715
rect 19993 6613 20027 6647
rect 24685 6613 24719 6647
rect 9321 6409 9355 6443
rect 20361 6409 20395 6443
rect 21281 6409 21315 6443
rect 23305 6341 23339 6375
rect 8677 6273 8711 6307
rect 20821 6273 20855 6307
rect 22109 6273 22143 6307
rect 24133 6273 24167 6307
rect 24777 6205 24811 6239
rect 20637 6069 20671 6103
rect 20637 5865 20671 5899
rect 25329 5865 25363 5899
rect 21281 5797 21315 5831
rect 25237 5797 25271 5831
rect 22017 5729 22051 5763
rect 20821 5661 20855 5695
rect 21465 5661 21499 5695
rect 22845 5661 22879 5695
rect 23857 5661 23891 5695
rect 24685 5593 24719 5627
rect 24869 5593 24903 5627
rect 21281 5321 21315 5355
rect 23305 5253 23339 5287
rect 21465 5185 21499 5219
rect 22293 5185 22327 5219
rect 23949 5185 23983 5219
rect 24685 5117 24719 5151
rect 8585 4777 8619 4811
rect 25145 4777 25179 4811
rect 21373 4709 21407 4743
rect 24685 4709 24719 4743
rect 7941 4573 7975 4607
rect 21557 4573 21591 4607
rect 22845 4573 22879 4607
rect 24869 4573 24903 4607
rect 23857 4505 23891 4539
rect 22017 4437 22051 4471
rect 20269 4097 20303 4131
rect 22293 4097 22327 4131
rect 23949 4097 23983 4131
rect 21281 4029 21315 4063
rect 23305 4029 23339 4063
rect 24777 4029 24811 4063
rect 6837 3485 6871 3519
rect 20821 3485 20855 3519
rect 22845 3485 22879 3519
rect 24869 3485 24903 3519
rect 22017 3417 22051 3451
rect 23857 3417 23891 3451
rect 7481 3349 7515 3383
rect 24685 3349 24719 3383
rect 7481 3145 7515 3179
rect 23305 3077 23339 3111
rect 25145 3077 25179 3111
rect 6837 3009 6871 3043
rect 18429 3009 18463 3043
rect 20085 3009 20119 3043
rect 22293 3009 22327 3043
rect 24041 3009 24075 3043
rect 19349 2941 19383 2975
rect 21281 2941 21315 2975
rect 6561 2805 6595 2839
rect 6561 2601 6595 2635
rect 7849 2465 7883 2499
rect 21281 2465 21315 2499
rect 6745 2397 6779 2431
rect 7205 2397 7239 2431
rect 20269 2397 20303 2431
rect 22845 2397 22879 2431
rect 24777 2397 24811 2431
rect 23857 2329 23891 2363
rect 24593 2261 24627 2295
<< metal1 >>
rect 3050 26392 3056 26444
rect 3108 26432 3114 26444
rect 3418 26432 3424 26444
rect 3108 26404 3424 26432
rect 3108 26392 3114 26404
rect 3418 26392 3424 26404
rect 3476 26392 3482 26444
rect 1946 26324 1952 26376
rect 2004 26364 2010 26376
rect 18690 26364 18696 26376
rect 2004 26336 18696 26364
rect 2004 26324 2010 26336
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 12802 24964 12808 25016
rect 12860 25004 12866 25016
rect 14918 25004 14924 25016
rect 12860 24976 14924 25004
rect 12860 24964 12866 24976
rect 14918 24964 14924 24976
rect 14976 24964 14982 25016
rect 15470 24964 15476 25016
rect 15528 25004 15534 25016
rect 20070 25004 20076 25016
rect 15528 24976 20076 25004
rect 15528 24964 15534 24976
rect 20070 24964 20076 24976
rect 20128 24964 20134 25016
rect 11606 24896 11612 24948
rect 11664 24936 11670 24948
rect 13078 24936 13084 24948
rect 11664 24908 13084 24936
rect 11664 24896 11670 24908
rect 13078 24896 13084 24908
rect 13136 24896 13142 24948
rect 16206 24896 16212 24948
rect 16264 24936 16270 24948
rect 18230 24936 18236 24948
rect 16264 24908 18236 24936
rect 16264 24896 16270 24908
rect 18230 24896 18236 24908
rect 18288 24896 18294 24948
rect 3694 24828 3700 24880
rect 3752 24868 3758 24880
rect 18414 24868 18420 24880
rect 3752 24840 18420 24868
rect 3752 24828 3758 24840
rect 18414 24828 18420 24840
rect 18472 24828 18478 24880
rect 11882 24760 11888 24812
rect 11940 24800 11946 24812
rect 12066 24800 12072 24812
rect 11940 24772 12072 24800
rect 11940 24760 11946 24772
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 13538 24760 13544 24812
rect 13596 24800 13602 24812
rect 18598 24800 18604 24812
rect 13596 24772 18604 24800
rect 13596 24760 13602 24772
rect 18598 24760 18604 24772
rect 18656 24760 18662 24812
rect 7466 24692 7472 24744
rect 7524 24732 7530 24744
rect 20530 24732 20536 24744
rect 7524 24704 20536 24732
rect 7524 24692 7530 24704
rect 20530 24692 20536 24704
rect 20588 24692 20594 24744
rect 4154 24624 4160 24676
rect 4212 24664 4218 24676
rect 13722 24664 13728 24676
rect 4212 24636 13728 24664
rect 4212 24624 4218 24636
rect 13722 24624 13728 24636
rect 13780 24624 13786 24676
rect 15010 24624 15016 24676
rect 15068 24664 15074 24676
rect 21450 24664 21456 24676
rect 15068 24636 21456 24664
rect 15068 24624 15074 24636
rect 21450 24624 21456 24636
rect 21508 24624 21514 24676
rect 5810 24556 5816 24608
rect 5868 24596 5874 24608
rect 12250 24596 12256 24608
rect 5868 24568 12256 24596
rect 5868 24556 5874 24568
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 14090 24556 14096 24608
rect 14148 24596 14154 24608
rect 17218 24596 17224 24608
rect 14148 24568 17224 24596
rect 14148 24556 14154 24568
rect 17218 24556 17224 24568
rect 17276 24556 17282 24608
rect 17586 24556 17592 24608
rect 17644 24596 17650 24608
rect 24118 24596 24124 24608
rect 17644 24568 24124 24596
rect 17644 24556 17650 24568
rect 24118 24556 24124 24568
rect 24176 24556 24182 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 1581 24395 1639 24401
rect 1581 24361 1593 24395
rect 1627 24392 1639 24395
rect 6730 24392 6736 24404
rect 1627 24364 6736 24392
rect 1627 24361 1639 24364
rect 1581 24355 1639 24361
rect 6730 24352 6736 24364
rect 6788 24352 6794 24404
rect 11790 24392 11796 24404
rect 6840 24364 11796 24392
rect 4706 24324 4712 24336
rect 2746 24296 4712 24324
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2746 24188 2774 24296
rect 4706 24284 4712 24296
rect 4764 24284 4770 24336
rect 5350 24284 5356 24336
rect 5408 24324 5414 24336
rect 6840 24324 6868 24364
rect 11790 24352 11796 24364
rect 11848 24352 11854 24404
rect 14090 24392 14096 24404
rect 11900 24364 14096 24392
rect 5408 24296 6868 24324
rect 5408 24284 5414 24296
rect 9766 24284 9772 24336
rect 9824 24324 9830 24336
rect 11701 24327 11759 24333
rect 11701 24324 11713 24327
rect 9824 24296 11713 24324
rect 9824 24284 9830 24296
rect 11701 24293 11713 24296
rect 11747 24293 11759 24327
rect 11701 24287 11759 24293
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 6454 24256 6460 24268
rect 3283 24228 6460 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 8205 24259 8263 24265
rect 6564 24228 7236 24256
rect 2271 24160 2774 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 4154 24148 4160 24200
rect 4212 24148 4218 24200
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 5258 24148 5264 24200
rect 5316 24188 5322 24200
rect 6564 24188 6592 24228
rect 5316 24160 6592 24188
rect 5316 24148 5322 24160
rect 6730 24148 6736 24200
rect 6788 24148 6794 24200
rect 7208 24197 7236 24228
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9674 24256 9680 24268
rect 8251 24228 9680 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 11238 24256 11244 24268
rect 11011 24228 11244 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 7742 24148 7748 24200
rect 7800 24188 7806 24200
rect 11900 24197 11928 24364
rect 14090 24352 14096 24364
rect 14148 24352 14154 24404
rect 14369 24395 14427 24401
rect 14369 24361 14381 24395
rect 14415 24392 14427 24395
rect 16850 24392 16856 24404
rect 14415 24364 16856 24392
rect 14415 24361 14427 24364
rect 14369 24355 14427 24361
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 16942 24352 16948 24404
rect 17000 24352 17006 24404
rect 19886 24392 19892 24404
rect 17420 24364 19892 24392
rect 13630 24284 13636 24336
rect 13688 24324 13694 24336
rect 15470 24324 15476 24336
rect 13688 24296 15476 24324
rect 13688 24284 13694 24296
rect 15470 24284 15476 24296
rect 15528 24284 15534 24336
rect 15562 24284 15568 24336
rect 15620 24284 15626 24336
rect 12342 24216 12348 24268
rect 12400 24256 12406 24268
rect 12805 24259 12863 24265
rect 12805 24256 12817 24259
rect 12400 24228 12817 24256
rect 12400 24216 12406 24228
rect 12805 24225 12817 24228
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 13998 24216 14004 24268
rect 14056 24256 14062 24268
rect 14550 24256 14556 24268
rect 14056 24228 14556 24256
rect 14056 24216 14062 24228
rect 14550 24216 14556 24228
rect 14608 24216 14614 24268
rect 15013 24259 15071 24265
rect 15013 24225 15025 24259
rect 15059 24256 15071 24259
rect 15059 24228 16160 24256
rect 15059 24225 15071 24228
rect 15013 24219 15071 24225
rect 9769 24191 9827 24197
rect 9769 24188 9781 24191
rect 7800 24160 9781 24188
rect 7800 24148 7806 24160
rect 9769 24157 9781 24160
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 12434 24148 12440 24200
rect 12492 24148 12498 24200
rect 16132 24188 16160 24228
rect 16206 24216 16212 24268
rect 16264 24216 16270 24268
rect 17420 24265 17448 24364
rect 19886 24352 19892 24364
rect 19944 24392 19950 24404
rect 21821 24395 21879 24401
rect 21821 24392 21833 24395
rect 19944 24364 21833 24392
rect 19944 24352 19950 24364
rect 21821 24361 21833 24364
rect 21867 24361 21879 24395
rect 23750 24392 23756 24404
rect 21821 24355 21879 24361
rect 22066 24364 23756 24392
rect 18141 24327 18199 24333
rect 18141 24293 18153 24327
rect 18187 24293 18199 24327
rect 18141 24287 18199 24293
rect 17405 24259 17463 24265
rect 17405 24225 17417 24259
rect 17451 24225 17463 24259
rect 17405 24219 17463 24225
rect 17497 24259 17555 24265
rect 17497 24225 17509 24259
rect 17543 24225 17555 24259
rect 17497 24219 17555 24225
rect 16482 24188 16488 24200
rect 16132 24160 16488 24188
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 17512 24188 17540 24219
rect 17954 24216 17960 24268
rect 18012 24256 18018 24268
rect 18156 24256 18184 24287
rect 18230 24284 18236 24336
rect 18288 24324 18294 24336
rect 22066 24324 22094 24364
rect 23750 24352 23756 24364
rect 23808 24352 23814 24404
rect 18288 24296 22094 24324
rect 18288 24284 18294 24296
rect 18012 24228 18184 24256
rect 18012 24216 18018 24228
rect 18322 24216 18328 24268
rect 18380 24256 18386 24268
rect 18693 24259 18751 24265
rect 18693 24256 18705 24259
rect 18380 24228 18705 24256
rect 18380 24216 18386 24228
rect 18693 24225 18705 24228
rect 18739 24225 18751 24259
rect 22646 24256 22652 24268
rect 18693 24219 18751 24225
rect 20088 24228 22652 24256
rect 17512 24160 17724 24188
rect 1673 24123 1731 24129
rect 1673 24089 1685 24123
rect 1719 24120 1731 24123
rect 5626 24120 5632 24132
rect 1719 24092 5632 24120
rect 1719 24089 1731 24092
rect 1673 24083 1731 24089
rect 5626 24080 5632 24092
rect 5684 24080 5690 24132
rect 5813 24123 5871 24129
rect 5813 24089 5825 24123
rect 5859 24120 5871 24123
rect 8386 24120 8392 24132
rect 5859 24092 8392 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 8386 24080 8392 24092
rect 8444 24080 8450 24132
rect 8570 24080 8576 24132
rect 8628 24120 8634 24132
rect 12158 24120 12164 24132
rect 8628 24092 12164 24120
rect 8628 24080 8634 24092
rect 12158 24080 12164 24092
rect 12216 24080 12222 24132
rect 12250 24080 12256 24132
rect 12308 24120 12314 24132
rect 13814 24120 13820 24132
rect 12308 24092 13820 24120
rect 12308 24080 12314 24092
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 16025 24123 16083 24129
rect 16025 24120 16037 24123
rect 14200 24092 16037 24120
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 4982 24052 4988 24064
rect 4019 24024 4988 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 4982 24012 4988 24024
rect 5040 24012 5046 24064
rect 6546 24012 6552 24064
rect 6604 24012 6610 24064
rect 9125 24055 9183 24061
rect 9125 24021 9137 24055
rect 9171 24052 9183 24055
rect 10962 24052 10968 24064
rect 9171 24024 10968 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 10962 24012 10968 24024
rect 11020 24012 11026 24064
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 14200 24052 14228 24092
rect 16025 24089 16037 24092
rect 16071 24089 16083 24123
rect 17696 24120 17724 24160
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 20088 24188 20116 24228
rect 22646 24216 22652 24228
rect 22704 24216 22710 24268
rect 25222 24216 25228 24268
rect 25280 24216 25286 24268
rect 18647 24160 20116 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 20162 24148 20168 24200
rect 20220 24148 20226 24200
rect 20530 24148 20536 24200
rect 20588 24148 20594 24200
rect 21450 24148 21456 24200
rect 21508 24148 21514 24200
rect 22278 24148 22284 24200
rect 22336 24148 22342 24200
rect 24949 24191 25007 24197
rect 24949 24157 24961 24191
rect 24995 24188 25007 24191
rect 25038 24188 25044 24200
rect 24995 24160 25044 24188
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 25038 24148 25044 24160
rect 25096 24148 25102 24200
rect 22462 24120 22468 24132
rect 16025 24083 16083 24089
rect 16132 24092 17448 24120
rect 17696 24092 22468 24120
rect 11848 24024 14228 24052
rect 11848 24012 11854 24024
rect 14734 24012 14740 24064
rect 14792 24012 14798 24064
rect 14826 24012 14832 24064
rect 14884 24012 14890 24064
rect 15562 24012 15568 24064
rect 15620 24052 15626 24064
rect 15933 24055 15991 24061
rect 15933 24052 15945 24055
rect 15620 24024 15945 24052
rect 15620 24012 15626 24024
rect 15933 24021 15945 24024
rect 15979 24052 15991 24055
rect 16132 24052 16160 24092
rect 15979 24024 16160 24052
rect 15979 24021 15991 24024
rect 15933 24015 15991 24021
rect 17310 24012 17316 24064
rect 17368 24012 17374 24064
rect 17420 24052 17448 24092
rect 22462 24080 22468 24092
rect 22520 24080 22526 24132
rect 22557 24123 22615 24129
rect 22557 24089 22569 24123
rect 22603 24089 22615 24123
rect 22557 24083 22615 24089
rect 18690 24052 18696 24064
rect 17420 24024 18696 24052
rect 18690 24012 18696 24024
rect 18748 24012 18754 24064
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 19518 24052 19524 24064
rect 19475 24024 19524 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 19518 24012 19524 24024
rect 19576 24012 19582 24064
rect 21266 24012 21272 24064
rect 21324 24012 21330 24064
rect 22572 24052 22600 24083
rect 23014 24080 23020 24132
rect 23072 24080 23078 24132
rect 23842 24052 23848 24064
rect 22572 24024 23848 24052
rect 23842 24012 23848 24024
rect 23900 24012 23906 24064
rect 24029 24055 24087 24061
rect 24029 24021 24041 24055
rect 24075 24052 24087 24055
rect 24118 24052 24124 24064
rect 24075 24024 24124 24052
rect 24075 24021 24087 24024
rect 24029 24015 24087 24021
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24578 24012 24584 24064
rect 24636 24012 24642 24064
rect 24670 24012 24676 24064
rect 24728 24052 24734 24064
rect 25041 24055 25099 24061
rect 25041 24052 25053 24055
rect 24728 24024 25053 24052
rect 24728 24012 24734 24024
rect 25041 24021 25053 24024
rect 25087 24021 25099 24055
rect 25041 24015 25099 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 3786 23808 3792 23860
rect 3844 23848 3850 23860
rect 3844 23820 9812 23848
rect 3844 23808 3850 23820
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 5166 23780 5172 23792
rect 4019 23752 5172 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 5166 23740 5172 23752
rect 5224 23740 5230 23792
rect 5813 23783 5871 23789
rect 5813 23749 5825 23783
rect 5859 23780 5871 23783
rect 7374 23780 7380 23792
rect 5859 23752 7380 23780
rect 5859 23749 5871 23752
rect 5813 23743 5871 23749
rect 7374 23740 7380 23752
rect 7432 23740 7438 23792
rect 9125 23783 9183 23789
rect 7484 23752 8064 23780
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 1854 23712 1860 23724
rect 1719 23684 1860 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 4154 23712 4160 23724
rect 3007 23684 4160 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 4154 23672 4160 23684
rect 4212 23672 4218 23724
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23681 4859 23715
rect 4801 23675 4859 23681
rect 4816 23644 4844 23675
rect 5626 23672 5632 23724
rect 5684 23712 5690 23724
rect 6825 23715 6883 23721
rect 6825 23712 6837 23715
rect 5684 23684 6837 23712
rect 5684 23672 5690 23684
rect 6825 23681 6837 23684
rect 6871 23712 6883 23715
rect 7484 23712 7512 23752
rect 6871 23684 7512 23712
rect 6871 23681 6883 23684
rect 6825 23675 6883 23681
rect 7558 23672 7564 23724
rect 7616 23712 7622 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7616 23684 7941 23712
rect 7616 23672 7622 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 8036 23712 8064 23752
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9171 23752 9536 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 8036 23684 9444 23712
rect 7929 23675 7987 23681
rect 9306 23644 9312 23656
rect 4816 23616 9312 23644
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 5166 23536 5172 23588
rect 5224 23576 5230 23588
rect 7469 23579 7527 23585
rect 7469 23576 7481 23579
rect 5224 23548 7481 23576
rect 5224 23536 5230 23548
rect 7469 23545 7481 23548
rect 7515 23545 7527 23579
rect 9416 23576 9444 23684
rect 9508 23644 9536 23752
rect 9784 23721 9812 23820
rect 10686 23808 10692 23860
rect 10744 23848 10750 23860
rect 16669 23851 16727 23857
rect 16669 23848 16681 23851
rect 10744 23820 16681 23848
rect 10744 23808 10750 23820
rect 16669 23817 16681 23820
rect 16715 23817 16727 23851
rect 16669 23811 16727 23817
rect 16853 23851 16911 23857
rect 16853 23817 16865 23851
rect 16899 23848 16911 23851
rect 24670 23848 24676 23860
rect 16899 23820 24676 23848
rect 16899 23817 16911 23820
rect 16853 23811 16911 23817
rect 10870 23740 10876 23792
rect 10928 23740 10934 23792
rect 14734 23780 14740 23792
rect 11716 23752 14740 23780
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 10134 23644 10140 23656
rect 9508 23616 10140 23644
rect 10134 23604 10140 23616
rect 10192 23604 10198 23656
rect 11422 23604 11428 23656
rect 11480 23644 11486 23656
rect 11716 23653 11744 23752
rect 14734 23740 14740 23752
rect 14792 23740 14798 23792
rect 15562 23740 15568 23792
rect 15620 23780 15626 23792
rect 15933 23783 15991 23789
rect 15933 23780 15945 23783
rect 15620 23752 15945 23780
rect 15620 23740 15626 23752
rect 15933 23749 15945 23752
rect 15979 23749 15991 23783
rect 15933 23743 15991 23749
rect 16025 23783 16083 23789
rect 16025 23749 16037 23783
rect 16071 23780 16083 23783
rect 16114 23780 16120 23792
rect 16071 23752 16120 23780
rect 16071 23749 16083 23752
rect 16025 23743 16083 23749
rect 16114 23740 16120 23752
rect 16172 23740 16178 23792
rect 16684 23780 16712 23811
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 17313 23783 17371 23789
rect 17313 23780 17325 23783
rect 16684 23752 17325 23780
rect 17313 23749 17325 23752
rect 17359 23749 17371 23783
rect 20073 23783 20131 23789
rect 20073 23780 20085 23783
rect 19550 23752 20085 23780
rect 17313 23743 17371 23749
rect 20073 23749 20085 23752
rect 20119 23780 20131 23783
rect 20254 23780 20260 23792
rect 20119 23752 20260 23780
rect 20119 23749 20131 23752
rect 20073 23743 20131 23749
rect 20254 23740 20260 23752
rect 20312 23780 20318 23792
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 20312 23752 21833 23780
rect 20312 23740 20318 23752
rect 21821 23749 21833 23752
rect 21867 23780 21879 23783
rect 23014 23780 23020 23792
rect 21867 23752 23020 23780
rect 21867 23749 21879 23752
rect 21821 23743 21879 23749
rect 11882 23672 11888 23724
rect 11940 23712 11946 23724
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 11940 23684 12081 23712
rect 11940 23672 11946 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12069 23675 12127 23681
rect 12158 23672 12164 23724
rect 12216 23712 12222 23724
rect 13909 23715 13967 23721
rect 13909 23712 13921 23715
rect 12216 23684 13921 23712
rect 12216 23672 12222 23684
rect 13909 23681 13921 23684
rect 13955 23712 13967 23715
rect 14461 23715 14519 23721
rect 14461 23712 14473 23715
rect 13955 23684 14473 23712
rect 13955 23681 13967 23684
rect 13909 23675 13967 23681
rect 14461 23681 14473 23684
rect 14507 23681 14519 23715
rect 14461 23675 14519 23681
rect 14553 23715 14611 23721
rect 14553 23681 14565 23715
rect 14599 23712 14611 23715
rect 14599 23684 15884 23712
rect 14599 23681 14611 23684
rect 14553 23675 14611 23681
rect 11701 23647 11759 23653
rect 11701 23644 11713 23647
rect 11480 23616 11713 23644
rect 11480 23604 11486 23616
rect 11701 23613 11713 23616
rect 11747 23613 11759 23647
rect 11701 23607 11759 23613
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12032 23616 12541 23644
rect 12032 23604 12038 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 13872 23616 14136 23644
rect 13872 23604 13878 23616
rect 13630 23576 13636 23588
rect 9416 23548 13636 23576
rect 7469 23539 7527 23545
rect 13630 23536 13636 23548
rect 13688 23536 13694 23588
rect 14108 23585 14136 23616
rect 14734 23604 14740 23656
rect 14792 23604 14798 23656
rect 15856 23644 15884 23684
rect 16040 23684 16988 23712
rect 16040 23644 16068 23684
rect 15856 23616 16068 23644
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 16960 23644 16988 23684
rect 17034 23672 17040 23724
rect 17092 23712 17098 23724
rect 17221 23715 17279 23721
rect 17221 23712 17233 23715
rect 17092 23684 17233 23712
rect 17092 23672 17098 23684
rect 17221 23681 17233 23684
rect 17267 23681 17279 23715
rect 17221 23675 17279 23681
rect 17420 23684 18000 23712
rect 17420 23644 17448 23684
rect 16255 23616 16896 23644
rect 16960 23616 17448 23644
rect 17497 23647 17555 23653
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 14093 23579 14151 23585
rect 14093 23545 14105 23579
rect 14139 23545 14151 23579
rect 14093 23539 14151 23545
rect 2222 23468 2228 23520
rect 2280 23508 2286 23520
rect 2317 23511 2375 23517
rect 2317 23508 2329 23511
rect 2280 23480 2329 23508
rect 2280 23468 2286 23480
rect 2317 23477 2329 23480
rect 2363 23477 2375 23511
rect 2317 23471 2375 23477
rect 6549 23511 6607 23517
rect 6549 23477 6561 23511
rect 6595 23508 6607 23511
rect 6914 23508 6920 23520
rect 6595 23480 6920 23508
rect 6595 23477 6607 23480
rect 6549 23471 6607 23477
rect 6914 23468 6920 23480
rect 6972 23468 6978 23520
rect 11609 23511 11667 23517
rect 11609 23477 11621 23511
rect 11655 23508 11667 23511
rect 11790 23508 11796 23520
rect 11655 23480 11796 23508
rect 11655 23477 11667 23480
rect 11609 23471 11667 23477
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 11974 23468 11980 23520
rect 12032 23508 12038 23520
rect 12434 23508 12440 23520
rect 12032 23480 12440 23508
rect 12032 23468 12038 23480
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 13817 23511 13875 23517
rect 13817 23477 13829 23511
rect 13863 23508 13875 23511
rect 14918 23508 14924 23520
rect 13863 23480 14924 23508
rect 13863 23477 13875 23480
rect 13817 23471 13875 23477
rect 14918 23468 14924 23480
rect 14976 23468 14982 23520
rect 15197 23511 15255 23517
rect 15197 23477 15209 23511
rect 15243 23508 15255 23511
rect 15378 23508 15384 23520
rect 15243 23480 15384 23508
rect 15243 23477 15255 23480
rect 15197 23471 15255 23477
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 15565 23511 15623 23517
rect 15565 23477 15577 23511
rect 15611 23508 15623 23511
rect 16390 23508 16396 23520
rect 15611 23480 16396 23508
rect 15611 23477 15623 23480
rect 15565 23471 15623 23477
rect 16390 23468 16396 23480
rect 16448 23468 16454 23520
rect 16868 23508 16896 23616
rect 17497 23613 17509 23647
rect 17543 23644 17555 23647
rect 17586 23644 17592 23656
rect 17543 23616 17592 23644
rect 17543 23613 17555 23616
rect 17497 23607 17555 23613
rect 17586 23604 17592 23616
rect 17644 23604 17650 23656
rect 17862 23508 17868 23520
rect 16868 23480 17868 23508
rect 17862 23468 17868 23480
rect 17920 23468 17926 23520
rect 17972 23508 18000 23684
rect 20622 23672 20628 23724
rect 20680 23672 20686 23724
rect 18046 23604 18052 23656
rect 18104 23604 18110 23656
rect 18322 23604 18328 23656
rect 18380 23604 18386 23656
rect 18690 23604 18696 23656
rect 18748 23644 18754 23656
rect 20901 23647 20959 23653
rect 20901 23644 20913 23647
rect 18748 23616 20913 23644
rect 18748 23604 18754 23616
rect 20901 23613 20913 23616
rect 20947 23644 20959 23647
rect 21818 23644 21824 23656
rect 20947 23616 21824 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 21818 23604 21824 23616
rect 21876 23604 21882 23656
rect 22204 23588 22232 23752
rect 23014 23740 23020 23752
rect 23072 23740 23078 23792
rect 24026 23740 24032 23792
rect 24084 23780 24090 23792
rect 24394 23780 24400 23792
rect 24084 23752 24400 23780
rect 24084 23740 24090 23752
rect 24394 23740 24400 23752
rect 24452 23780 24458 23792
rect 24581 23783 24639 23789
rect 24581 23780 24593 23783
rect 24452 23752 24593 23780
rect 24452 23740 24458 23752
rect 24581 23749 24593 23752
rect 24627 23749 24639 23783
rect 24581 23743 24639 23749
rect 25130 23740 25136 23792
rect 25188 23780 25194 23792
rect 25774 23780 25780 23792
rect 25188 23752 25780 23780
rect 25188 23740 25194 23752
rect 25774 23740 25780 23752
rect 25832 23740 25838 23792
rect 23842 23672 23848 23724
rect 23900 23712 23906 23724
rect 25314 23712 25320 23724
rect 23900 23684 25320 23712
rect 23900 23672 23906 23684
rect 22278 23604 22284 23656
rect 22336 23604 22342 23656
rect 22554 23604 22560 23656
rect 22612 23604 22618 23656
rect 24044 23653 24072 23684
rect 25314 23672 25320 23684
rect 25372 23672 25378 23724
rect 24029 23647 24087 23653
rect 24029 23613 24041 23647
rect 24075 23613 24087 23647
rect 24029 23607 24087 23613
rect 20349 23579 20407 23585
rect 20349 23576 20361 23579
rect 19352 23548 20361 23576
rect 18506 23508 18512 23520
rect 17972 23480 18512 23508
rect 18506 23468 18512 23480
rect 18564 23468 18570 23520
rect 18782 23468 18788 23520
rect 18840 23508 18846 23520
rect 19352 23508 19380 23548
rect 20349 23545 20361 23548
rect 20395 23545 20407 23579
rect 20349 23539 20407 23545
rect 21910 23536 21916 23588
rect 21968 23576 21974 23588
rect 21968 23548 22094 23576
rect 21968 23536 21974 23548
rect 18840 23480 19380 23508
rect 18840 23468 18846 23480
rect 19794 23468 19800 23520
rect 19852 23468 19858 23520
rect 22066 23508 22094 23548
rect 22186 23536 22192 23588
rect 22244 23536 22250 23588
rect 25317 23579 25375 23585
rect 25317 23576 25329 23579
rect 23584 23548 25329 23576
rect 23584 23508 23612 23548
rect 25317 23545 25329 23548
rect 25363 23545 25375 23579
rect 25317 23539 25375 23545
rect 22066 23480 23612 23508
rect 24394 23468 24400 23520
rect 24452 23468 24458 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 1762 23264 1768 23316
rect 1820 23264 1826 23316
rect 9306 23264 9312 23316
rect 9364 23264 9370 23316
rect 11330 23264 11336 23316
rect 11388 23304 11394 23316
rect 13354 23304 13360 23316
rect 11388 23276 13360 23304
rect 11388 23264 11394 23276
rect 13354 23264 13360 23276
rect 13412 23264 13418 23316
rect 14182 23304 14188 23316
rect 13464 23276 14188 23304
rect 8478 23196 8484 23248
rect 8536 23236 8542 23248
rect 8536 23208 10640 23236
rect 8536 23196 8542 23208
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 4249 23171 4307 23177
rect 1627 23140 4200 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 2314 23100 2320 23112
rect 2271 23072 2320 23100
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 3970 23060 3976 23112
rect 4028 23060 4034 23112
rect 4172 23100 4200 23140
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 4295 23140 9996 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 5442 23100 5448 23112
rect 4172 23072 5448 23100
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 5552 23072 7205 23100
rect 3237 23035 3295 23041
rect 3237 23001 3249 23035
rect 3283 23032 3295 23035
rect 4614 23032 4620 23044
rect 3283 23004 4620 23032
rect 3283 23001 3295 23004
rect 3237 22995 3295 23001
rect 4614 22992 4620 23004
rect 4672 22992 4678 23044
rect 4890 22992 4896 23044
rect 4948 23032 4954 23044
rect 5552 23032 5580 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23100 8263 23103
rect 9398 23100 9404 23112
rect 8251 23072 9404 23100
rect 8251 23069 8263 23072
rect 8205 23063 8263 23069
rect 9398 23060 9404 23072
rect 9456 23060 9462 23112
rect 9490 23060 9496 23112
rect 9548 23100 9554 23112
rect 9861 23103 9919 23109
rect 9861 23100 9873 23103
rect 9548 23072 9873 23100
rect 9548 23060 9554 23072
rect 9861 23069 9873 23072
rect 9907 23069 9919 23103
rect 9968 23100 9996 23140
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 10612 23168 10640 23208
rect 11054 23196 11060 23248
rect 11112 23236 11118 23248
rect 13464 23236 13492 23276
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 14918 23264 14924 23316
rect 14976 23304 14982 23316
rect 16298 23304 16304 23316
rect 14976 23276 16304 23304
rect 14976 23264 14982 23276
rect 16298 23264 16304 23276
rect 16356 23264 16362 23316
rect 16942 23264 16948 23316
rect 17000 23304 17006 23316
rect 18046 23304 18052 23316
rect 17000 23276 18052 23304
rect 17000 23264 17006 23276
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 18322 23264 18328 23316
rect 18380 23304 18386 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 18380 23276 21189 23304
rect 18380 23264 18386 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 21266 23264 21272 23316
rect 21324 23304 21330 23316
rect 22370 23304 22376 23316
rect 21324 23276 22376 23304
rect 21324 23264 21330 23276
rect 22370 23264 22376 23276
rect 22428 23264 22434 23316
rect 22554 23264 22560 23316
rect 22612 23304 22618 23316
rect 23385 23307 23443 23313
rect 23385 23304 23397 23307
rect 22612 23276 23397 23304
rect 22612 23264 22618 23276
rect 23385 23273 23397 23276
rect 23431 23273 23443 23307
rect 23385 23267 23443 23273
rect 24302 23264 24308 23316
rect 24360 23304 24366 23316
rect 24397 23307 24455 23313
rect 24397 23304 24409 23307
rect 24360 23276 24409 23304
rect 24360 23264 24366 23276
rect 24397 23273 24409 23276
rect 24443 23304 24455 23307
rect 24443 23276 25084 23304
rect 24443 23273 24455 23276
rect 24397 23267 24455 23273
rect 11112 23208 13492 23236
rect 13541 23239 13599 23245
rect 11112 23196 11118 23208
rect 13541 23205 13553 23239
rect 13587 23236 13599 23239
rect 14642 23236 14648 23248
rect 13587 23208 14648 23236
rect 13587 23205 13599 23208
rect 13541 23199 13599 23205
rect 14642 23196 14648 23208
rect 14700 23196 14706 23248
rect 16758 23196 16764 23248
rect 16816 23236 16822 23248
rect 18690 23236 18696 23248
rect 16816 23208 18696 23236
rect 16816 23196 16822 23208
rect 18690 23196 18696 23208
rect 18748 23196 18754 23248
rect 23934 23196 23940 23248
rect 23992 23236 23998 23248
rect 24581 23239 24639 23245
rect 24581 23236 24593 23239
rect 23992 23208 24593 23236
rect 23992 23196 23998 23208
rect 24581 23205 24593 23208
rect 24627 23205 24639 23239
rect 24581 23199 24639 23205
rect 10612 23140 11836 23168
rect 11701 23103 11759 23109
rect 11701 23100 11713 23103
rect 9968 23072 11713 23100
rect 9861 23063 9919 23069
rect 11701 23069 11713 23072
rect 11747 23069 11759 23103
rect 11808 23100 11836 23140
rect 12066 23128 12072 23180
rect 12124 23168 12130 23180
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 12124 23140 12173 23168
rect 12124 23128 12130 23140
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 13906 23168 13912 23180
rect 12161 23131 12219 23137
rect 12268 23140 13912 23168
rect 12268 23100 12296 23140
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 17770 23168 17776 23180
rect 15335 23140 17776 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18966 23168 18972 23180
rect 18012 23140 18972 23168
rect 18012 23128 18018 23140
rect 18966 23128 18972 23140
rect 19024 23128 19030 23180
rect 19242 23128 19248 23180
rect 19300 23168 19306 23180
rect 19705 23171 19763 23177
rect 19300 23140 19472 23168
rect 19300 23128 19334 23140
rect 13725 23103 13783 23109
rect 13725 23100 13737 23103
rect 11808 23072 12296 23100
rect 12406 23072 13737 23100
rect 11701 23063 11759 23069
rect 4948 23004 5580 23032
rect 6549 23035 6607 23041
rect 4948 22992 4954 23004
rect 6549 23001 6561 23035
rect 6595 23032 6607 23035
rect 7650 23032 7656 23044
rect 6595 23004 7656 23032
rect 6595 23001 6607 23004
rect 6549 22995 6607 23001
rect 7650 22992 7656 23004
rect 7708 22992 7714 23044
rect 8386 22992 8392 23044
rect 8444 23032 8450 23044
rect 9217 23035 9275 23041
rect 9217 23032 9229 23035
rect 8444 23004 9229 23032
rect 8444 22992 8450 23004
rect 9217 23001 9229 23004
rect 9263 23001 9275 23035
rect 9217 22995 9275 23001
rect 9306 22992 9312 23044
rect 9364 23032 9370 23044
rect 12406 23032 12434 23072
rect 13725 23069 13737 23072
rect 13771 23069 13783 23103
rect 13725 23063 13783 23069
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 14240 23072 15025 23100
rect 14240 23060 14246 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 16666 23100 16672 23112
rect 16422 23072 16672 23100
rect 15013 23063 15071 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17589 23103 17647 23109
rect 17589 23100 17601 23103
rect 16908 23072 17601 23100
rect 16908 23060 16914 23072
rect 17589 23069 17601 23072
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 18046 23060 18052 23112
rect 18104 23100 18110 23112
rect 19306 23100 19334 23128
rect 19444 23109 19472 23140
rect 19705 23137 19717 23171
rect 19751 23168 19763 23171
rect 21174 23168 21180 23180
rect 19751 23140 21180 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 21174 23128 21180 23140
rect 21232 23128 21238 23180
rect 21637 23171 21695 23177
rect 21637 23137 21649 23171
rect 21683 23168 21695 23171
rect 22278 23168 22284 23180
rect 21683 23140 22284 23168
rect 21683 23137 21695 23140
rect 21637 23131 21695 23137
rect 22278 23128 22284 23140
rect 22336 23168 22342 23180
rect 23290 23168 23296 23180
rect 22336 23140 23296 23168
rect 22336 23128 22342 23140
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 25056 23177 25084 23276
rect 25041 23171 25099 23177
rect 25041 23137 25053 23171
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 18104 23072 19334 23100
rect 19429 23103 19487 23109
rect 18104 23060 18110 23072
rect 19429 23069 19441 23103
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23100 24087 23103
rect 25498 23100 25504 23112
rect 24075 23072 25504 23100
rect 24075 23069 24087 23072
rect 24029 23063 24087 23069
rect 25498 23060 25504 23072
rect 25556 23060 25562 23112
rect 14369 23035 14427 23041
rect 9364 23004 12434 23032
rect 13464 23004 13676 23032
rect 9364 22992 9370 23004
rect 9398 22924 9404 22976
rect 9456 22964 9462 22976
rect 13464 22964 13492 23004
rect 9456 22936 13492 22964
rect 13648 22964 13676 23004
rect 14369 23001 14381 23035
rect 14415 23032 14427 23035
rect 17126 23032 17132 23044
rect 14415 23004 14964 23032
rect 14415 23001 14427 23004
rect 14369 22995 14427 23001
rect 14461 22967 14519 22973
rect 14461 22964 14473 22967
rect 13648 22936 14473 22964
rect 9456 22924 9462 22936
rect 14461 22933 14473 22936
rect 14507 22933 14519 22967
rect 14936 22964 14964 23004
rect 16592 23004 17132 23032
rect 15378 22964 15384 22976
rect 14936 22936 15384 22964
rect 14461 22927 14519 22933
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 15470 22924 15476 22976
rect 15528 22964 15534 22976
rect 16592 22964 16620 23004
rect 17126 22992 17132 23004
rect 17184 22992 17190 23044
rect 18322 22992 18328 23044
rect 18380 23032 18386 23044
rect 18509 23035 18567 23041
rect 18509 23032 18521 23035
rect 18380 23004 18521 23032
rect 18380 22992 18386 23004
rect 18509 23001 18521 23004
rect 18555 23032 18567 23035
rect 18782 23032 18788 23044
rect 18555 23004 18788 23032
rect 18555 23001 18567 23004
rect 18509 22995 18567 23001
rect 18782 22992 18788 23004
rect 18840 22992 18846 23044
rect 18984 23004 19334 23032
rect 15528 22936 16620 22964
rect 15528 22924 15534 22936
rect 16758 22924 16764 22976
rect 16816 22924 16822 22976
rect 17221 22967 17279 22973
rect 17221 22933 17233 22967
rect 17267 22964 17279 22967
rect 17402 22964 17408 22976
rect 17267 22936 17408 22964
rect 17267 22933 17279 22936
rect 17221 22927 17279 22933
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 17678 22924 17684 22976
rect 17736 22924 17742 22976
rect 18414 22924 18420 22976
rect 18472 22964 18478 22976
rect 18601 22967 18659 22973
rect 18601 22964 18613 22967
rect 18472 22936 18613 22964
rect 18472 22924 18478 22936
rect 18601 22933 18613 22936
rect 18647 22933 18659 22967
rect 18601 22927 18659 22933
rect 18690 22924 18696 22976
rect 18748 22964 18754 22976
rect 18984 22964 19012 23004
rect 18748 22936 19012 22964
rect 19061 22967 19119 22973
rect 18748 22924 18754 22936
rect 19061 22933 19073 22967
rect 19107 22964 19119 22967
rect 19150 22964 19156 22976
rect 19107 22936 19156 22964
rect 19107 22933 19119 22936
rect 19061 22927 19119 22933
rect 19150 22924 19156 22936
rect 19208 22924 19214 22976
rect 19306 22964 19334 23004
rect 20254 22992 20260 23044
rect 20312 22992 20318 23044
rect 21634 22992 21640 23044
rect 21692 23032 21698 23044
rect 21913 23035 21971 23041
rect 21913 23032 21925 23035
rect 21692 23004 21925 23032
rect 21692 22992 21698 23004
rect 21913 23001 21925 23004
rect 21959 23001 21971 23035
rect 21913 22995 21971 23001
rect 22186 22992 22192 23044
rect 22244 23032 22250 23044
rect 22244 23004 22402 23032
rect 22244 22992 22250 23004
rect 23658 22992 23664 23044
rect 23716 23032 23722 23044
rect 24949 23035 25007 23041
rect 24949 23032 24961 23035
rect 23716 23004 24961 23032
rect 23716 22992 23722 23004
rect 24949 23001 24961 23004
rect 24995 23001 25007 23035
rect 24949 22995 25007 23001
rect 20990 22964 20996 22976
rect 19306 22936 20996 22964
rect 20990 22924 20996 22936
rect 21048 22924 21054 22976
rect 22922 22924 22928 22976
rect 22980 22964 22986 22976
rect 23845 22967 23903 22973
rect 23845 22964 23857 22967
rect 22980 22936 23857 22964
rect 22980 22924 22986 22936
rect 23845 22933 23857 22936
rect 23891 22933 23903 22967
rect 23845 22927 23903 22933
rect 24118 22924 24124 22976
rect 24176 22964 24182 22976
rect 24302 22964 24308 22976
rect 24176 22936 24308 22964
rect 24176 22924 24182 22936
rect 24302 22924 24308 22936
rect 24360 22964 24366 22976
rect 25590 22964 25596 22976
rect 24360 22936 25596 22964
rect 24360 22924 24366 22936
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 9398 22760 9404 22772
rect 4816 22732 9404 22760
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 4246 22692 4252 22704
rect 4019 22664 4252 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 1394 22584 1400 22636
rect 1452 22624 1458 22636
rect 1673 22627 1731 22633
rect 1673 22624 1685 22627
rect 1452 22596 1685 22624
rect 1452 22584 1458 22596
rect 1673 22593 1685 22596
rect 1719 22624 1731 22627
rect 1946 22624 1952 22636
rect 1719 22596 1952 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 1946 22584 1952 22596
rect 2004 22584 2010 22636
rect 2774 22584 2780 22636
rect 2832 22584 2838 22636
rect 4816 22633 4844 22732
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 12342 22760 12348 22772
rect 9508 22732 12348 22760
rect 5718 22652 5724 22704
rect 5776 22652 5782 22704
rect 6914 22652 6920 22704
rect 6972 22692 6978 22704
rect 7098 22692 7104 22704
rect 6972 22664 7104 22692
rect 6972 22652 6978 22664
rect 7098 22652 7104 22664
rect 7156 22652 7162 22704
rect 8754 22652 8760 22704
rect 8812 22652 8818 22704
rect 9508 22692 9536 22732
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 14734 22720 14740 22772
rect 14792 22760 14798 22772
rect 15381 22763 15439 22769
rect 15381 22760 15393 22763
rect 14792 22732 15393 22760
rect 14792 22720 14798 22732
rect 15381 22729 15393 22732
rect 15427 22729 15439 22763
rect 15381 22723 15439 22729
rect 16298 22720 16304 22772
rect 16356 22760 16362 22772
rect 16666 22760 16672 22772
rect 16356 22732 16672 22760
rect 16356 22720 16362 22732
rect 16666 22720 16672 22732
rect 16724 22760 16730 22772
rect 19245 22763 19303 22769
rect 16724 22732 18460 22760
rect 16724 22720 16730 22732
rect 11698 22692 11704 22704
rect 8864 22664 9536 22692
rect 10902 22664 11704 22692
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 4154 22516 4160 22568
rect 4212 22556 4218 22568
rect 7101 22559 7159 22565
rect 7101 22556 7113 22559
rect 4212 22528 7113 22556
rect 4212 22516 4218 22528
rect 7101 22525 7113 22528
rect 7147 22525 7159 22559
rect 7101 22519 7159 22525
rect 4614 22448 4620 22500
rect 4672 22488 4678 22500
rect 7576 22488 7604 22587
rect 7650 22584 7656 22636
rect 7708 22624 7714 22636
rect 8864 22624 8892 22664
rect 11698 22652 11704 22664
rect 11756 22652 11762 22704
rect 12069 22695 12127 22701
rect 12069 22661 12081 22695
rect 12115 22692 12127 22695
rect 12158 22692 12164 22704
rect 12115 22664 12164 22692
rect 12115 22661 12127 22664
rect 12069 22655 12127 22661
rect 12158 22652 12164 22664
rect 12216 22652 12222 22704
rect 13538 22692 13544 22704
rect 12636 22664 13544 22692
rect 12636 22624 12664 22664
rect 13538 22652 13544 22664
rect 13596 22652 13602 22704
rect 14182 22692 14188 22704
rect 13648 22664 14188 22692
rect 7708 22596 8892 22624
rect 11992 22596 12296 22624
rect 7708 22584 7714 22596
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 9088 22528 9413 22556
rect 9088 22516 9094 22528
rect 9401 22525 9413 22528
rect 9447 22525 9459 22559
rect 9401 22519 9459 22525
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 11992 22556 12020 22596
rect 12268 22568 12296 22596
rect 12360 22596 12664 22624
rect 12989 22627 13047 22633
rect 9723 22528 12020 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 12066 22516 12072 22568
rect 12124 22556 12130 22568
rect 12161 22559 12219 22565
rect 12161 22556 12173 22559
rect 12124 22528 12173 22556
rect 12124 22516 12130 22528
rect 12161 22525 12173 22528
rect 12207 22525 12219 22559
rect 12161 22519 12219 22525
rect 12250 22516 12256 22568
rect 12308 22516 12314 22568
rect 11701 22491 11759 22497
rect 11701 22488 11713 22491
rect 4672 22460 7604 22488
rect 10704 22460 11713 22488
rect 4672 22448 4678 22460
rect 2317 22423 2375 22429
rect 2317 22389 2329 22423
rect 2363 22420 2375 22423
rect 2682 22420 2688 22432
rect 2363 22392 2688 22420
rect 2363 22389 2375 22392
rect 2317 22383 2375 22389
rect 2682 22380 2688 22392
rect 2740 22380 2746 22432
rect 5994 22380 6000 22432
rect 6052 22420 6058 22432
rect 6457 22423 6515 22429
rect 6457 22420 6469 22423
rect 6052 22392 6469 22420
rect 6052 22380 6058 22392
rect 6457 22389 6469 22392
rect 6503 22420 6515 22423
rect 9398 22420 9404 22432
rect 6503 22392 9404 22420
rect 6503 22389 6515 22392
rect 6457 22383 6515 22389
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 10704 22420 10732 22460
rect 11701 22457 11713 22460
rect 11747 22457 11759 22491
rect 11701 22451 11759 22457
rect 9732 22392 10732 22420
rect 11149 22423 11207 22429
rect 9732 22380 9738 22392
rect 11149 22389 11161 22423
rect 11195 22420 11207 22423
rect 11238 22420 11244 22432
rect 11195 22392 11244 22420
rect 11195 22389 11207 22392
rect 11149 22383 11207 22389
rect 11238 22380 11244 22392
rect 11296 22380 11302 22432
rect 11514 22380 11520 22432
rect 11572 22420 11578 22432
rect 12360 22420 12388 22596
rect 12989 22593 13001 22627
rect 13035 22624 13047 22627
rect 13354 22624 13360 22636
rect 13035 22596 13360 22624
rect 13035 22593 13047 22596
rect 12989 22587 13047 22593
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 13648 22633 13676 22664
rect 14182 22652 14188 22664
rect 14240 22652 14246 22704
rect 14918 22652 14924 22704
rect 14976 22652 14982 22704
rect 15654 22652 15660 22704
rect 15712 22692 15718 22704
rect 16482 22692 16488 22704
rect 15712 22664 16488 22692
rect 15712 22652 15718 22664
rect 16482 22652 16488 22664
rect 16540 22692 16546 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16540 22664 17141 22692
rect 16540 22652 16546 22664
rect 17129 22661 17141 22664
rect 17175 22692 17187 22695
rect 17218 22692 17224 22704
rect 17175 22664 17224 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 17218 22652 17224 22664
rect 17276 22652 17282 22704
rect 18432 22692 18460 22732
rect 19245 22729 19257 22763
rect 19291 22760 19303 22763
rect 19610 22760 19616 22772
rect 19291 22732 19616 22760
rect 19291 22729 19303 22732
rect 19245 22723 19303 22729
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 20254 22720 20260 22772
rect 20312 22760 20318 22772
rect 21082 22760 21088 22772
rect 20312 22732 21088 22760
rect 20312 22720 20318 22732
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 21634 22720 21640 22772
rect 21692 22760 21698 22772
rect 22370 22760 22376 22772
rect 21692 22732 22376 22760
rect 21692 22720 21698 22732
rect 22370 22720 22376 22732
rect 22428 22720 22434 22772
rect 24302 22760 24308 22772
rect 23584 22732 24308 22760
rect 18598 22692 18604 22704
rect 18354 22664 18604 22692
rect 18598 22652 18604 22664
rect 18656 22652 18662 22704
rect 19153 22695 19211 22701
rect 19153 22661 19165 22695
rect 19199 22692 19211 22695
rect 22922 22692 22928 22704
rect 19199 22664 22928 22692
rect 19199 22661 19211 22664
rect 19153 22655 19211 22661
rect 22922 22652 22928 22664
rect 22980 22652 22986 22704
rect 23584 22701 23612 22732
rect 24302 22720 24308 22732
rect 24360 22720 24366 22772
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 25041 22763 25099 22769
rect 25041 22760 25053 22763
rect 24912 22732 25053 22760
rect 24912 22720 24918 22732
rect 25041 22729 25053 22732
rect 25087 22760 25099 22763
rect 25222 22760 25228 22772
rect 25087 22732 25228 22760
rect 25087 22729 25099 22732
rect 25041 22723 25099 22729
rect 25222 22720 25228 22732
rect 25280 22720 25286 22772
rect 23569 22695 23627 22701
rect 23569 22661 23581 22695
rect 23615 22661 23627 22695
rect 23569 22655 23627 22661
rect 23842 22652 23848 22704
rect 23900 22692 23906 22704
rect 23900 22664 24058 22692
rect 23900 22652 23906 22664
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22624 15991 22627
rect 16758 22624 16764 22636
rect 15979 22596 16764 22624
rect 15979 22593 15991 22596
rect 15933 22587 15991 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 16850 22584 16856 22636
rect 16908 22584 16914 22636
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 19484 22596 20177 22624
rect 19484 22584 19490 22596
rect 20165 22593 20177 22596
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22624 20775 22627
rect 22646 22624 22652 22636
rect 20763 22596 22652 22624
rect 20763 22593 20775 22596
rect 20717 22587 20775 22593
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 13909 22559 13967 22565
rect 13909 22525 13921 22559
rect 13955 22556 13967 22559
rect 14550 22556 14556 22568
rect 13955 22528 14556 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 14550 22516 14556 22528
rect 14608 22516 14614 22568
rect 14642 22516 14648 22568
rect 14700 22556 14706 22568
rect 14700 22528 16896 22556
rect 14700 22516 14706 22528
rect 16868 22500 16896 22528
rect 17770 22516 17776 22568
rect 17828 22556 17834 22568
rect 18601 22559 18659 22565
rect 18601 22556 18613 22559
rect 17828 22528 18613 22556
rect 17828 22516 17834 22528
rect 18601 22525 18613 22528
rect 18647 22525 18659 22559
rect 18601 22519 18659 22525
rect 19610 22516 19616 22568
rect 19668 22556 19674 22568
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 19668 22528 21281 22556
rect 19668 22516 19674 22528
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 21358 22516 21364 22568
rect 21416 22556 21422 22568
rect 22005 22559 22063 22565
rect 22005 22556 22017 22559
rect 21416 22528 22017 22556
rect 21416 22516 21422 22528
rect 22005 22525 22017 22528
rect 22051 22556 22063 22559
rect 22051 22528 22140 22556
rect 22051 22525 22063 22528
rect 22005 22519 22063 22525
rect 14918 22448 14924 22500
rect 14976 22488 14982 22500
rect 16117 22491 16175 22497
rect 16117 22488 16129 22491
rect 14976 22460 16129 22488
rect 14976 22448 14982 22460
rect 16117 22457 16129 22460
rect 16163 22457 16175 22491
rect 16117 22451 16175 22457
rect 16482 22448 16488 22500
rect 16540 22448 16546 22500
rect 16850 22448 16856 22500
rect 16908 22448 16914 22500
rect 19702 22488 19708 22500
rect 19306 22460 19708 22488
rect 11572 22392 12388 22420
rect 11572 22380 11578 22392
rect 12710 22380 12716 22432
rect 12768 22420 12774 22432
rect 13081 22423 13139 22429
rect 13081 22420 13093 22423
rect 12768 22392 13093 22420
rect 12768 22380 12774 22392
rect 13081 22389 13093 22392
rect 13127 22389 13139 22423
rect 13081 22383 13139 22389
rect 13538 22380 13544 22432
rect 13596 22420 13602 22432
rect 17126 22420 17132 22432
rect 13596 22392 17132 22420
rect 13596 22380 13602 22392
rect 17126 22380 17132 22392
rect 17184 22380 17190 22432
rect 17586 22380 17592 22432
rect 17644 22420 17650 22432
rect 19306 22420 19334 22460
rect 19702 22448 19708 22460
rect 19760 22448 19766 22500
rect 22112 22488 22140 22528
rect 22278 22516 22284 22568
rect 22336 22516 22342 22568
rect 23290 22516 23296 22568
rect 23348 22516 23354 22568
rect 24946 22556 24952 22568
rect 23400 22528 24952 22556
rect 23400 22488 23428 22528
rect 24946 22516 24952 22528
rect 25004 22516 25010 22568
rect 22112 22460 23428 22488
rect 25222 22448 25228 22500
rect 25280 22488 25286 22500
rect 25317 22491 25375 22497
rect 25317 22488 25329 22491
rect 25280 22460 25329 22488
rect 25280 22448 25286 22460
rect 25317 22457 25329 22460
rect 25363 22457 25375 22491
rect 25317 22451 25375 22457
rect 17644 22392 19334 22420
rect 17644 22380 17650 22392
rect 19426 22380 19432 22432
rect 19484 22420 19490 22432
rect 19613 22423 19671 22429
rect 19613 22420 19625 22423
rect 19484 22392 19625 22420
rect 19484 22380 19490 22392
rect 19613 22389 19625 22392
rect 19659 22389 19671 22423
rect 19613 22383 19671 22389
rect 21450 22380 21456 22432
rect 21508 22380 21514 22432
rect 22830 22380 22836 22432
rect 22888 22420 22894 22432
rect 25406 22420 25412 22432
rect 22888 22392 25412 22420
rect 22888 22380 22894 22392
rect 25406 22380 25412 22392
rect 25464 22380 25470 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 2406 22176 2412 22228
rect 2464 22216 2470 22228
rect 2958 22216 2964 22228
rect 2464 22188 2964 22216
rect 2464 22176 2470 22188
rect 2958 22176 2964 22188
rect 3016 22176 3022 22228
rect 10952 22219 11010 22225
rect 10952 22185 10964 22219
rect 10998 22216 11010 22219
rect 13538 22216 13544 22228
rect 10998 22188 13544 22216
rect 10998 22185 11010 22188
rect 10952 22179 11010 22185
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 14540 22219 14598 22225
rect 14540 22185 14552 22219
rect 14586 22216 14598 22219
rect 14734 22216 14740 22228
rect 14586 22188 14740 22216
rect 14586 22185 14598 22188
rect 14540 22179 14598 22185
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 14918 22176 14924 22228
rect 14976 22216 14982 22228
rect 16206 22216 16212 22228
rect 14976 22188 16212 22216
rect 14976 22176 14982 22188
rect 16206 22176 16212 22188
rect 16264 22176 16270 22228
rect 16485 22219 16543 22225
rect 16485 22216 16497 22219
rect 16408 22188 16497 22216
rect 2314 22108 2320 22160
rect 2372 22148 2378 22160
rect 9766 22148 9772 22160
rect 2372 22120 9772 22148
rect 2372 22108 2378 22120
rect 9766 22108 9772 22120
rect 9824 22108 9830 22160
rect 12066 22108 12072 22160
rect 12124 22148 12130 22160
rect 12124 22120 12572 22148
rect 12124 22108 12130 22120
rect 2866 22040 2872 22092
rect 2924 22040 2930 22092
rect 3878 22040 3884 22092
rect 3936 22080 3942 22092
rect 3973 22083 4031 22089
rect 3973 22080 3985 22083
rect 3936 22052 3985 22080
rect 3936 22040 3942 22052
rect 3973 22049 3985 22052
rect 4019 22080 4031 22083
rect 4019 22052 5672 22080
rect 4019 22049 4031 22052
rect 3973 22043 4031 22049
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 1762 21904 1768 21956
rect 1820 21904 1826 21956
rect 2240 21944 2268 21975
rect 4246 21972 4252 22024
rect 4304 21972 4310 22024
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 4522 21944 4528 21956
rect 2240 21916 4528 21944
rect 4522 21904 4528 21916
rect 4580 21904 4586 21956
rect 5552 21888 5580 21975
rect 5644 21944 5672 22052
rect 6086 22040 6092 22092
rect 6144 22040 6150 22092
rect 8294 22040 8300 22092
rect 8352 22040 8358 22092
rect 9030 22040 9036 22092
rect 9088 22080 9094 22092
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 9088 22052 10701 22080
rect 9088 22040 9094 22052
rect 10689 22049 10701 22052
rect 10735 22080 10747 22083
rect 11054 22080 11060 22092
rect 10735 22052 11060 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12437 22083 12495 22089
rect 12437 22080 12449 22083
rect 12308 22052 12449 22080
rect 12308 22040 12314 22052
rect 12437 22049 12449 22052
rect 12483 22049 12495 22083
rect 12544 22080 12572 22120
rect 12710 22108 12716 22160
rect 12768 22148 12774 22160
rect 13906 22148 13912 22160
rect 12768 22120 13912 22148
rect 12768 22108 12774 22120
rect 13906 22108 13912 22120
rect 13964 22108 13970 22160
rect 14200 22120 14412 22148
rect 14200 22080 14228 22120
rect 12544 22052 14228 22080
rect 14384 22080 14412 22120
rect 16408 22080 16436 22188
rect 16485 22185 16497 22188
rect 16531 22185 16543 22219
rect 16485 22179 16543 22185
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 17276 22188 18552 22216
rect 17276 22176 17282 22188
rect 18524 22148 18552 22188
rect 18598 22176 18604 22228
rect 18656 22216 18662 22228
rect 18693 22219 18751 22225
rect 18693 22216 18705 22219
rect 18656 22188 18705 22216
rect 18656 22176 18662 22188
rect 18693 22185 18705 22188
rect 18739 22185 18751 22219
rect 18693 22179 18751 22185
rect 18966 22176 18972 22228
rect 19024 22216 19030 22228
rect 20438 22216 20444 22228
rect 19024 22188 20444 22216
rect 19024 22176 19030 22188
rect 20438 22176 20444 22188
rect 20496 22216 20502 22228
rect 20606 22219 20664 22225
rect 20606 22216 20618 22219
rect 20496 22188 20618 22216
rect 20496 22176 20502 22188
rect 20606 22185 20618 22188
rect 20652 22185 20664 22219
rect 20606 22179 20664 22185
rect 21174 22176 21180 22228
rect 21232 22216 21238 22228
rect 21232 22188 25176 22216
rect 21232 22176 21238 22188
rect 19794 22148 19800 22160
rect 14384 22052 16436 22080
rect 16500 22120 18276 22148
rect 18524 22120 19800 22148
rect 12437 22043 12495 22049
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7834 22012 7840 22024
rect 7423 21984 7840 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 9596 22015 9654 22021
rect 9596 21981 9608 22015
rect 9642 21981 9654 22015
rect 12894 22012 12900 22024
rect 12098 21984 12900 22012
rect 9596 21975 9654 21981
rect 9398 21944 9404 21956
rect 5644 21916 9404 21944
rect 9398 21904 9404 21916
rect 9456 21904 9462 21956
rect 9600 21944 9628 21975
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 13078 21972 13084 22024
rect 13136 22012 13142 22024
rect 13630 22012 13636 22024
rect 13136 21984 13636 22012
rect 13136 21972 13142 21984
rect 13630 21972 13636 21984
rect 13688 21972 13694 22024
rect 14182 21972 14188 22024
rect 14240 22012 14246 22024
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 14240 21984 14289 22012
rect 14240 21972 14246 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 9766 21944 9772 21956
rect 9600 21916 9772 21944
rect 9766 21904 9772 21916
rect 9824 21904 9830 21956
rect 12728 21916 13124 21944
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 1946 21876 1952 21888
rect 1627 21848 1952 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 1946 21836 1952 21848
rect 2004 21836 2010 21888
rect 4430 21836 4436 21888
rect 4488 21876 4494 21888
rect 4893 21879 4951 21885
rect 4893 21876 4905 21879
rect 4488 21848 4905 21876
rect 4488 21836 4494 21848
rect 4893 21845 4905 21848
rect 4939 21845 4951 21879
rect 4893 21839 4951 21845
rect 5534 21836 5540 21888
rect 5592 21836 5598 21888
rect 6730 21836 6736 21888
rect 6788 21876 6794 21888
rect 8386 21876 8392 21888
rect 6788 21848 8392 21876
rect 6788 21836 6794 21848
rect 8386 21836 8392 21848
rect 8444 21836 8450 21888
rect 9309 21879 9367 21885
rect 9309 21845 9321 21879
rect 9355 21876 9367 21879
rect 9858 21876 9864 21888
rect 9355 21848 9864 21876
rect 9355 21845 9367 21848
rect 9309 21839 9367 21845
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 10229 21879 10287 21885
rect 10229 21876 10241 21879
rect 10008 21848 10241 21876
rect 10008 21836 10014 21848
rect 10229 21845 10241 21848
rect 10275 21845 10287 21879
rect 10229 21839 10287 21845
rect 11882 21836 11888 21888
rect 11940 21876 11946 21888
rect 12728 21876 12756 21916
rect 11940 21848 12756 21876
rect 12805 21879 12863 21885
rect 11940 21836 11946 21848
rect 12805 21845 12817 21879
rect 12851 21876 12863 21879
rect 12894 21876 12900 21888
rect 12851 21848 12900 21876
rect 12851 21845 12863 21848
rect 12805 21839 12863 21845
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 13096 21876 13124 21916
rect 13170 21904 13176 21956
rect 13228 21944 13234 21956
rect 13725 21947 13783 21953
rect 13725 21944 13737 21947
rect 13228 21916 13737 21944
rect 13228 21904 13234 21916
rect 13725 21913 13737 21916
rect 13771 21913 13783 21947
rect 15838 21944 15844 21956
rect 15778 21916 15844 21944
rect 13725 21907 13783 21913
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 13814 21876 13820 21888
rect 13096 21848 13820 21876
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14090 21836 14096 21888
rect 14148 21876 14154 21888
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 14148 21848 16037 21876
rect 14148 21836 14154 21848
rect 16025 21845 16037 21848
rect 16071 21876 16083 21879
rect 16500 21876 16528 22120
rect 17126 22040 17132 22092
rect 17184 22040 17190 22092
rect 18138 22080 18144 22092
rect 17236 22052 18144 22080
rect 17236 22012 17264 22052
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 18248 22089 18276 22120
rect 19794 22108 19800 22120
rect 19852 22108 19858 22160
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22049 18291 22083
rect 19981 22083 20039 22089
rect 19981 22080 19993 22083
rect 18233 22043 18291 22049
rect 18432 22052 19993 22080
rect 16960 21984 17264 22012
rect 16758 21904 16764 21956
rect 16816 21944 16822 21956
rect 16960 21953 16988 21984
rect 17494 21972 17500 22024
rect 17552 22012 17558 22024
rect 18432 22012 18460 22052
rect 19981 22049 19993 22052
rect 20027 22049 20039 22083
rect 19981 22043 20039 22049
rect 20714 22040 20720 22092
rect 20772 22080 20778 22092
rect 25148 22089 25176 22188
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 20772 22052 25053 22080
rect 20772 22040 20778 22052
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25041 22043 25099 22049
rect 25133 22083 25191 22089
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 17552 21984 18460 22012
rect 17552 21972 17558 21984
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19392 21984 20361 22012
rect 19392 21972 19398 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 22646 21972 22652 22024
rect 22704 21972 22710 22024
rect 24946 21972 24952 22024
rect 25004 21972 25010 22024
rect 16945 21947 17003 21953
rect 16945 21944 16957 21947
rect 16816 21916 16957 21944
rect 16816 21904 16822 21916
rect 16945 21913 16957 21916
rect 16991 21913 17003 21947
rect 16945 21907 17003 21913
rect 17126 21904 17132 21956
rect 17184 21944 17190 21956
rect 19150 21944 19156 21956
rect 17184 21916 19156 21944
rect 17184 21904 17190 21916
rect 16071 21848 16528 21876
rect 16071 21845 16083 21848
rect 16025 21839 16083 21845
rect 16850 21836 16856 21888
rect 16908 21836 16914 21888
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 18156 21885 18184 21916
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21944 19579 21947
rect 19610 21944 19616 21956
rect 19567 21916 19616 21944
rect 19567 21913 19579 21916
rect 19521 21907 19579 21913
rect 19610 21904 19616 21916
rect 19668 21904 19674 21956
rect 19702 21904 19708 21956
rect 19760 21904 19766 21956
rect 21082 21904 21088 21956
rect 21140 21904 21146 21956
rect 22186 21904 22192 21956
rect 22244 21944 22250 21956
rect 23474 21944 23480 21956
rect 22244 21916 23480 21944
rect 22244 21904 22250 21916
rect 23474 21904 23480 21916
rect 23532 21944 23538 21956
rect 23569 21947 23627 21953
rect 23569 21944 23581 21947
rect 23532 21916 23581 21944
rect 23532 21904 23538 21916
rect 23569 21913 23581 21916
rect 23615 21944 23627 21947
rect 23842 21944 23848 21956
rect 23615 21916 23848 21944
rect 23615 21913 23627 21916
rect 23569 21907 23627 21913
rect 23842 21904 23848 21916
rect 23900 21944 23906 21956
rect 24118 21944 24124 21956
rect 23900 21916 24124 21944
rect 23900 21904 23906 21916
rect 24118 21904 24124 21916
rect 24176 21944 24182 21956
rect 25222 21944 25228 21956
rect 24176 21916 25228 21944
rect 24176 21904 24182 21916
rect 25222 21904 25228 21916
rect 25280 21904 25286 21956
rect 18049 21879 18107 21885
rect 18049 21876 18061 21879
rect 17828 21848 18061 21876
rect 17828 21836 17834 21848
rect 18049 21845 18061 21848
rect 18095 21845 18107 21879
rect 18049 21839 18107 21845
rect 18141 21879 18199 21885
rect 18141 21845 18153 21879
rect 18187 21845 18199 21879
rect 18141 21839 18199 21845
rect 18230 21836 18236 21888
rect 18288 21876 18294 21888
rect 18877 21879 18935 21885
rect 18877 21876 18889 21879
rect 18288 21848 18889 21876
rect 18288 21836 18294 21848
rect 18877 21845 18889 21848
rect 18923 21876 18935 21879
rect 18966 21876 18972 21888
rect 18923 21848 18972 21876
rect 18923 21845 18935 21848
rect 18877 21839 18935 21845
rect 18966 21836 18972 21848
rect 19024 21836 19030 21888
rect 19168 21876 19196 21904
rect 20714 21876 20720 21888
rect 19168 21848 20720 21876
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 21910 21876 21916 21888
rect 21324 21848 21916 21876
rect 21324 21836 21330 21848
rect 21910 21836 21916 21848
rect 21968 21836 21974 21888
rect 22097 21879 22155 21885
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22370 21876 22376 21888
rect 22143 21848 22376 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22370 21836 22376 21848
rect 22428 21836 22434 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 22612 21848 24593 21876
rect 22612 21836 22618 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25406 21836 25412 21888
rect 25464 21876 25470 21888
rect 26142 21876 26148 21888
rect 25464 21848 26148 21876
rect 25464 21836 25470 21848
rect 26142 21836 26148 21848
rect 26200 21836 26206 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 1765 21675 1823 21681
rect 1765 21641 1777 21675
rect 1811 21672 1823 21675
rect 1811 21644 10916 21672
rect 1811 21641 1823 21644
rect 1765 21635 1823 21641
rect 1578 21564 1584 21616
rect 1636 21604 1642 21616
rect 1673 21607 1731 21613
rect 1673 21604 1685 21607
rect 1636 21576 1685 21604
rect 1636 21564 1642 21576
rect 1673 21573 1685 21576
rect 1719 21573 1731 21607
rect 1673 21567 1731 21573
rect 6549 21607 6607 21613
rect 6549 21573 6561 21607
rect 6595 21604 6607 21607
rect 9398 21604 9404 21616
rect 6595 21576 9404 21604
rect 6595 21573 6607 21576
rect 6549 21567 6607 21573
rect 9398 21564 9404 21576
rect 9456 21564 9462 21616
rect 10318 21564 10324 21616
rect 10376 21564 10382 21616
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21536 3019 21539
rect 3326 21536 3332 21548
rect 3007 21508 3332 21536
rect 3007 21505 3019 21508
rect 2961 21499 3019 21505
rect 3326 21496 3332 21508
rect 3384 21496 3390 21548
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 7374 21496 7380 21548
rect 7432 21496 7438 21548
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 10888 21536 10916 21644
rect 10962 21632 10968 21684
rect 11020 21672 11026 21684
rect 12621 21675 12679 21681
rect 12621 21672 12633 21675
rect 11020 21644 12633 21672
rect 11020 21632 11026 21644
rect 12621 21641 12633 21644
rect 12667 21641 12679 21675
rect 12621 21635 12679 21641
rect 12710 21632 12716 21684
rect 12768 21632 12774 21684
rect 13722 21632 13728 21684
rect 13780 21672 13786 21684
rect 13817 21675 13875 21681
rect 13817 21672 13829 21675
rect 13780 21644 13829 21672
rect 13780 21632 13786 21644
rect 13817 21641 13829 21644
rect 13863 21641 13875 21675
rect 13817 21635 13875 21641
rect 13906 21632 13912 21684
rect 13964 21672 13970 21684
rect 16666 21672 16672 21684
rect 13964 21644 16672 21672
rect 13964 21632 13970 21644
rect 16666 21632 16672 21644
rect 16724 21632 16730 21684
rect 18506 21632 18512 21684
rect 18564 21672 18570 21684
rect 20441 21675 20499 21681
rect 20441 21672 20453 21675
rect 18564 21644 20453 21672
rect 18564 21632 18570 21644
rect 20441 21641 20453 21644
rect 20487 21641 20499 21675
rect 20441 21635 20499 21641
rect 20530 21632 20536 21684
rect 20588 21672 20594 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 20588 21644 22017 21672
rect 20588 21632 20594 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22005 21635 22063 21641
rect 22373 21675 22431 21681
rect 22373 21641 22385 21675
rect 22419 21672 22431 21675
rect 23658 21672 23664 21684
rect 22419 21644 23664 21672
rect 22419 21641 22431 21644
rect 22373 21635 22431 21641
rect 11146 21564 11152 21616
rect 11204 21564 11210 21616
rect 11977 21607 12035 21613
rect 11977 21573 11989 21607
rect 12023 21604 12035 21607
rect 13078 21604 13084 21616
rect 12023 21576 13084 21604
rect 12023 21573 12035 21576
rect 11977 21567 12035 21573
rect 13078 21564 13084 21576
rect 13136 21564 13142 21616
rect 14277 21607 14335 21613
rect 14277 21573 14289 21607
rect 14323 21604 14335 21607
rect 17678 21604 17684 21616
rect 14323 21576 17684 21604
rect 14323 21573 14335 21576
rect 14277 21567 14335 21573
rect 17678 21564 17684 21576
rect 17736 21564 17742 21616
rect 20622 21564 20628 21616
rect 20680 21564 20686 21616
rect 20809 21607 20867 21613
rect 20809 21604 20821 21607
rect 20732 21576 20821 21604
rect 11882 21536 11888 21548
rect 10888 21508 11888 21536
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 13170 21536 13176 21548
rect 12912 21508 13176 21536
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 5074 21428 5080 21480
rect 5132 21428 5138 21480
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7340 21440 7665 21468
rect 7340 21428 7346 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 9309 21471 9367 21477
rect 9309 21437 9321 21471
rect 9355 21468 9367 21471
rect 11238 21468 11244 21480
rect 9355 21440 11244 21468
rect 9355 21437 9367 21440
rect 9309 21431 9367 21437
rect 11238 21428 11244 21440
rect 11296 21428 11302 21480
rect 11330 21428 11336 21480
rect 11388 21428 11394 21480
rect 11609 21471 11667 21477
rect 11609 21437 11621 21471
rect 11655 21468 11667 21471
rect 11698 21468 11704 21480
rect 11655 21440 11704 21468
rect 11655 21437 11667 21440
rect 11609 21431 11667 21437
rect 2317 21403 2375 21409
rect 2317 21369 2329 21403
rect 2363 21400 2375 21403
rect 4062 21400 4068 21412
rect 2363 21372 4068 21400
rect 2363 21369 2375 21372
rect 2317 21363 2375 21369
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 4246 21360 4252 21412
rect 4304 21400 4310 21412
rect 11348 21400 11376 21428
rect 4304 21372 7144 21400
rect 4304 21360 4310 21372
rect 2501 21335 2559 21341
rect 2501 21301 2513 21335
rect 2547 21332 2559 21335
rect 7006 21332 7012 21344
rect 2547 21304 7012 21332
rect 2547 21301 2559 21304
rect 2501 21295 2559 21301
rect 7006 21292 7012 21304
rect 7064 21292 7070 21344
rect 7116 21332 7144 21372
rect 10336 21372 11376 21400
rect 10336 21332 10364 21372
rect 7116 21304 10364 21332
rect 10502 21292 10508 21344
rect 10560 21332 10566 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 10560 21304 10793 21332
rect 10560 21292 10566 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 10781 21295 10839 21301
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11624 21332 11652 21431
rect 11698 21428 11704 21440
rect 11756 21468 11762 21480
rect 11756 21440 11836 21468
rect 11756 21428 11762 21440
rect 11808 21400 11836 21440
rect 12066 21428 12072 21480
rect 12124 21468 12130 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12124 21440 12817 21468
rect 12124 21428 12130 21440
rect 12805 21437 12817 21440
rect 12851 21437 12863 21471
rect 12805 21431 12863 21437
rect 11808 21372 12388 21400
rect 11808 21341 11836 21372
rect 11379 21304 11652 21332
rect 11793 21335 11851 21341
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11793 21301 11805 21335
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 12250 21292 12256 21344
rect 12308 21292 12314 21344
rect 12360 21332 12388 21372
rect 12434 21360 12440 21412
rect 12492 21400 12498 21412
rect 12912 21400 12940 21508
rect 13170 21496 13176 21508
rect 13228 21496 13234 21548
rect 14185 21539 14243 21545
rect 14185 21505 14197 21539
rect 14231 21536 14243 21539
rect 15102 21536 15108 21548
rect 14231 21508 15108 21536
rect 14231 21505 14243 21508
rect 14185 21499 14243 21505
rect 15102 21496 15108 21508
rect 15160 21496 15166 21548
rect 15194 21496 15200 21548
rect 15252 21536 15258 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 15252 21508 15393 21536
rect 15252 21496 15258 21508
rect 15381 21505 15393 21508
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 13446 21428 13452 21480
rect 13504 21468 13510 21480
rect 14369 21471 14427 21477
rect 14369 21468 14381 21471
rect 13504 21440 14381 21468
rect 13504 21428 13510 21440
rect 14369 21437 14381 21440
rect 14415 21437 14427 21471
rect 15488 21468 15516 21499
rect 15562 21496 15568 21548
rect 15620 21536 15626 21548
rect 15838 21536 15844 21548
rect 15620 21508 15844 21536
rect 15620 21496 15626 21508
rect 15838 21496 15844 21508
rect 15896 21536 15902 21548
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15896 21508 16129 21536
rect 15896 21496 15902 21508
rect 16117 21505 16129 21508
rect 16163 21536 16175 21539
rect 16298 21536 16304 21548
rect 16163 21508 16304 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 16298 21496 16304 21508
rect 16356 21496 16362 21548
rect 17034 21496 17040 21548
rect 17092 21536 17098 21548
rect 17405 21539 17463 21545
rect 17405 21536 17417 21539
rect 17092 21508 17417 21536
rect 17092 21496 17098 21508
rect 14369 21431 14427 21437
rect 14476 21440 15516 21468
rect 12492 21372 12940 21400
rect 13357 21403 13415 21409
rect 12492 21360 12498 21372
rect 13357 21369 13369 21403
rect 13403 21400 13415 21403
rect 13906 21400 13912 21412
rect 13403 21372 13912 21400
rect 13403 21369 13415 21372
rect 13357 21363 13415 21369
rect 13906 21360 13912 21372
rect 13964 21400 13970 21412
rect 14476 21400 14504 21440
rect 13964 21372 14504 21400
rect 15488 21400 15516 21440
rect 15654 21428 15660 21480
rect 15712 21428 15718 21480
rect 16482 21468 16488 21480
rect 16040 21440 16488 21468
rect 16040 21412 16068 21440
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 16022 21400 16028 21412
rect 15488 21372 16028 21400
rect 13964 21360 13970 21372
rect 16022 21360 16028 21372
rect 16080 21360 16086 21412
rect 16298 21360 16304 21412
rect 16356 21360 16362 21412
rect 16758 21360 16764 21412
rect 16816 21400 16822 21412
rect 17126 21400 17132 21412
rect 16816 21372 17132 21400
rect 16816 21360 16822 21372
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 17236 21400 17264 21508
rect 17405 21505 17417 21508
rect 17451 21505 17463 21539
rect 17405 21499 17463 21505
rect 17494 21496 17500 21548
rect 17552 21496 17558 21548
rect 18233 21539 18291 21545
rect 18233 21505 18245 21539
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 17310 21428 17316 21480
rect 17368 21468 17374 21480
rect 17589 21471 17647 21477
rect 17589 21468 17601 21471
rect 17368 21440 17601 21468
rect 17368 21428 17374 21440
rect 17589 21437 17601 21440
rect 17635 21437 17647 21471
rect 17589 21431 17647 21437
rect 17862 21400 17868 21412
rect 17236 21372 17868 21400
rect 17862 21360 17868 21372
rect 17920 21360 17926 21412
rect 18248 21400 18276 21499
rect 18966 21496 18972 21548
rect 19024 21536 19030 21548
rect 20640 21536 20668 21564
rect 19024 21508 20668 21536
rect 19024 21496 19030 21508
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 20257 21471 20315 21477
rect 20257 21468 20269 21471
rect 18380 21440 20269 21468
rect 18380 21428 18386 21440
rect 20257 21437 20269 21440
rect 20303 21468 20315 21471
rect 20732 21468 20760 21576
rect 20809 21573 20821 21576
rect 20855 21573 20867 21607
rect 20809 21567 20867 21573
rect 20898 21564 20904 21616
rect 20956 21604 20962 21616
rect 21450 21604 21456 21616
rect 20956 21576 21456 21604
rect 20956 21564 20962 21576
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 21726 21564 21732 21616
rect 21784 21604 21790 21616
rect 22388 21604 22416 21635
rect 23658 21632 23664 21644
rect 23716 21672 23722 21684
rect 23842 21672 23848 21684
rect 23716 21644 23848 21672
rect 23716 21632 23722 21644
rect 23842 21632 23848 21644
rect 23900 21632 23906 21684
rect 21784 21576 22416 21604
rect 21784 21564 21790 21576
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 23290 21496 23296 21548
rect 23348 21536 23354 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23348 21508 23397 21536
rect 23348 21496 23354 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 20303 21440 20760 21468
rect 20303 21437 20315 21440
rect 20257 21431 20315 21437
rect 20990 21428 20996 21480
rect 21048 21428 21054 21480
rect 21726 21428 21732 21480
rect 21784 21468 21790 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 21784 21440 22477 21468
rect 21784 21428 21790 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22557 21471 22615 21477
rect 22557 21437 22569 21471
rect 22603 21437 22615 21471
rect 22557 21431 22615 21437
rect 23661 21471 23719 21477
rect 23661 21437 23673 21471
rect 23707 21468 23719 21471
rect 24854 21468 24860 21480
rect 23707 21440 24860 21468
rect 23707 21437 23719 21440
rect 23661 21431 23719 21437
rect 21542 21400 21548 21412
rect 18248 21372 21548 21400
rect 21542 21360 21548 21372
rect 21600 21360 21606 21412
rect 12526 21332 12532 21344
rect 12360 21304 12532 21332
rect 12526 21292 12532 21304
rect 12584 21332 12590 21344
rect 12894 21332 12900 21344
rect 12584 21304 12900 21332
rect 12584 21292 12590 21304
rect 12894 21292 12900 21304
rect 12952 21332 12958 21344
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 12952 21304 13553 21332
rect 12952 21292 12958 21304
rect 13541 21301 13553 21304
rect 13587 21332 13599 21335
rect 14734 21332 14740 21344
rect 13587 21304 14740 21332
rect 13587 21301 13599 21304
rect 13541 21295 13599 21301
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 14918 21292 14924 21344
rect 14976 21332 14982 21344
rect 15013 21335 15071 21341
rect 15013 21332 15025 21335
rect 14976 21304 15025 21332
rect 14976 21292 14982 21304
rect 15013 21301 15025 21304
rect 15059 21301 15071 21335
rect 15013 21295 15071 21301
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 16393 21335 16451 21341
rect 16393 21332 16405 21335
rect 16264 21304 16405 21332
rect 16264 21292 16270 21304
rect 16393 21301 16405 21304
rect 16439 21301 16451 21335
rect 16393 21295 16451 21301
rect 17034 21292 17040 21344
rect 17092 21292 17098 21344
rect 17144 21332 17172 21360
rect 17494 21332 17500 21344
rect 17144 21304 17500 21332
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19392 21304 19533 21332
rect 19392 21292 19398 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 19521 21295 19579 21301
rect 20254 21292 20260 21344
rect 20312 21332 20318 21344
rect 22572 21332 22600 21431
rect 24854 21428 24860 21440
rect 24912 21428 24918 21480
rect 20312 21304 22600 21332
rect 20312 21292 20318 21304
rect 22830 21292 22836 21344
rect 22888 21332 22894 21344
rect 23017 21335 23075 21341
rect 23017 21332 23029 21335
rect 22888 21304 23029 21332
rect 22888 21292 22894 21304
rect 23017 21301 23029 21304
rect 23063 21301 23075 21335
rect 23017 21295 23075 21301
rect 23750 21292 23756 21344
rect 23808 21332 23814 21344
rect 25133 21335 25191 21341
rect 25133 21332 25145 21335
rect 23808 21304 25145 21332
rect 23808 21292 23814 21304
rect 25133 21301 25145 21304
rect 25179 21301 25191 21335
rect 25133 21295 25191 21301
rect 25406 21292 25412 21344
rect 25464 21292 25470 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 1581 21131 1639 21137
rect 1581 21097 1593 21131
rect 1627 21128 1639 21131
rect 1627 21100 3280 21128
rect 1627 21097 1639 21100
rect 1581 21091 1639 21097
rect 2240 20964 2774 20992
rect 2240 20933 2268 20964
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 2746 20856 2774 20964
rect 2866 20952 2872 21004
rect 2924 20952 2930 21004
rect 3252 20992 3280 21100
rect 3326 21088 3332 21140
rect 3384 21128 3390 21140
rect 9309 21131 9367 21137
rect 9309 21128 9321 21131
rect 3384 21100 9321 21128
rect 3384 21088 3390 21100
rect 9309 21097 9321 21100
rect 9355 21097 9367 21131
rect 12897 21131 12955 21137
rect 9309 21091 9367 21097
rect 10520 21100 12848 21128
rect 8478 21020 8484 21072
rect 8536 21060 8542 21072
rect 9953 21063 10011 21069
rect 9953 21060 9965 21063
rect 8536 21032 9965 21060
rect 8536 21020 8542 21032
rect 9953 21029 9965 21032
rect 9999 21029 10011 21063
rect 10520 21060 10548 21100
rect 9953 21023 10011 21029
rect 10428 21032 10548 21060
rect 12820 21060 12848 21100
rect 12897 21097 12909 21131
rect 12943 21128 12955 21131
rect 13538 21128 13544 21140
rect 12943 21100 13544 21128
rect 12943 21097 12955 21100
rect 12897 21091 12955 21097
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 13630 21088 13636 21140
rect 13688 21088 13694 21140
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 16206 21128 16212 21140
rect 15252 21100 16212 21128
rect 15252 21088 15258 21100
rect 16206 21088 16212 21100
rect 16264 21088 16270 21140
rect 16666 21088 16672 21140
rect 16724 21088 16730 21140
rect 17218 21088 17224 21140
rect 17276 21128 17282 21140
rect 17865 21131 17923 21137
rect 17865 21128 17877 21131
rect 17276 21100 17877 21128
rect 17276 21088 17282 21100
rect 17865 21097 17877 21100
rect 17911 21097 17923 21131
rect 17865 21091 17923 21097
rect 18414 21088 18420 21140
rect 18472 21128 18478 21140
rect 18966 21128 18972 21140
rect 18472 21100 18972 21128
rect 18472 21088 18478 21100
rect 18966 21088 18972 21100
rect 19024 21088 19030 21140
rect 19518 21088 19524 21140
rect 19576 21088 19582 21140
rect 21174 21088 21180 21140
rect 21232 21088 21238 21140
rect 21358 21088 21364 21140
rect 21416 21128 21422 21140
rect 21416 21100 25176 21128
rect 21416 21088 21422 21100
rect 15473 21063 15531 21069
rect 15473 21060 15485 21063
rect 12820 21032 15485 21060
rect 4246 20992 4252 21004
rect 3252 20964 4252 20992
rect 4246 20952 4252 20964
rect 4304 20952 4310 21004
rect 4338 20952 4344 21004
rect 4396 20992 4402 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4396 20964 4445 20992
rect 4396 20952 4402 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 6972 20964 7389 20992
rect 6972 20952 6978 20964
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 7377 20955 7435 20961
rect 8754 20952 8760 21004
rect 8812 20952 8818 21004
rect 10428 21001 10456 21032
rect 15473 21029 15485 21032
rect 15519 21029 15531 21063
rect 18322 21060 18328 21072
rect 15473 21023 15531 21029
rect 16224 21032 18328 21060
rect 16224 21004 16252 21032
rect 18322 21020 18328 21032
rect 18380 21020 18386 21072
rect 19536 21060 19564 21088
rect 18432 21032 19564 21060
rect 10413 20995 10471 21001
rect 10413 20961 10425 20995
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 10502 20952 10508 21004
rect 10560 20952 10566 21004
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 11112 20964 11161 20992
rect 11112 20952 11118 20964
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20992 11483 20995
rect 12066 20992 12072 21004
rect 11471 20964 12072 20992
rect 11471 20961 11483 20964
rect 11425 20955 11483 20961
rect 12066 20952 12072 20964
rect 12124 20992 12130 21004
rect 12802 20992 12808 21004
rect 12124 20964 12808 20992
rect 12124 20952 12130 20964
rect 12802 20952 12808 20964
rect 12860 20952 12866 21004
rect 12894 20952 12900 21004
rect 12952 20992 12958 21004
rect 16025 20995 16083 21001
rect 16025 20992 16037 20995
rect 12952 20964 16037 20992
rect 12952 20952 12958 20964
rect 16025 20961 16037 20964
rect 16071 20961 16083 20995
rect 16025 20955 16083 20961
rect 16206 20952 16212 21004
rect 16264 20952 16270 21004
rect 16390 20952 16396 21004
rect 16448 20992 16454 21004
rect 17221 20995 17279 21001
rect 17221 20992 17233 20995
rect 16448 20964 17233 20992
rect 16448 20952 16454 20964
rect 17221 20961 17233 20964
rect 17267 20961 17279 20995
rect 17221 20955 17279 20961
rect 4154 20884 4160 20936
rect 4212 20884 4218 20936
rect 5813 20927 5871 20933
rect 5813 20893 5825 20927
rect 5859 20924 5871 20927
rect 7006 20924 7012 20936
rect 5859 20896 7012 20924
rect 5859 20893 5871 20896
rect 5813 20887 5871 20893
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 7098 20884 7104 20936
rect 7156 20884 7162 20936
rect 12526 20884 12532 20936
rect 12584 20884 12590 20936
rect 12710 20884 12716 20936
rect 12768 20924 12774 20936
rect 12768 20896 13308 20924
rect 12768 20884 12774 20896
rect 2746 20828 6592 20856
rect 1765 20791 1823 20797
rect 1765 20757 1777 20791
rect 1811 20788 1823 20791
rect 1946 20788 1952 20800
rect 1811 20760 1952 20788
rect 1811 20757 1823 20760
rect 1765 20751 1823 20757
rect 1946 20748 1952 20760
rect 2004 20788 2010 20800
rect 2406 20788 2412 20800
rect 2004 20760 2412 20788
rect 2004 20748 2010 20760
rect 2406 20748 2412 20760
rect 2464 20748 2470 20800
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 5626 20788 5632 20800
rect 3108 20760 5632 20788
rect 3108 20748 3114 20760
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 6454 20748 6460 20800
rect 6512 20748 6518 20800
rect 6564 20788 6592 20828
rect 6638 20816 6644 20868
rect 6696 20856 6702 20868
rect 9217 20859 9275 20865
rect 9217 20856 9229 20859
rect 6696 20828 9229 20856
rect 6696 20816 6702 20828
rect 9217 20825 9229 20828
rect 9263 20825 9275 20859
rect 13280 20856 13308 20896
rect 13998 20884 14004 20936
rect 14056 20924 14062 20936
rect 14274 20924 14280 20936
rect 14056 20896 14280 20924
rect 14056 20884 14062 20896
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 16298 20924 16304 20936
rect 14415 20896 16304 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 17126 20884 17132 20936
rect 17184 20924 17190 20936
rect 17402 20924 17408 20936
rect 17184 20896 17408 20924
rect 17184 20884 17190 20896
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 18233 20927 18291 20933
rect 18233 20893 18245 20927
rect 18279 20924 18291 20927
rect 18432 20924 18460 21032
rect 21450 21020 21456 21072
rect 21508 21060 21514 21072
rect 24581 21063 24639 21069
rect 21508 21032 24440 21060
rect 21508 21020 21514 21032
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18690 20992 18696 21004
rect 18555 20964 18696 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18690 20952 18696 20964
rect 18748 20992 18754 21004
rect 19705 20995 19763 21001
rect 19705 20992 19717 20995
rect 18748 20964 19717 20992
rect 18748 20952 18754 20964
rect 19705 20961 19717 20964
rect 19751 20961 19763 20995
rect 19705 20955 19763 20961
rect 21634 20952 21640 21004
rect 21692 20992 21698 21004
rect 22189 20995 22247 21001
rect 22189 20992 22201 20995
rect 21692 20964 22201 20992
rect 21692 20952 21698 20964
rect 22189 20961 22201 20964
rect 22235 20961 22247 20995
rect 22189 20955 22247 20961
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 23017 20995 23075 21001
rect 23017 20992 23029 20995
rect 22787 20964 23029 20992
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 23017 20961 23029 20964
rect 23063 20992 23075 20995
rect 23474 20992 23480 21004
rect 23063 20964 23480 20992
rect 23063 20961 23075 20964
rect 23017 20955 23075 20961
rect 23474 20952 23480 20964
rect 23532 20952 23538 21004
rect 24412 20992 24440 21032
rect 24581 21029 24593 21063
rect 24627 21060 24639 21063
rect 24670 21060 24676 21072
rect 24627 21032 24676 21060
rect 24627 21029 24639 21032
rect 24581 21023 24639 21029
rect 24670 21020 24676 21032
rect 24728 21020 24734 21072
rect 25148 21001 25176 21100
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 24412 20964 25053 20992
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 18279 20896 18460 20924
rect 18279 20893 18291 20896
rect 18233 20887 18291 20893
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19392 20896 19441 20924
rect 19392 20884 19398 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20924 23903 20927
rect 24026 20924 24032 20936
rect 23891 20896 24032 20924
rect 23891 20893 23903 20896
rect 23845 20887 23903 20893
rect 24026 20884 24032 20896
rect 24084 20884 24090 20936
rect 13541 20859 13599 20865
rect 13541 20856 13553 20859
rect 13280 20828 13553 20856
rect 9217 20819 9275 20825
rect 13541 20825 13553 20828
rect 13587 20825 13599 20859
rect 15194 20856 15200 20868
rect 13541 20819 13599 20825
rect 13924 20828 15200 20856
rect 8294 20788 8300 20800
rect 6564 20760 8300 20788
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 9950 20788 9956 20800
rect 9824 20760 9956 20788
rect 9824 20748 9830 20760
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 10321 20791 10379 20797
rect 10321 20757 10333 20791
rect 10367 20788 10379 20791
rect 10410 20788 10416 20800
rect 10367 20760 10416 20788
rect 10367 20757 10379 20760
rect 10321 20751 10379 20757
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 11238 20748 11244 20800
rect 11296 20788 11302 20800
rect 12894 20788 12900 20800
rect 11296 20760 12900 20788
rect 11296 20748 11302 20760
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 13170 20748 13176 20800
rect 13228 20788 13234 20800
rect 13924 20788 13952 20828
rect 15194 20816 15200 20828
rect 15252 20816 15258 20868
rect 15933 20859 15991 20865
rect 15933 20825 15945 20859
rect 15979 20856 15991 20859
rect 16758 20856 16764 20868
rect 15979 20828 16764 20856
rect 15979 20825 15991 20828
rect 15933 20819 15991 20825
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 17037 20859 17095 20865
rect 17037 20825 17049 20859
rect 17083 20856 17095 20859
rect 17678 20856 17684 20868
rect 17083 20828 17684 20856
rect 17083 20825 17095 20828
rect 17037 20819 17095 20825
rect 17678 20816 17684 20828
rect 17736 20816 17742 20868
rect 18325 20859 18383 20865
rect 18325 20825 18337 20859
rect 18371 20856 18383 20859
rect 19978 20856 19984 20868
rect 18371 20828 19984 20856
rect 18371 20825 18383 20828
rect 18325 20819 18383 20825
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 21082 20856 21088 20868
rect 20930 20828 21088 20856
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 21266 20816 21272 20868
rect 21324 20856 21330 20868
rect 22097 20859 22155 20865
rect 22097 20856 22109 20859
rect 21324 20828 22109 20856
rect 21324 20816 21330 20828
rect 22097 20825 22109 20828
rect 22143 20856 22155 20859
rect 22833 20859 22891 20865
rect 22833 20856 22845 20859
rect 22143 20828 22845 20856
rect 22143 20825 22155 20828
rect 22097 20819 22155 20825
rect 22833 20825 22845 20828
rect 22879 20825 22891 20859
rect 22833 20819 22891 20825
rect 23198 20816 23204 20868
rect 23256 20816 23262 20868
rect 24489 20859 24547 20865
rect 24489 20825 24501 20859
rect 24535 20856 24547 20859
rect 24578 20856 24584 20868
rect 24535 20828 24584 20856
rect 24535 20825 24547 20828
rect 24489 20819 24547 20825
rect 24578 20816 24584 20828
rect 24636 20856 24642 20868
rect 24949 20859 25007 20865
rect 24949 20856 24961 20859
rect 24636 20828 24961 20856
rect 24636 20816 24642 20828
rect 24949 20825 24961 20828
rect 24995 20825 25007 20859
rect 24949 20819 25007 20825
rect 13228 20760 13952 20788
rect 13228 20748 13234 20760
rect 13998 20748 14004 20800
rect 14056 20788 14062 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 14056 20760 15025 20788
rect 14056 20748 14062 20760
rect 15013 20757 15025 20760
rect 15059 20757 15071 20791
rect 15013 20751 15071 20757
rect 15838 20748 15844 20800
rect 15896 20748 15902 20800
rect 16022 20748 16028 20800
rect 16080 20788 16086 20800
rect 17129 20791 17187 20797
rect 17129 20788 17141 20791
rect 16080 20760 17141 20788
rect 16080 20748 16086 20760
rect 17129 20757 17141 20760
rect 17175 20757 17187 20791
rect 17129 20751 17187 20757
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21450 20788 21456 20800
rect 21232 20760 21456 20788
rect 21232 20748 21238 20760
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 21637 20791 21695 20797
rect 21637 20757 21649 20791
rect 21683 20788 21695 20791
rect 21910 20788 21916 20800
rect 21683 20760 21916 20788
rect 21683 20757 21695 20760
rect 21637 20751 21695 20757
rect 21910 20748 21916 20760
rect 21968 20748 21974 20800
rect 22002 20748 22008 20800
rect 22060 20748 22066 20800
rect 23477 20791 23535 20797
rect 23477 20757 23489 20791
rect 23523 20788 23535 20791
rect 23658 20788 23664 20800
rect 23523 20760 23664 20788
rect 23523 20757 23535 20760
rect 23477 20751 23535 20757
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 23842 20748 23848 20800
rect 23900 20788 23906 20800
rect 23937 20791 23995 20797
rect 23937 20788 23949 20791
rect 23900 20760 23949 20788
rect 23900 20748 23906 20760
rect 23937 20757 23949 20760
rect 23983 20788 23995 20791
rect 24118 20788 24124 20800
rect 23983 20760 24124 20788
rect 23983 20757 23995 20760
rect 23937 20751 23995 20757
rect 24118 20748 24124 20760
rect 24176 20748 24182 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 26050 20680 26056 20732
rect 26108 20720 26114 20732
rect 26418 20720 26424 20732
rect 26108 20692 26424 20720
rect 26108 20680 26114 20692
rect 26418 20680 26424 20692
rect 26476 20680 26482 20732
rect 1104 20624 25852 20646
rect 2225 20587 2283 20593
rect 2225 20553 2237 20587
rect 2271 20584 2283 20587
rect 6549 20587 6607 20593
rect 2271 20556 2774 20584
rect 2271 20553 2283 20556
rect 2225 20547 2283 20553
rect 1670 20476 1676 20528
rect 1728 20476 1734 20528
rect 2746 20516 2774 20556
rect 6549 20553 6561 20587
rect 6595 20584 6607 20587
rect 7466 20584 7472 20596
rect 6595 20556 7472 20584
rect 6595 20553 6607 20556
rect 6549 20547 6607 20553
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 11514 20584 11520 20596
rect 8496 20556 11520 20584
rect 3602 20516 3608 20528
rect 2746 20488 3608 20516
rect 3602 20476 3608 20488
rect 3660 20516 3666 20528
rect 4801 20519 4859 20525
rect 4801 20516 4813 20519
rect 3660 20488 4813 20516
rect 3660 20476 3666 20488
rect 4801 20485 4813 20488
rect 4847 20485 4859 20519
rect 8386 20516 8392 20528
rect 4801 20479 4859 20485
rect 6840 20488 8392 20516
rect 3050 20408 3056 20460
rect 3108 20408 3114 20460
rect 6840 20457 6868 20488
rect 8386 20476 8392 20488
rect 8444 20476 8450 20528
rect 6181 20451 6239 20457
rect 6181 20417 6193 20451
rect 6227 20448 6239 20451
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 6227 20420 6837 20448
rect 6227 20417 6239 20420
rect 6181 20411 6239 20417
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20448 7987 20451
rect 8496 20448 8524 20556
rect 11514 20544 11520 20556
rect 11572 20544 11578 20596
rect 11698 20544 11704 20596
rect 11756 20544 11762 20596
rect 12434 20544 12440 20596
rect 12492 20544 12498 20596
rect 13170 20584 13176 20596
rect 13004 20556 13176 20584
rect 8573 20519 8631 20525
rect 8573 20485 8585 20519
rect 8619 20516 8631 20519
rect 9306 20516 9312 20528
rect 8619 20488 9312 20516
rect 8619 20485 8631 20488
rect 8573 20479 8631 20485
rect 9306 20476 9312 20488
rect 9364 20476 9370 20528
rect 10594 20476 10600 20528
rect 10652 20516 10658 20528
rect 11149 20519 11207 20525
rect 11149 20516 11161 20519
rect 10652 20488 11161 20516
rect 10652 20476 10658 20488
rect 11149 20485 11161 20488
rect 11195 20516 11207 20519
rect 11606 20516 11612 20528
rect 11195 20488 11612 20516
rect 11195 20485 11207 20488
rect 11149 20479 11207 20485
rect 11606 20476 11612 20488
rect 11664 20476 11670 20528
rect 7975 20420 8524 20448
rect 7975 20417 7987 20420
rect 7929 20411 7987 20417
rect 9030 20408 9036 20460
rect 9088 20408 9094 20460
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 11241 20451 11299 20457
rect 11241 20448 11253 20451
rect 10376 20420 11253 20448
rect 10376 20408 10382 20420
rect 11241 20417 11253 20420
rect 11287 20448 11299 20451
rect 11716 20448 11744 20544
rect 11882 20476 11888 20528
rect 11940 20516 11946 20528
rect 13004 20516 13032 20556
rect 13170 20544 13176 20556
rect 13228 20544 13234 20596
rect 13906 20584 13912 20596
rect 13464 20556 13912 20584
rect 11940 20488 13032 20516
rect 11940 20476 11946 20488
rect 13464 20448 13492 20556
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 15470 20584 15476 20596
rect 14792 20556 15476 20584
rect 14792 20544 14798 20556
rect 13804 20519 13862 20525
rect 13804 20485 13816 20519
rect 13850 20516 13862 20519
rect 14090 20516 14096 20528
rect 13850 20488 14096 20516
rect 13850 20485 13862 20488
rect 13804 20479 13862 20485
rect 14090 20476 14096 20488
rect 14148 20476 14154 20528
rect 15120 20516 15148 20556
rect 15470 20544 15476 20556
rect 15528 20544 15534 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18012 20556 18368 20584
rect 18012 20544 18018 20556
rect 15042 20488 15148 20516
rect 15194 20476 15200 20528
rect 15252 20516 15258 20528
rect 15565 20519 15623 20525
rect 15565 20516 15577 20519
rect 15252 20488 15577 20516
rect 15252 20476 15258 20488
rect 15565 20485 15577 20488
rect 15611 20485 15623 20519
rect 15565 20479 15623 20485
rect 16758 20476 16764 20528
rect 16816 20516 16822 20528
rect 16816 20488 16988 20516
rect 16816 20476 16822 20488
rect 11287 20420 11744 20448
rect 12268 20420 13492 20448
rect 11287 20417 11299 20420
rect 11241 20411 11299 20417
rect 2590 20340 2596 20392
rect 2648 20340 2654 20392
rect 3418 20340 3424 20392
rect 3476 20340 3482 20392
rect 5537 20383 5595 20389
rect 5537 20349 5549 20383
rect 5583 20380 5595 20383
rect 8938 20380 8944 20392
rect 5583 20352 8944 20380
rect 5583 20349 5595 20352
rect 5537 20343 5595 20349
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 9309 20383 9367 20389
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 10502 20380 10508 20392
rect 9355 20352 10508 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 1857 20315 1915 20321
rect 1857 20281 1869 20315
rect 1903 20312 1915 20315
rect 12268 20312 12296 20420
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 16960 20457 16988 20488
rect 18340 20460 18368 20556
rect 18690 20544 18696 20596
rect 18748 20544 18754 20596
rect 20438 20544 20444 20596
rect 20496 20584 20502 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20496 20556 21005 20584
rect 20496 20544 20502 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 20993 20547 21051 20553
rect 21082 20544 21088 20596
rect 21140 20584 21146 20596
rect 21269 20587 21327 20593
rect 21269 20584 21281 20587
rect 21140 20556 21281 20584
rect 21140 20544 21146 20556
rect 21269 20553 21281 20556
rect 21315 20584 21327 20587
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 21315 20556 21465 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 22002 20584 22008 20596
rect 21876 20556 22008 20584
rect 21876 20544 21882 20556
rect 22002 20544 22008 20556
rect 22060 20584 22066 20596
rect 22465 20587 22523 20593
rect 22465 20584 22477 20587
rect 22060 20556 22477 20584
rect 22060 20544 22066 20556
rect 22465 20553 22477 20556
rect 22511 20553 22523 20587
rect 22465 20547 22523 20553
rect 23198 20544 23204 20596
rect 23256 20584 23262 20596
rect 23382 20584 23388 20596
rect 23256 20556 23388 20584
rect 23256 20544 23262 20556
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 23474 20544 23480 20596
rect 23532 20584 23538 20596
rect 23532 20556 23888 20584
rect 23532 20544 23538 20556
rect 18598 20476 18604 20528
rect 18656 20516 18662 20528
rect 19978 20516 19984 20528
rect 18656 20488 19984 20516
rect 18656 20476 18662 20488
rect 19978 20476 19984 20488
rect 20036 20476 20042 20528
rect 21100 20516 21128 20544
rect 20746 20502 21128 20516
rect 20732 20488 21128 20502
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 16945 20451 17003 20457
rect 16163 20420 16896 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 12529 20383 12587 20389
rect 12529 20380 12541 20383
rect 1903 20284 8708 20312
rect 1903 20281 1915 20284
rect 1857 20275 1915 20281
rect 2406 20204 2412 20256
rect 2464 20204 2470 20256
rect 4062 20204 4068 20256
rect 4120 20244 4126 20256
rect 4893 20247 4951 20253
rect 4893 20244 4905 20247
rect 4120 20216 4905 20244
rect 4120 20204 4126 20216
rect 4893 20213 4905 20216
rect 4939 20244 4951 20247
rect 5350 20244 5356 20256
rect 4939 20216 5356 20244
rect 4939 20213 4951 20216
rect 4893 20207 4951 20213
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7469 20247 7527 20253
rect 7469 20244 7481 20247
rect 6972 20216 7481 20244
rect 6972 20204 6978 20216
rect 7469 20213 7481 20216
rect 7515 20213 7527 20247
rect 8680 20244 8708 20284
rect 10704 20284 12296 20312
rect 12360 20352 12541 20380
rect 10704 20244 10732 20284
rect 8680 20216 10732 20244
rect 7469 20207 7527 20213
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 11940 20216 12081 20244
rect 11940 20204 11946 20216
rect 12069 20213 12081 20216
rect 12115 20213 12127 20247
rect 12360 20244 12388 20352
rect 12529 20349 12541 20352
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 12621 20383 12679 20389
rect 12621 20349 12633 20383
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 12434 20272 12440 20324
rect 12492 20312 12498 20324
rect 12636 20312 12664 20343
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 15289 20383 15347 20389
rect 15289 20380 15301 20383
rect 13504 20352 15301 20380
rect 13504 20340 13510 20352
rect 15289 20349 15301 20352
rect 15335 20349 15347 20383
rect 15289 20343 15347 20349
rect 12492 20284 12664 20312
rect 12492 20272 12498 20284
rect 16022 20244 16028 20256
rect 12360 20216 16028 20244
rect 12069 20207 12127 20213
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 16206 20204 16212 20256
rect 16264 20204 16270 20256
rect 16868 20244 16896 20420
rect 16945 20417 16957 20451
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 18322 20408 18328 20460
rect 18380 20408 18386 20460
rect 20732 20392 20760 20488
rect 23750 20476 23756 20528
rect 23808 20476 23814 20528
rect 23860 20516 23888 20556
rect 24026 20516 24032 20528
rect 23860 20488 24032 20516
rect 24026 20476 24032 20488
rect 24084 20516 24090 20528
rect 24084 20488 24242 20516
rect 24084 20476 24090 20488
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23477 20451 23535 20457
rect 23477 20448 23489 20451
rect 23348 20420 23489 20448
rect 23348 20408 23354 20420
rect 23477 20417 23489 20420
rect 23523 20417 23535 20451
rect 23477 20411 23535 20417
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 17276 20352 18828 20380
rect 17276 20340 17282 20352
rect 18230 20244 18236 20256
rect 16868 20216 18236 20244
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 18800 20244 18828 20352
rect 19242 20340 19248 20392
rect 19300 20340 19306 20392
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19886 20380 19892 20392
rect 19567 20352 19892 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 19978 20340 19984 20392
rect 20036 20380 20042 20392
rect 20714 20380 20720 20392
rect 20036 20352 20720 20380
rect 20036 20340 20042 20352
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 22646 20340 22652 20392
rect 22704 20340 22710 20392
rect 21358 20312 21364 20324
rect 20548 20284 21364 20312
rect 20548 20244 20576 20284
rect 21358 20272 21364 20284
rect 21416 20272 21422 20324
rect 22572 20312 22600 20340
rect 23109 20315 23167 20321
rect 23109 20312 23121 20315
rect 22572 20284 23121 20312
rect 23109 20281 23121 20284
rect 23155 20281 23167 20315
rect 23109 20275 23167 20281
rect 18800 20216 20576 20244
rect 22097 20247 22155 20253
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 23842 20244 23848 20256
rect 22143 20216 23848 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 25222 20204 25228 20256
rect 25280 20204 25286 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 1394 20000 1400 20052
rect 1452 20040 1458 20052
rect 1489 20043 1547 20049
rect 1489 20040 1501 20043
rect 1452 20012 1501 20040
rect 1452 20000 1458 20012
rect 1489 20009 1501 20012
rect 1535 20009 1547 20043
rect 1489 20003 1547 20009
rect 1670 20000 1676 20052
rect 1728 20000 1734 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 5261 20043 5319 20049
rect 5261 20040 5273 20043
rect 4212 20012 5273 20040
rect 4212 20000 4218 20012
rect 5261 20009 5273 20012
rect 5307 20009 5319 20043
rect 5261 20003 5319 20009
rect 6638 20000 6644 20052
rect 6696 20000 6702 20052
rect 7282 20000 7288 20052
rect 7340 20000 7346 20052
rect 9033 20043 9091 20049
rect 9033 20009 9045 20043
rect 9079 20040 9091 20043
rect 9214 20040 9220 20052
rect 9079 20012 9220 20040
rect 9079 20009 9091 20012
rect 9033 20003 9091 20009
rect 9214 20000 9220 20012
rect 9272 20000 9278 20052
rect 9306 20000 9312 20052
rect 9364 20040 9370 20052
rect 10778 20040 10784 20052
rect 9364 20012 10784 20040
rect 9364 20000 9370 20012
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 11204 20012 14933 20040
rect 11204 20000 11210 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 16080 20012 17693 20040
rect 16080 20000 16086 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 20533 20043 20591 20049
rect 17681 20003 17739 20009
rect 17788 20012 20024 20040
rect 6822 19972 6828 19984
rect 2746 19944 6828 19972
rect 2746 19904 2774 19944
rect 6822 19932 6828 19944
rect 6880 19932 6886 19984
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 10594 19972 10600 19984
rect 8904 19944 10600 19972
rect 8904 19932 8910 19944
rect 10594 19932 10600 19944
rect 10652 19932 10658 19984
rect 10796 19972 10824 20000
rect 10796 19944 11100 19972
rect 2240 19876 2774 19904
rect 3973 19907 4031 19913
rect 2240 19845 2268 19876
rect 3973 19873 3985 19907
rect 4019 19904 4031 19907
rect 4430 19904 4436 19916
rect 4019 19876 4436 19904
rect 4019 19873 4031 19876
rect 3973 19867 4031 19873
rect 4430 19864 4436 19876
rect 4488 19864 4494 19916
rect 6086 19864 6092 19916
rect 6144 19904 6150 19916
rect 6144 19876 6868 19904
rect 6144 19864 6150 19876
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 4246 19796 4252 19848
rect 4304 19796 4310 19848
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 6546 19836 6552 19848
rect 5491 19808 6552 19836
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 6840 19845 6868 19876
rect 8938 19864 8944 19916
rect 8996 19904 9002 19916
rect 8996 19876 10824 19904
rect 8996 19864 9002 19876
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 7466 19796 7472 19848
rect 7524 19796 7530 19848
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 8754 19836 8760 19848
rect 7975 19808 8760 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 8754 19796 8760 19808
rect 8812 19796 8818 19848
rect 9214 19796 9220 19848
rect 9272 19836 9278 19848
rect 10796 19845 10824 19876
rect 10962 19864 10968 19916
rect 11020 19864 11026 19916
rect 11072 19904 11100 19944
rect 12894 19932 12900 19984
rect 12952 19972 12958 19984
rect 13357 19975 13415 19981
rect 13357 19972 13369 19975
rect 12952 19944 13369 19972
rect 12952 19932 12958 19944
rect 13357 19941 13369 19944
rect 13403 19941 13415 19975
rect 13357 19935 13415 19941
rect 13722 19932 13728 19984
rect 13780 19972 13786 19984
rect 13909 19975 13967 19981
rect 13909 19972 13921 19975
rect 13780 19944 13921 19972
rect 13780 19932 13786 19944
rect 13909 19941 13921 19944
rect 13955 19972 13967 19975
rect 14090 19972 14096 19984
rect 13955 19944 14096 19972
rect 13955 19941 13967 19944
rect 13909 19935 13967 19941
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 14458 19932 14464 19984
rect 14516 19972 14522 19984
rect 16390 19972 16396 19984
rect 14516 19944 16396 19972
rect 14516 19932 14522 19944
rect 16390 19932 16396 19944
rect 16448 19932 16454 19984
rect 16666 19932 16672 19984
rect 16724 19972 16730 19984
rect 17788 19972 17816 20012
rect 16724 19944 17816 19972
rect 16724 19932 16730 19944
rect 18046 19932 18052 19984
rect 18104 19972 18110 19984
rect 18782 19972 18788 19984
rect 18104 19944 18788 19972
rect 18104 19932 18110 19944
rect 18782 19932 18788 19944
rect 18840 19932 18846 19984
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 11072 19876 15485 19904
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 17129 19907 17187 19913
rect 15473 19867 15531 19873
rect 16132 19876 16896 19904
rect 9309 19839 9367 19845
rect 9309 19836 9321 19839
rect 9272 19808 9321 19836
rect 9272 19796 9278 19808
rect 9309 19805 9321 19808
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 11606 19796 11612 19848
rect 11664 19796 11670 19848
rect 13538 19836 13544 19848
rect 13018 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19836 13783 19839
rect 13906 19836 13912 19848
rect 13771 19808 13912 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 13906 19796 13912 19808
rect 13964 19836 13970 19848
rect 14642 19836 14648 19848
rect 13964 19808 14648 19836
rect 13964 19796 13970 19808
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 16132 19845 16160 19876
rect 15381 19839 15439 19845
rect 15381 19836 15393 19839
rect 15252 19808 15393 19836
rect 15252 19796 15258 19808
rect 15381 19805 15393 19808
rect 15427 19805 15439 19839
rect 15381 19799 15439 19805
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16758 19796 16764 19848
rect 16816 19796 16822 19848
rect 16868 19836 16896 19876
rect 17129 19873 17141 19907
rect 17175 19904 17187 19907
rect 17494 19904 17500 19916
rect 17175 19876 17500 19904
rect 17175 19873 17187 19876
rect 17129 19867 17187 19873
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17586 19864 17592 19916
rect 17644 19904 17650 19916
rect 18138 19904 18144 19916
rect 17644 19876 18144 19904
rect 17644 19864 17650 19876
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18690 19904 18696 19916
rect 18371 19876 18696 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18690 19864 18696 19876
rect 18748 19864 18754 19916
rect 19334 19864 19340 19916
rect 19392 19904 19398 19916
rect 19996 19913 20024 20012
rect 20533 20009 20545 20043
rect 20579 20040 20591 20043
rect 20714 20040 20720 20052
rect 20579 20012 20720 20040
rect 20579 20009 20591 20012
rect 20533 20003 20591 20009
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 21348 20043 21406 20049
rect 21348 20009 21360 20043
rect 21394 20040 21406 20043
rect 23566 20040 23572 20052
rect 21394 20012 23572 20040
rect 21394 20009 21406 20012
rect 21348 20003 21406 20009
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 24210 20000 24216 20052
rect 24268 20040 24274 20052
rect 24581 20043 24639 20049
rect 24581 20040 24593 20043
rect 24268 20012 24593 20040
rect 24268 20000 24274 20012
rect 24581 20009 24593 20012
rect 24627 20009 24639 20043
rect 24581 20003 24639 20009
rect 22370 19932 22376 19984
rect 22428 19972 22434 19984
rect 22428 19944 25176 19972
rect 22428 19932 22434 19944
rect 19889 19907 19947 19913
rect 19889 19904 19901 19907
rect 19392 19876 19901 19904
rect 19392 19864 19398 19876
rect 19889 19873 19901 19876
rect 19935 19873 19947 19907
rect 19889 19867 19947 19873
rect 19981 19907 20039 19913
rect 19981 19873 19993 19907
rect 20027 19904 20039 19907
rect 20625 19907 20683 19913
rect 20625 19904 20637 19907
rect 20027 19876 20637 19904
rect 20027 19873 20039 19876
rect 19981 19867 20039 19873
rect 20625 19873 20637 19876
rect 20671 19873 20683 19907
rect 20625 19867 20683 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 23290 19904 23296 19916
rect 21131 19876 23296 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19904 23995 19907
rect 24762 19904 24768 19916
rect 23983 19876 24768 19904
rect 23983 19873 23995 19876
rect 23937 19867 23995 19873
rect 24762 19864 24768 19876
rect 24820 19864 24826 19916
rect 25038 19864 25044 19916
rect 25096 19864 25102 19916
rect 25148 19913 25176 19944
rect 25133 19907 25191 19913
rect 25133 19873 25145 19907
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 18969 19839 19027 19845
rect 18969 19836 18981 19839
rect 16868 19808 18981 19836
rect 18969 19805 18981 19808
rect 19015 19836 19027 19839
rect 20070 19836 20076 19848
rect 19015 19808 20076 19836
rect 19015 19805 19027 19808
rect 18969 19799 19027 19805
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 23382 19796 23388 19848
rect 23440 19836 23446 19848
rect 23753 19839 23811 19845
rect 23753 19836 23765 19839
rect 23440 19808 23765 19836
rect 23440 19796 23446 19808
rect 23753 19805 23765 19808
rect 23799 19805 23811 19839
rect 23753 19799 23811 19805
rect 2038 19728 2044 19780
rect 2096 19768 2102 19780
rect 2961 19771 3019 19777
rect 2961 19768 2973 19771
rect 2096 19740 2973 19768
rect 2096 19728 2102 19740
rect 2961 19737 2973 19740
rect 3007 19737 3019 19771
rect 2961 19731 3019 19737
rect 5997 19771 6055 19777
rect 5997 19737 6009 19771
rect 6043 19768 6055 19771
rect 9490 19768 9496 19780
rect 6043 19740 9496 19768
rect 6043 19737 6055 19740
rect 5997 19731 6055 19737
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 10873 19771 10931 19777
rect 10873 19737 10885 19771
rect 10919 19768 10931 19771
rect 11146 19768 11152 19780
rect 10919 19740 11152 19768
rect 10919 19737 10931 19740
rect 10873 19731 10931 19737
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 11885 19771 11943 19777
rect 11885 19737 11897 19771
rect 11931 19737 11943 19771
rect 14458 19768 14464 19780
rect 11885 19731 11943 19737
rect 13556 19740 14464 19768
rect 4430 19660 4436 19712
rect 4488 19700 4494 19712
rect 6270 19700 6276 19712
rect 4488 19672 6276 19700
rect 4488 19660 4494 19672
rect 6270 19660 6276 19672
rect 6328 19660 6334 19712
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19700 8631 19703
rect 9122 19700 9128 19712
rect 8619 19672 9128 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 9950 19660 9956 19712
rect 10008 19660 10014 19712
rect 10410 19660 10416 19712
rect 10468 19660 10474 19712
rect 11900 19700 11928 19731
rect 13556 19700 13584 19740
rect 14458 19728 14464 19740
rect 14516 19728 14522 19780
rect 14918 19728 14924 19780
rect 14976 19768 14982 19780
rect 14976 19740 15424 19768
rect 14976 19728 14982 19740
rect 11900 19672 13584 19700
rect 13906 19660 13912 19712
rect 13964 19700 13970 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 13964 19672 14289 19700
rect 13964 19660 13970 19672
rect 14277 19669 14289 19672
rect 14323 19669 14335 19703
rect 14277 19663 14335 19669
rect 15286 19660 15292 19712
rect 15344 19660 15350 19712
rect 15396 19700 15424 19740
rect 15470 19728 15476 19780
rect 15528 19768 15534 19780
rect 15528 19740 19472 19768
rect 15528 19728 15534 19740
rect 16666 19700 16672 19712
rect 15396 19672 16672 19700
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 17405 19703 17463 19709
rect 17405 19700 17417 19703
rect 16816 19672 17417 19700
rect 16816 19660 16822 19672
rect 17405 19669 17417 19672
rect 17451 19700 17463 19703
rect 17954 19700 17960 19712
rect 17451 19672 17960 19700
rect 17451 19669 17463 19672
rect 17405 19663 17463 19669
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 18046 19660 18052 19712
rect 18104 19660 18110 19712
rect 18230 19660 18236 19712
rect 18288 19700 18294 19712
rect 18785 19703 18843 19709
rect 18785 19700 18797 19703
rect 18288 19672 18797 19700
rect 18288 19660 18294 19672
rect 18785 19669 18797 19672
rect 18831 19700 18843 19703
rect 18966 19700 18972 19712
rect 18831 19672 18972 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 18966 19660 18972 19672
rect 19024 19660 19030 19712
rect 19334 19660 19340 19712
rect 19392 19660 19398 19712
rect 19444 19709 19472 19740
rect 20714 19728 20720 19780
rect 20772 19768 20778 19780
rect 21358 19768 21364 19780
rect 20772 19740 21364 19768
rect 20772 19728 20778 19740
rect 21358 19728 21364 19740
rect 21416 19768 21422 19780
rect 21416 19740 21850 19768
rect 21416 19728 21422 19740
rect 19429 19703 19487 19709
rect 19429 19669 19441 19703
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 19797 19703 19855 19709
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 20346 19700 20352 19712
rect 19843 19672 20352 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 20346 19660 20352 19672
rect 20404 19660 20410 19712
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 21692 19672 22845 19700
rect 21692 19660 21698 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 22833 19663 22891 19669
rect 23293 19703 23351 19709
rect 23293 19669 23305 19703
rect 23339 19700 23351 19703
rect 23474 19700 23480 19712
rect 23339 19672 23480 19700
rect 23339 19669 23351 19672
rect 23293 19663 23351 19669
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 23661 19703 23719 19709
rect 23661 19669 23673 19703
rect 23707 19700 23719 19703
rect 24118 19700 24124 19712
rect 23707 19672 24124 19700
rect 23707 19669 23719 19672
rect 23661 19663 23719 19669
rect 24118 19660 24124 19672
rect 24176 19660 24182 19712
rect 24394 19660 24400 19712
rect 24452 19700 24458 19712
rect 24949 19703 25007 19709
rect 24949 19700 24961 19703
rect 24452 19672 24961 19700
rect 24452 19660 24458 19672
rect 24949 19669 24961 19672
rect 24995 19669 25007 19703
rect 24949 19663 25007 19669
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 4522 19456 4528 19508
rect 4580 19456 4586 19508
rect 6546 19456 6552 19508
rect 6604 19456 6610 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 8573 19499 8631 19505
rect 8573 19496 8585 19499
rect 6788 19468 8585 19496
rect 6788 19456 6794 19468
rect 8573 19465 8585 19468
rect 8619 19465 8631 19499
rect 8573 19459 8631 19465
rect 9214 19456 9220 19508
rect 9272 19496 9278 19508
rect 10781 19499 10839 19505
rect 10781 19496 10793 19499
rect 9272 19468 10793 19496
rect 9272 19456 9278 19468
rect 10781 19465 10793 19468
rect 10827 19496 10839 19499
rect 10962 19496 10968 19508
rect 10827 19468 10968 19496
rect 10827 19465 10839 19468
rect 10781 19459 10839 19465
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 13814 19496 13820 19508
rect 11664 19468 13820 19496
rect 11664 19456 11670 19468
rect 7742 19428 7748 19440
rect 4080 19400 5396 19428
rect 4080 19369 4108 19400
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19360 2007 19363
rect 4065 19363 4123 19369
rect 1995 19332 3556 19360
rect 1995 19329 2007 19332
rect 1949 19323 2007 19329
rect 1489 19295 1547 19301
rect 1489 19261 1501 19295
rect 1535 19292 1547 19295
rect 1578 19292 1584 19304
rect 1535 19264 1584 19292
rect 1535 19261 1547 19264
rect 1489 19255 1547 19261
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 1854 19252 1860 19304
rect 1912 19292 1918 19304
rect 3528 19301 3556 19332
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4154 19320 4160 19372
rect 4212 19360 4218 19372
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4212 19332 4721 19360
rect 4212 19320 4218 19332
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1912 19264 2237 19292
rect 1912 19252 1918 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 3694 19292 3700 19304
rect 3559 19264 3700 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3694 19252 3700 19264
rect 3752 19252 3758 19304
rect 5166 19252 5172 19304
rect 5224 19252 5230 19304
rect 5368 19292 5396 19400
rect 5460 19400 7748 19428
rect 5460 19369 5488 19400
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 8754 19428 8760 19440
rect 7852 19400 8760 19428
rect 5445 19363 5503 19369
rect 5445 19329 5457 19363
rect 5491 19329 5503 19363
rect 6733 19363 6791 19369
rect 5445 19323 5503 19329
rect 5552 19332 6684 19360
rect 5552 19292 5580 19332
rect 6546 19292 6552 19304
rect 5368 19264 5580 19292
rect 5644 19264 6552 19292
rect 2774 19184 2780 19236
rect 2832 19224 2838 19236
rect 3881 19227 3939 19233
rect 3881 19224 3893 19227
rect 2832 19196 3893 19224
rect 2832 19184 2838 19196
rect 3881 19193 3893 19196
rect 3927 19193 3939 19227
rect 3881 19187 3939 19193
rect 4982 19184 4988 19236
rect 5040 19224 5046 19236
rect 5644 19224 5672 19264
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 6656 19292 6684 19332
rect 6733 19329 6745 19363
rect 6779 19360 6791 19363
rect 7285 19363 7343 19369
rect 6779 19332 6960 19360
rect 6779 19329 6791 19332
rect 6733 19323 6791 19329
rect 6822 19292 6828 19304
rect 6656 19264 6828 19292
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 5040 19196 5672 19224
rect 5040 19184 5046 19196
rect 6270 19184 6276 19236
rect 6328 19224 6334 19236
rect 6932 19224 6960 19332
rect 7285 19329 7297 19363
rect 7331 19360 7343 19363
rect 7852 19360 7880 19400
rect 8754 19388 8760 19400
rect 8812 19388 8818 19440
rect 9306 19388 9312 19440
rect 9364 19388 9370 19440
rect 7331 19332 7880 19360
rect 7929 19363 7987 19369
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7929 19329 7941 19363
rect 7975 19360 7987 19363
rect 8846 19360 8852 19372
rect 7975 19332 8852 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 11149 19363 11207 19369
rect 11149 19360 11161 19363
rect 10442 19332 11161 19360
rect 11149 19329 11161 19332
rect 11195 19360 11207 19363
rect 11609 19363 11667 19369
rect 11609 19360 11621 19363
rect 11195 19332 11621 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11609 19329 11621 19332
rect 11655 19360 11667 19363
rect 11698 19360 11704 19372
rect 11655 19332 11704 19360
rect 11655 19329 11667 19332
rect 11609 19323 11667 19329
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 12158 19320 12164 19372
rect 12216 19360 12222 19372
rect 12728 19369 12756 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14458 19456 14464 19508
rect 14516 19456 14522 19508
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14608 19468 14933 19496
rect 14608 19456 14614 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 14921 19459 14979 19465
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 15470 19496 15476 19508
rect 15335 19468 15476 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 16206 19456 16212 19508
rect 16264 19496 16270 19508
rect 16758 19496 16764 19508
rect 16264 19468 16764 19496
rect 16264 19456 16270 19468
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 17034 19456 17040 19508
rect 17092 19496 17098 19508
rect 18785 19499 18843 19505
rect 17092 19468 18644 19496
rect 17092 19456 17098 19468
rect 14274 19388 14280 19440
rect 14332 19428 14338 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14332 19400 15393 19428
rect 14332 19388 14338 19400
rect 15381 19397 15393 19400
rect 15427 19397 15439 19431
rect 15381 19391 15439 19397
rect 18322 19388 18328 19440
rect 18380 19388 18386 19440
rect 12253 19363 12311 19369
rect 12253 19360 12265 19363
rect 12216 19332 12265 19360
rect 12216 19320 12222 19332
rect 12253 19329 12265 19332
rect 12299 19329 12311 19363
rect 12253 19323 12311 19329
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 14734 19360 14740 19372
rect 14148 19332 14740 19360
rect 14148 19320 14154 19332
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15102 19320 15108 19372
rect 15160 19360 15166 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15160 19332 16129 19360
rect 15160 19320 15166 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16908 19332 17049 19360
rect 16908 19320 16914 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 18616 19360 18644 19468
rect 18785 19465 18797 19499
rect 18831 19465 18843 19499
rect 18785 19459 18843 19465
rect 19245 19499 19303 19505
rect 19245 19465 19257 19499
rect 19291 19496 19303 19499
rect 19518 19496 19524 19508
rect 19291 19468 19524 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 18800 19428 18828 19459
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19659 19468 20453 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 20990 19496 20996 19508
rect 20947 19468 20996 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21174 19456 21180 19508
rect 21232 19496 21238 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21232 19468 22017 19496
rect 21232 19456 21238 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 23382 19456 23388 19508
rect 23440 19456 23446 19508
rect 25041 19499 25099 19505
rect 25041 19465 25053 19499
rect 25087 19496 25099 19499
rect 25130 19496 25136 19508
rect 25087 19468 25136 19496
rect 25087 19465 25099 19468
rect 25041 19459 25099 19465
rect 25130 19456 25136 19468
rect 25188 19496 25194 19508
rect 25682 19496 25688 19508
rect 25188 19468 25688 19496
rect 25188 19456 25194 19468
rect 25682 19456 25688 19468
rect 25740 19456 25746 19508
rect 19886 19428 19892 19440
rect 18800 19400 19892 19428
rect 19886 19388 19892 19400
rect 19944 19388 19950 19440
rect 20070 19388 20076 19440
rect 20128 19428 20134 19440
rect 23400 19428 23428 19456
rect 20128 19400 23428 19428
rect 20128 19388 20134 19400
rect 24026 19388 24032 19440
rect 24084 19388 24090 19440
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 18616 19332 19717 19360
rect 17037 19323 17095 19329
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19978 19320 19984 19372
rect 20036 19360 20042 19372
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20036 19332 20821 19360
rect 20036 19320 20042 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 22094 19360 22100 19372
rect 21140 19332 22100 19360
rect 21140 19320 21146 19332
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 22186 19320 22192 19372
rect 22244 19360 22250 19372
rect 22373 19363 22431 19369
rect 22373 19360 22385 19363
rect 22244 19332 22385 19360
rect 22244 19320 22250 19332
rect 22373 19329 22385 19332
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 8386 19292 8392 19304
rect 7524 19264 8392 19292
rect 7524 19252 7530 19264
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 10962 19252 10968 19304
rect 11020 19292 11026 19304
rect 12526 19292 12532 19304
rect 11020 19264 12532 19292
rect 11020 19252 11026 19264
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 13446 19292 13452 19304
rect 13035 19264 13452 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16022 19292 16028 19304
rect 15611 19264 16028 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 17368 19264 19840 19292
rect 17368 19252 17374 19264
rect 6328 19196 6960 19224
rect 6328 19184 6334 19196
rect 7282 19184 7288 19236
rect 7340 19224 7346 19236
rect 7340 19196 8984 19224
rect 7340 19184 7346 19196
rect 3418 19116 3424 19168
rect 3476 19156 3482 19168
rect 8846 19156 8852 19168
rect 3476 19128 8852 19156
rect 3476 19116 3482 19128
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 8956 19156 8984 19196
rect 10410 19184 10416 19236
rect 10468 19224 10474 19236
rect 10468 19196 12434 19224
rect 10468 19184 10474 19196
rect 9858 19156 9864 19168
rect 8956 19128 9864 19156
rect 9858 19116 9864 19128
rect 9916 19156 9922 19168
rect 10318 19156 10324 19168
rect 9916 19128 10324 19156
rect 9916 19116 9922 19128
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 11330 19116 11336 19168
rect 11388 19116 11394 19168
rect 11698 19116 11704 19168
rect 11756 19116 11762 19168
rect 12066 19116 12072 19168
rect 12124 19116 12130 19168
rect 12406 19156 12434 19196
rect 14090 19184 14096 19236
rect 14148 19224 14154 19236
rect 14734 19224 14740 19236
rect 14148 19196 14740 19224
rect 14148 19184 14154 19196
rect 14734 19184 14740 19196
rect 14792 19224 14798 19236
rect 14918 19224 14924 19236
rect 14792 19196 14924 19224
rect 14792 19184 14798 19196
rect 14918 19184 14924 19196
rect 14976 19184 14982 19236
rect 19812 19224 19840 19264
rect 19886 19252 19892 19304
rect 19944 19252 19950 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 19996 19264 21005 19292
rect 19996 19224 20024 19264
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21358 19252 21364 19304
rect 21416 19292 21422 19304
rect 21545 19295 21603 19301
rect 21545 19292 21557 19295
rect 21416 19264 21557 19292
rect 21416 19252 21422 19264
rect 21545 19261 21557 19264
rect 21591 19261 21603 19295
rect 21545 19255 21603 19261
rect 22002 19252 22008 19304
rect 22060 19292 22066 19304
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 22060 19264 22477 19292
rect 22060 19252 22066 19264
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 25222 19292 25228 19304
rect 23615 19264 25228 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 19812 19196 20024 19224
rect 20162 19184 20168 19236
rect 20220 19224 20226 19236
rect 20220 19196 20392 19224
rect 20220 19184 20226 19196
rect 13722 19156 13728 19168
rect 12406 19128 13728 19156
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 15654 19116 15660 19168
rect 15712 19156 15718 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 15712 19128 16681 19156
rect 15712 19116 15718 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 16669 19119 16727 19125
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 19242 19156 19248 19168
rect 18380 19128 19248 19156
rect 18380 19116 18386 19128
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19978 19156 19984 19168
rect 19484 19128 19984 19156
rect 19484 19116 19490 19128
rect 19978 19116 19984 19128
rect 20036 19156 20042 19168
rect 20257 19159 20315 19165
rect 20257 19156 20269 19159
rect 20036 19128 20269 19156
rect 20036 19116 20042 19128
rect 20257 19125 20269 19128
rect 20303 19125 20315 19159
rect 20364 19156 20392 19196
rect 20806 19184 20812 19236
rect 20864 19224 20870 19236
rect 22572 19224 22600 19255
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 20864 19196 22600 19224
rect 20864 19184 20870 19196
rect 21818 19156 21824 19168
rect 20364 19128 21824 19156
rect 20257 19119 20315 19125
rect 21818 19116 21824 19128
rect 21876 19116 21882 19168
rect 21913 19159 21971 19165
rect 21913 19125 21925 19159
rect 21959 19156 21971 19159
rect 22002 19156 22008 19168
rect 21959 19128 22008 19156
rect 21959 19125 21971 19128
rect 21913 19119 21971 19125
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 25130 19116 25136 19168
rect 25188 19156 25194 19168
rect 25317 19159 25375 19165
rect 25317 19156 25329 19159
rect 25188 19128 25329 19156
rect 25188 19116 25194 19128
rect 25317 19125 25329 19128
rect 25363 19125 25375 19159
rect 25317 19119 25375 19125
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 1765 18955 1823 18961
rect 1765 18921 1777 18955
rect 1811 18952 1823 18955
rect 3878 18952 3884 18964
rect 1811 18924 3884 18952
rect 1811 18921 1823 18924
rect 1765 18915 1823 18921
rect 3878 18912 3884 18924
rect 3936 18912 3942 18964
rect 4065 18955 4123 18961
rect 4065 18921 4077 18955
rect 4111 18952 4123 18955
rect 7282 18952 7288 18964
rect 4111 18924 7288 18952
rect 4111 18921 4123 18924
rect 4065 18915 4123 18921
rect 2406 18844 2412 18896
rect 2464 18884 2470 18896
rect 2464 18856 3924 18884
rect 2464 18844 2470 18856
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 3786 18816 3792 18828
rect 2915 18788 3792 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 3786 18776 3792 18788
rect 3844 18776 3850 18828
rect 3896 18825 3924 18856
rect 3881 18819 3939 18825
rect 3881 18785 3893 18819
rect 3927 18816 3939 18819
rect 4080 18816 4108 18915
rect 7282 18912 7288 18924
rect 7340 18912 7346 18964
rect 14090 18952 14096 18964
rect 7392 18924 12434 18952
rect 4249 18887 4307 18893
rect 4249 18853 4261 18887
rect 4295 18884 4307 18887
rect 4982 18884 4988 18896
rect 4295 18856 4988 18884
rect 4295 18853 4307 18856
rect 4249 18847 4307 18853
rect 4982 18844 4988 18856
rect 5040 18844 5046 18896
rect 5350 18844 5356 18896
rect 5408 18884 5414 18896
rect 7392 18884 7420 18924
rect 5408 18856 7420 18884
rect 5408 18844 5414 18856
rect 7834 18844 7840 18896
rect 7892 18884 7898 18896
rect 10962 18884 10968 18896
rect 7892 18856 10968 18884
rect 7892 18844 7898 18856
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 12406 18884 12434 18924
rect 13556 18924 14096 18952
rect 12989 18887 13047 18893
rect 12989 18884 13001 18887
rect 12406 18856 13001 18884
rect 12989 18853 13001 18856
rect 13035 18853 13047 18887
rect 12989 18847 13047 18853
rect 3927 18788 4108 18816
rect 4801 18819 4859 18825
rect 3927 18785 3939 18788
rect 3881 18779 3939 18785
rect 4801 18785 4813 18819
rect 4847 18816 4859 18819
rect 4890 18816 4896 18828
rect 4847 18788 4896 18816
rect 4847 18785 4859 18788
rect 4801 18779 4859 18785
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 5902 18776 5908 18828
rect 5960 18816 5966 18828
rect 6457 18819 6515 18825
rect 5960 18788 6040 18816
rect 5960 18776 5966 18788
rect 1486 18708 1492 18760
rect 1544 18748 1550 18760
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1544 18720 1685 18748
rect 1544 18708 1550 18720
rect 1673 18717 1685 18720
rect 1719 18748 1731 18751
rect 2133 18751 2191 18757
rect 2133 18748 2145 18751
rect 1719 18720 2145 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 2133 18717 2145 18720
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 2590 18708 2596 18760
rect 2648 18708 2654 18760
rect 6012 18757 6040 18788
rect 6457 18785 6469 18819
rect 6503 18816 6515 18819
rect 6546 18816 6552 18828
rect 6503 18788 6552 18816
rect 6503 18785 6515 18788
rect 6457 18779 6515 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 6733 18819 6791 18825
rect 6733 18785 6745 18819
rect 6779 18816 6791 18819
rect 9398 18816 9404 18828
rect 6779 18788 9404 18816
rect 6779 18785 6791 18788
rect 6733 18779 6791 18785
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 9582 18776 9588 18828
rect 9640 18816 9646 18828
rect 9769 18819 9827 18825
rect 9769 18816 9781 18819
rect 9640 18788 9781 18816
rect 9640 18776 9646 18788
rect 9769 18785 9781 18788
rect 9815 18785 9827 18819
rect 13556 18816 13584 18924
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 15562 18952 15568 18964
rect 14384 18924 15568 18952
rect 14384 18884 14412 18924
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 16758 18912 16764 18964
rect 16816 18952 16822 18964
rect 19613 18955 19671 18961
rect 19613 18952 19625 18955
rect 16816 18924 19625 18952
rect 16816 18912 16822 18924
rect 19613 18921 19625 18924
rect 19659 18921 19671 18955
rect 19613 18915 19671 18921
rect 19720 18924 21680 18952
rect 13648 18856 14412 18884
rect 13648 18825 13676 18856
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 14792 18856 14872 18884
rect 14792 18844 14798 18856
rect 9769 18779 9827 18785
rect 13188 18788 13584 18816
rect 13633 18819 13691 18825
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 5997 18751 6055 18757
rect 5997 18717 6009 18751
rect 6043 18717 6055 18751
rect 5997 18711 6055 18717
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18748 7987 18751
rect 10226 18748 10232 18760
rect 7975 18720 10232 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 2682 18640 2688 18692
rect 2740 18680 2746 18692
rect 4338 18680 4344 18692
rect 2740 18652 4344 18680
rect 2740 18640 2746 18652
rect 4338 18640 4344 18652
rect 4396 18640 4402 18692
rect 4540 18680 4568 18711
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11698 18748 11704 18760
rect 10459 18720 11704 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18748 12587 18751
rect 13188 18748 13216 18788
rect 13633 18785 13645 18819
rect 13679 18785 13691 18819
rect 14458 18816 14464 18828
rect 13633 18779 13691 18785
rect 13740 18788 14464 18816
rect 13740 18748 13768 18788
rect 14458 18776 14464 18788
rect 14516 18776 14522 18828
rect 14844 18825 14872 18856
rect 17218 18844 17224 18896
rect 17276 18844 17282 18896
rect 17586 18844 17592 18896
rect 17644 18844 17650 18896
rect 18049 18887 18107 18893
rect 18049 18853 18061 18887
rect 18095 18884 18107 18887
rect 19058 18884 19064 18896
rect 18095 18856 19064 18884
rect 18095 18853 18107 18856
rect 18049 18847 18107 18853
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 19150 18844 19156 18896
rect 19208 18884 19214 18896
rect 19208 18856 19334 18884
rect 19208 18844 19214 18856
rect 14829 18819 14887 18825
rect 14829 18785 14841 18819
rect 14875 18785 14887 18819
rect 14829 18779 14887 18785
rect 16942 18776 16948 18828
rect 17000 18816 17006 18828
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 17000 18788 18521 18816
rect 17000 18776 17006 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 18598 18776 18604 18828
rect 18656 18776 18662 18828
rect 19306 18816 19334 18856
rect 19720 18816 19748 18924
rect 21652 18884 21680 18924
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 22830 18952 22836 18964
rect 21876 18924 22836 18952
rect 21876 18912 21882 18924
rect 22830 18912 22836 18924
rect 22888 18952 22894 18964
rect 24670 18952 24676 18964
rect 22888 18924 24676 18952
rect 22888 18912 22894 18924
rect 24670 18912 24676 18924
rect 24728 18912 24734 18964
rect 23382 18884 23388 18896
rect 21652 18856 23388 18884
rect 23382 18844 23388 18856
rect 23440 18844 23446 18896
rect 26050 18884 26056 18896
rect 23768 18856 26056 18884
rect 19306 18788 19748 18816
rect 19794 18776 19800 18828
rect 19852 18816 19858 18828
rect 19981 18819 20039 18825
rect 19981 18816 19993 18819
rect 19852 18788 19993 18816
rect 19852 18776 19858 18788
rect 19981 18785 19993 18788
rect 20027 18785 20039 18819
rect 19981 18779 20039 18785
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18816 20683 18819
rect 21634 18816 21640 18828
rect 20671 18788 21640 18816
rect 20671 18785 20683 18788
rect 20625 18779 20683 18785
rect 21634 18776 21640 18788
rect 21692 18776 21698 18828
rect 22462 18776 22468 18828
rect 22520 18816 22526 18828
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22520 18788 23121 18816
rect 22520 18776 22526 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 12575 18720 13216 18748
rect 13280 18720 13768 18748
rect 12575 18717 12587 18720
rect 12529 18711 12587 18717
rect 8294 18680 8300 18692
rect 4540 18652 8300 18680
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 9490 18640 9496 18692
rect 9548 18680 9554 18692
rect 9585 18683 9643 18689
rect 9585 18680 9597 18683
rect 9548 18652 9597 18680
rect 9548 18640 9554 18652
rect 9585 18649 9597 18652
rect 9631 18649 9643 18683
rect 9585 18643 9643 18649
rect 9677 18683 9735 18689
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 13280 18680 13308 18720
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14918 18748 14924 18760
rect 13872 18720 14924 18748
rect 13872 18708 13878 18720
rect 14918 18708 14924 18720
rect 14976 18748 14982 18760
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 14976 18720 15485 18748
rect 14976 18708 14982 18720
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 19300 18720 20361 18748
rect 19300 18708 19306 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 23768 18748 23796 18856
rect 26050 18844 26056 18856
rect 26108 18844 26114 18896
rect 24029 18819 24087 18825
rect 24029 18785 24041 18819
rect 24075 18816 24087 18819
rect 25038 18816 25044 18828
rect 24075 18788 25044 18816
rect 24075 18785 24087 18788
rect 24029 18779 24087 18785
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 25222 18776 25228 18828
rect 25280 18776 25286 18828
rect 25130 18748 25136 18760
rect 20349 18711 20407 18717
rect 22572 18720 23796 18748
rect 23860 18720 25136 18748
rect 9723 18652 13308 18680
rect 13357 18683 13415 18689
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 13906 18680 13912 18692
rect 13403 18652 13912 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13906 18640 13912 18652
rect 13964 18640 13970 18692
rect 14550 18640 14556 18692
rect 14608 18680 14614 18692
rect 14737 18683 14795 18689
rect 14737 18680 14749 18683
rect 14608 18652 14749 18680
rect 14608 18640 14614 18652
rect 14737 18649 14749 18652
rect 14783 18680 14795 18683
rect 15194 18680 15200 18692
rect 14783 18652 15200 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 15194 18640 15200 18652
rect 15252 18680 15258 18692
rect 15654 18680 15660 18692
rect 15252 18652 15660 18680
rect 15252 18640 15258 18652
rect 15654 18640 15660 18652
rect 15712 18640 15718 18692
rect 15749 18683 15807 18689
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 16022 18680 16028 18692
rect 15795 18652 16028 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 16206 18640 16212 18692
rect 16264 18640 16270 18692
rect 17218 18640 17224 18692
rect 17276 18680 17282 18692
rect 19150 18680 19156 18692
rect 17276 18652 19156 18680
rect 17276 18640 17282 18652
rect 19150 18640 19156 18652
rect 19208 18640 19214 18692
rect 19518 18640 19524 18692
rect 19576 18640 19582 18692
rect 20714 18680 20720 18692
rect 19904 18652 20720 18680
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 5350 18612 5356 18624
rect 2188 18584 5356 18612
rect 2188 18572 2194 18584
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 5810 18572 5816 18624
rect 5868 18572 5874 18624
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 7745 18615 7803 18621
rect 7745 18612 7757 18615
rect 5960 18584 7757 18612
rect 5960 18572 5966 18584
rect 7745 18581 7757 18584
rect 7791 18581 7803 18615
rect 7745 18575 7803 18581
rect 8386 18572 8392 18624
rect 8444 18572 8450 18624
rect 8846 18572 8852 18624
rect 8904 18612 8910 18624
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 8904 18584 9229 18612
rect 8904 18572 8910 18584
rect 9217 18581 9229 18584
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 9858 18572 9864 18624
rect 9916 18612 9922 18624
rect 10134 18612 10140 18624
rect 9916 18584 10140 18612
rect 9916 18572 9922 18584
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 12621 18615 12679 18621
rect 12621 18612 12633 18615
rect 12308 18584 12633 18612
rect 12308 18572 12314 18584
rect 12621 18581 12633 18584
rect 12667 18581 12679 18615
rect 12621 18575 12679 18581
rect 13446 18572 13452 18624
rect 13504 18572 13510 18624
rect 14645 18615 14703 18621
rect 14645 18581 14657 18615
rect 14691 18612 14703 18615
rect 15102 18612 15108 18624
rect 14691 18584 15108 18612
rect 14691 18581 14703 18584
rect 14645 18575 14703 18581
rect 15102 18572 15108 18584
rect 15160 18612 15166 18624
rect 17681 18615 17739 18621
rect 17681 18612 17693 18615
rect 15160 18584 17693 18612
rect 15160 18572 15166 18584
rect 17681 18581 17693 18584
rect 17727 18612 17739 18615
rect 17770 18612 17776 18624
rect 17727 18584 17776 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 17770 18572 17776 18584
rect 17828 18572 17834 18624
rect 18417 18615 18475 18621
rect 18417 18581 18429 18615
rect 18463 18612 18475 18615
rect 19904 18612 19932 18652
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 21358 18640 21364 18692
rect 21416 18640 21422 18692
rect 18463 18584 19932 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 20990 18612 20996 18624
rect 20036 18584 20996 18612
rect 20036 18572 20042 18584
rect 20990 18572 20996 18584
rect 21048 18612 21054 18624
rect 21634 18612 21640 18624
rect 21048 18584 21640 18612
rect 21048 18572 21054 18584
rect 21634 18572 21640 18584
rect 21692 18572 21698 18624
rect 22097 18615 22155 18621
rect 22097 18581 22109 18615
rect 22143 18612 22155 18615
rect 22186 18612 22192 18624
rect 22143 18584 22192 18612
rect 22143 18581 22155 18584
rect 22097 18575 22155 18581
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 22572 18621 22600 18720
rect 22830 18640 22836 18692
rect 22888 18680 22894 18692
rect 23017 18683 23075 18689
rect 23017 18680 23029 18683
rect 22888 18652 23029 18680
rect 22888 18640 22894 18652
rect 23017 18649 23029 18652
rect 23063 18649 23075 18683
rect 23017 18643 23075 18649
rect 23198 18640 23204 18692
rect 23256 18680 23262 18692
rect 23860 18689 23888 18720
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 23845 18683 23903 18689
rect 23845 18680 23857 18683
rect 23256 18652 23857 18680
rect 23256 18640 23262 18652
rect 23845 18649 23857 18652
rect 23891 18649 23903 18683
rect 25041 18683 25099 18689
rect 25041 18680 25053 18683
rect 23845 18643 23903 18649
rect 24412 18652 25053 18680
rect 24412 18624 24440 18652
rect 25041 18649 25053 18652
rect 25087 18649 25099 18683
rect 25041 18643 25099 18649
rect 22557 18615 22615 18621
rect 22557 18581 22569 18615
rect 22603 18581 22615 18615
rect 22557 18575 22615 18581
rect 22738 18572 22744 18624
rect 22796 18612 22802 18624
rect 22925 18615 22983 18621
rect 22925 18612 22937 18615
rect 22796 18584 22937 18612
rect 22796 18572 22802 18584
rect 22925 18581 22937 18584
rect 22971 18581 22983 18615
rect 22925 18575 22983 18581
rect 24394 18572 24400 18624
rect 24452 18572 24458 18624
rect 24578 18572 24584 18624
rect 24636 18572 24642 18624
rect 24670 18572 24676 18624
rect 24728 18612 24734 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24728 18584 24961 18612
rect 24728 18572 24734 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18377 2007 18411
rect 1949 18371 2007 18377
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18408 2651 18411
rect 2866 18408 2872 18420
rect 2639 18380 2872 18408
rect 2639 18377 2651 18380
rect 2593 18371 2651 18377
rect 1964 18340 1992 18371
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3881 18411 3939 18417
rect 3881 18377 3893 18411
rect 3927 18408 3939 18411
rect 5626 18408 5632 18420
rect 3927 18380 5632 18408
rect 3927 18377 3939 18380
rect 3881 18371 3939 18377
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 6236 18380 6377 18408
rect 6236 18368 6242 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 6733 18411 6791 18417
rect 6733 18377 6745 18411
rect 6779 18408 6791 18411
rect 7006 18408 7012 18420
rect 6779 18380 7012 18408
rect 6779 18377 6791 18380
rect 6733 18371 6791 18377
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 8294 18368 8300 18420
rect 8352 18368 8358 18420
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 8444 18380 12173 18408
rect 8444 18368 8450 18380
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 13354 18408 13360 18420
rect 12584 18380 13360 18408
rect 12584 18368 12590 18380
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13872 18380 14289 18408
rect 13872 18368 13878 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14516 18380 15209 18408
rect 14516 18368 14522 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 15528 18380 21312 18408
rect 15528 18368 15534 18380
rect 4154 18340 4160 18352
rect 1964 18312 4160 18340
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 9214 18300 9220 18352
rect 9272 18300 9278 18352
rect 10870 18300 10876 18352
rect 10928 18340 10934 18352
rect 10928 18312 15792 18340
rect 10928 18300 10934 18312
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 2038 18272 2044 18284
rect 1719 18244 2044 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 2130 18232 2136 18284
rect 2188 18232 2194 18284
rect 2774 18232 2780 18284
rect 2832 18232 2838 18284
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 3436 18136 3464 18235
rect 4062 18232 4068 18284
rect 4120 18232 4126 18284
rect 4338 18232 4344 18284
rect 4396 18272 4402 18284
rect 5997 18275 6055 18281
rect 5997 18272 6009 18275
rect 4396 18244 6009 18272
rect 4396 18232 4402 18244
rect 5997 18241 6009 18244
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 7193 18275 7251 18281
rect 7193 18241 7205 18275
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 4430 18164 4436 18216
rect 4488 18204 4494 18216
rect 4525 18207 4583 18213
rect 4525 18204 4537 18207
rect 4488 18176 4537 18204
rect 4488 18164 4494 18176
rect 4525 18173 4537 18176
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 4801 18207 4859 18213
rect 4801 18173 4813 18207
rect 4847 18204 4859 18207
rect 6362 18204 6368 18216
rect 4847 18176 6368 18204
rect 4847 18173 4859 18176
rect 4801 18167 4859 18173
rect 6362 18164 6368 18176
rect 6420 18164 6426 18216
rect 7208 18204 7236 18235
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 8478 18232 8484 18284
rect 8536 18232 8542 18284
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 11054 18272 11060 18284
rect 10376 18244 11060 18272
rect 10376 18232 10382 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 11848 18244 13001 18272
rect 11848 18232 11854 18244
rect 12989 18241 13001 18244
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 9766 18204 9772 18216
rect 7208 18176 9772 18204
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 9858 18164 9864 18216
rect 9916 18204 9922 18216
rect 10502 18204 10508 18216
rect 9916 18176 10508 18204
rect 9916 18164 9922 18176
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10962 18164 10968 18216
rect 11020 18204 11026 18216
rect 11241 18207 11299 18213
rect 11241 18204 11253 18207
rect 11020 18176 11253 18204
rect 11020 18164 11026 18176
rect 11241 18173 11253 18176
rect 11287 18204 11299 18207
rect 12253 18207 12311 18213
rect 11287 18176 11928 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 7190 18136 7196 18148
rect 3436 18108 7196 18136
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 7650 18096 7656 18148
rect 7708 18096 7714 18148
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 11793 18139 11851 18145
rect 11793 18136 11805 18139
rect 10284 18108 11805 18136
rect 10284 18096 10290 18108
rect 11793 18105 11805 18108
rect 11839 18105 11851 18139
rect 11793 18099 11851 18105
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 3326 18068 3332 18080
rect 3283 18040 3332 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 5810 18028 5816 18080
rect 5868 18028 5874 18080
rect 7009 18071 7067 18077
rect 7009 18037 7021 18071
rect 7055 18068 7067 18071
rect 9398 18068 9404 18080
rect 7055 18040 9404 18068
rect 7055 18037 7067 18040
rect 7009 18031 7067 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 9824 18040 10701 18068
rect 9824 18028 9830 18040
rect 10689 18037 10701 18040
rect 10735 18068 10747 18071
rect 10870 18068 10876 18080
rect 10735 18040 10876 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11900 18068 11928 18176
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 12268 18136 12296 18167
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 13004 18136 13032 18235
rect 13998 18232 14004 18284
rect 14056 18272 14062 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 14056 18244 15577 18272
rect 14056 18232 14062 18244
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15654 18232 15660 18284
rect 15712 18232 15718 18284
rect 13078 18164 13084 18216
rect 13136 18204 13142 18216
rect 15470 18204 15476 18216
rect 13136 18176 15476 18204
rect 13136 18164 13142 18176
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15764 18213 15792 18312
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 18509 18343 18567 18349
rect 18509 18340 18521 18343
rect 15896 18312 18521 18340
rect 15896 18300 15902 18312
rect 18509 18309 18521 18312
rect 18555 18309 18567 18343
rect 18509 18303 18567 18309
rect 18874 18300 18880 18352
rect 18932 18340 18938 18352
rect 18932 18312 21220 18340
rect 18932 18300 18938 18312
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 16393 18275 16451 18281
rect 16393 18272 16405 18275
rect 16264 18244 16405 18272
rect 16264 18232 16270 18244
rect 16393 18241 16405 18244
rect 16439 18241 16451 18275
rect 16393 18235 16451 18241
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16816 18244 17233 18272
rect 16816 18232 16822 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 17494 18272 17500 18284
rect 17359 18244 17500 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 17494 18232 17500 18244
rect 17552 18272 17558 18284
rect 17552 18244 17908 18272
rect 17552 18232 17558 18244
rect 15749 18207 15807 18213
rect 15749 18173 15761 18207
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 17880 18204 17908 18244
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 18012 18244 18429 18272
rect 18012 18232 18018 18244
rect 18417 18241 18429 18244
rect 18463 18272 18475 18275
rect 19613 18275 19671 18281
rect 18463 18244 19564 18272
rect 18463 18241 18475 18244
rect 18417 18235 18475 18241
rect 18601 18207 18659 18213
rect 17880 18176 18368 18204
rect 16209 18139 16267 18145
rect 16209 18136 16221 18139
rect 12268 18108 12940 18136
rect 13004 18108 16221 18136
rect 12802 18068 12808 18080
rect 11900 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 12912 18068 12940 18108
rect 16209 18105 16221 18108
rect 16255 18136 16267 18139
rect 18230 18136 18236 18148
rect 16255 18108 18236 18136
rect 16255 18105 16267 18108
rect 16209 18099 16267 18105
rect 18230 18096 18236 18108
rect 18288 18096 18294 18148
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 12912 18040 16865 18068
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 17494 18028 17500 18080
rect 17552 18068 17558 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17552 18040 18061 18068
rect 17552 18028 17558 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18340 18068 18368 18176
rect 18601 18173 18613 18207
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 19306 18176 19472 18204
rect 18506 18096 18512 18148
rect 18564 18136 18570 18148
rect 18616 18136 18644 18167
rect 19306 18136 19334 18176
rect 18564 18108 18644 18136
rect 18708 18108 19334 18136
rect 18564 18096 18570 18108
rect 18708 18068 18736 18108
rect 18340 18040 18736 18068
rect 18049 18031 18107 18037
rect 19242 18028 19248 18080
rect 19300 18028 19306 18080
rect 19444 18068 19472 18176
rect 19536 18136 19564 18244
rect 19613 18241 19625 18275
rect 19659 18272 19671 18275
rect 19978 18272 19984 18284
rect 19659 18244 19984 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 19702 18164 19708 18216
rect 19760 18164 19766 18216
rect 19886 18164 19892 18216
rect 19944 18164 19950 18216
rect 20824 18204 20852 18235
rect 20640 18176 20852 18204
rect 20640 18136 20668 18176
rect 20898 18164 20904 18216
rect 20956 18164 20962 18216
rect 21082 18164 21088 18216
rect 21140 18164 21146 18216
rect 21192 18204 21220 18312
rect 21284 18272 21312 18380
rect 21542 18368 21548 18420
rect 21600 18368 21606 18420
rect 21634 18368 21640 18420
rect 21692 18408 21698 18420
rect 22738 18408 22744 18420
rect 21692 18380 22744 18408
rect 21692 18368 21698 18380
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 23290 18408 23296 18420
rect 22848 18380 23296 18408
rect 21560 18340 21588 18368
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21560 18312 22017 18340
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22005 18303 22063 18309
rect 22554 18300 22560 18352
rect 22612 18340 22618 18352
rect 22848 18340 22876 18380
rect 23290 18368 23296 18380
rect 23348 18368 23354 18420
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 24949 18411 25007 18417
rect 24949 18408 24961 18411
rect 23716 18380 24961 18408
rect 23716 18368 23722 18380
rect 24949 18377 24961 18380
rect 24995 18377 25007 18411
rect 24949 18371 25007 18377
rect 22612 18312 22876 18340
rect 22612 18300 22618 18312
rect 22922 18300 22928 18352
rect 22980 18340 22986 18352
rect 25041 18343 25099 18349
rect 25041 18340 25053 18343
rect 22980 18312 25053 18340
rect 22980 18300 22986 18312
rect 25041 18309 25053 18312
rect 25087 18309 25099 18343
rect 25041 18303 25099 18309
rect 23382 18272 23388 18284
rect 21284 18244 23388 18272
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 24394 18204 24400 18216
rect 21192 18176 24400 18204
rect 24394 18164 24400 18176
rect 24452 18164 24458 18216
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25314 18204 25320 18216
rect 25271 18176 25320 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 19536 18108 20668 18136
rect 19978 18068 19984 18080
rect 19444 18040 19984 18068
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 20438 18028 20444 18080
rect 20496 18028 20502 18080
rect 20640 18068 20668 18108
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 24581 18139 24639 18145
rect 24581 18136 24593 18139
rect 20772 18108 24593 18136
rect 20772 18096 20778 18108
rect 24581 18105 24593 18108
rect 24627 18105 24639 18139
rect 24581 18099 24639 18105
rect 21450 18068 21456 18080
rect 20640 18040 21456 18068
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 23382 18028 23388 18080
rect 23440 18068 23446 18080
rect 23750 18068 23756 18080
rect 23440 18040 23756 18068
rect 23440 18028 23446 18040
rect 23750 18028 23756 18040
rect 23808 18028 23814 18080
rect 24026 18028 24032 18080
rect 24084 18028 24090 18080
rect 24210 18028 24216 18080
rect 24268 18028 24274 18080
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25866 18068 25872 18080
rect 25096 18040 25872 18068
rect 25096 18028 25102 18040
rect 25866 18028 25872 18040
rect 25924 18028 25930 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 4062 17864 4068 17876
rect 3927 17836 4068 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 4249 17867 4307 17873
rect 4249 17833 4261 17867
rect 4295 17864 4307 17867
rect 4430 17864 4436 17876
rect 4295 17836 4436 17864
rect 4295 17833 4307 17836
rect 4249 17827 4307 17833
rect 4430 17824 4436 17836
rect 4488 17824 4494 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 5592 17836 6469 17864
rect 5592 17824 5598 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 6457 17827 6515 17833
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7156 17836 7757 17864
rect 7156 17824 7162 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 7745 17827 7803 17833
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 8570 17864 8576 17876
rect 8444 17836 8576 17864
rect 8444 17824 8450 17836
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 8662 17824 8668 17876
rect 8720 17864 8726 17876
rect 13998 17864 14004 17876
rect 8720 17836 14004 17864
rect 8720 17824 8726 17836
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 17129 17867 17187 17873
rect 17129 17864 17141 17867
rect 15028 17836 17141 17864
rect 5350 17756 5356 17808
rect 5408 17796 5414 17808
rect 9125 17799 9183 17805
rect 9125 17796 9137 17799
rect 5408 17768 9137 17796
rect 5408 17756 5414 17768
rect 9125 17765 9137 17768
rect 9171 17765 9183 17799
rect 9125 17759 9183 17765
rect 13446 17756 13452 17808
rect 13504 17796 13510 17808
rect 15028 17796 15056 17836
rect 17129 17833 17141 17836
rect 17175 17833 17187 17867
rect 17129 17827 17187 17833
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 17862 17864 17868 17876
rect 17644 17836 17868 17864
rect 17644 17824 17650 17836
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 20980 17867 21038 17873
rect 20980 17833 20992 17867
rect 21026 17864 21038 17867
rect 22186 17864 22192 17876
rect 21026 17836 22192 17864
rect 21026 17833 21038 17836
rect 20980 17827 21038 17833
rect 22186 17824 22192 17836
rect 22244 17824 22250 17876
rect 22465 17867 22523 17873
rect 22465 17833 22477 17867
rect 22511 17864 22523 17867
rect 22646 17864 22652 17876
rect 22511 17836 22652 17864
rect 22511 17833 22523 17836
rect 22465 17827 22523 17833
rect 22646 17824 22652 17836
rect 22704 17824 22710 17876
rect 23014 17824 23020 17876
rect 23072 17864 23078 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 23072 17836 23305 17864
rect 23072 17824 23078 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 24581 17867 24639 17873
rect 24581 17833 24593 17867
rect 24627 17864 24639 17867
rect 24946 17864 24952 17876
rect 24627 17836 24952 17864
rect 24627 17833 24639 17836
rect 24581 17827 24639 17833
rect 24946 17824 24952 17836
rect 25004 17824 25010 17876
rect 18693 17799 18751 17805
rect 18693 17796 18705 17799
rect 13504 17768 15056 17796
rect 16224 17768 18705 17796
rect 13504 17756 13510 17768
rect 1946 17688 1952 17740
rect 2004 17688 2010 17740
rect 5074 17728 5080 17740
rect 3436 17700 5080 17728
rect 3436 17669 3464 17700
rect 5074 17688 5080 17700
rect 5132 17688 5138 17740
rect 5442 17688 5448 17740
rect 5500 17688 5506 17740
rect 8938 17688 8944 17740
rect 8996 17728 9002 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 8996 17700 9781 17728
rect 8996 17688 9002 17700
rect 9769 17697 9781 17700
rect 9815 17728 9827 17731
rect 11698 17728 11704 17740
rect 9815 17700 11704 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11756 17700 11989 17728
rect 11756 17688 11762 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12618 17728 12624 17740
rect 12299 17700 12624 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 14918 17688 14924 17740
rect 14976 17688 14982 17740
rect 15197 17731 15255 17737
rect 15197 17697 15209 17731
rect 15243 17728 15255 17731
rect 15562 17728 15568 17740
rect 15243 17700 15568 17728
rect 15243 17697 15255 17700
rect 15197 17691 15255 17697
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 15930 17688 15936 17740
rect 15988 17728 15994 17740
rect 16224 17728 16252 17768
rect 18693 17765 18705 17768
rect 18739 17765 18751 17799
rect 24118 17796 24124 17808
rect 18693 17759 18751 17765
rect 22848 17768 24124 17796
rect 15988 17700 16252 17728
rect 15988 17688 15994 17700
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 16724 17700 17693 17728
rect 16724 17688 16730 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 20070 17688 20076 17740
rect 20128 17688 20134 17740
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 22554 17728 22560 17740
rect 20763 17700 22560 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 22554 17688 22560 17700
rect 22612 17688 22618 17740
rect 22848 17728 22876 17768
rect 24118 17756 24124 17768
rect 24176 17756 24182 17808
rect 22664 17700 22876 17728
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17629 2835 17663
rect 2777 17623 2835 17629
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17629 3479 17663
rect 3421 17623 3479 17629
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17660 4123 17663
rect 4709 17663 4767 17669
rect 4709 17660 4721 17663
rect 4111 17632 4721 17660
rect 4111 17629 4123 17632
rect 4065 17623 4123 17629
rect 4709 17629 4721 17632
rect 4755 17660 4767 17663
rect 4798 17660 4804 17672
rect 4755 17632 4804 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 2792 17592 2820 17623
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 4982 17620 4988 17672
rect 5040 17660 5046 17672
rect 5169 17663 5227 17669
rect 5169 17660 5181 17663
rect 5040 17632 5181 17660
rect 5040 17620 5046 17632
rect 5169 17629 5181 17632
rect 5215 17629 5227 17663
rect 5169 17623 5227 17629
rect 6638 17620 6644 17672
rect 6696 17620 6702 17672
rect 7006 17620 7012 17672
rect 7064 17660 7070 17672
rect 7285 17663 7343 17669
rect 7285 17660 7297 17663
rect 7064 17632 7297 17660
rect 7064 17620 7070 17632
rect 7285 17629 7297 17632
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7524 17632 7941 17660
rect 7524 17620 7530 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17660 9367 17663
rect 9674 17660 9680 17672
rect 9355 17632 9680 17660
rect 9355 17629 9367 17632
rect 9309 17623 9367 17629
rect 6730 17592 6736 17604
rect 2792 17564 6736 17592
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 2593 17527 2651 17533
rect 2593 17493 2605 17527
rect 2639 17524 2651 17527
rect 2682 17524 2688 17536
rect 2639 17496 2688 17524
rect 2639 17493 2651 17496
rect 2593 17487 2651 17493
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 3234 17484 3240 17536
rect 3292 17484 3298 17536
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17524 4583 17527
rect 5442 17524 5448 17536
rect 4571 17496 5448 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 7098 17484 7104 17536
rect 7156 17484 7162 17536
rect 8386 17484 8392 17536
rect 8444 17484 8450 17536
rect 8588 17524 8616 17623
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 17402 17660 17408 17672
rect 16500 17632 17408 17660
rect 9582 17552 9588 17604
rect 9640 17592 9646 17604
rect 10042 17592 10048 17604
rect 9640 17564 10048 17592
rect 9640 17552 9646 17564
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 10318 17592 10324 17604
rect 10192 17564 10324 17592
rect 10192 17552 10198 17564
rect 10318 17552 10324 17564
rect 10376 17592 10382 17604
rect 10376 17564 10534 17592
rect 10376 17552 10382 17564
rect 12250 17552 12256 17604
rect 12308 17592 12314 17604
rect 12710 17592 12716 17604
rect 12308 17564 12716 17592
rect 12308 17552 12314 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 13740 17564 14583 17592
rect 11330 17524 11336 17536
rect 8588 17496 11336 17524
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 11517 17527 11575 17533
rect 11517 17493 11529 17527
rect 11563 17524 11575 17527
rect 12434 17524 12440 17536
rect 11563 17496 12440 17524
rect 11563 17493 11575 17496
rect 11517 17487 11575 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 13740 17533 13768 17564
rect 13725 17527 13783 17533
rect 13725 17524 13737 17527
rect 12584 17496 13737 17524
rect 12584 17484 12590 17496
rect 13725 17493 13737 17496
rect 13771 17493 13783 17527
rect 13725 17487 13783 17493
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14277 17527 14335 17533
rect 14277 17524 14289 17527
rect 14056 17496 14289 17524
rect 14056 17484 14062 17496
rect 14277 17493 14289 17496
rect 14323 17493 14335 17527
rect 14555 17524 14583 17564
rect 15102 17552 15108 17604
rect 15160 17592 15166 17604
rect 15470 17592 15476 17604
rect 15160 17564 15476 17592
rect 15160 17552 15166 17564
rect 15470 17552 15476 17564
rect 15528 17552 15534 17604
rect 15654 17552 15660 17604
rect 15712 17552 15718 17604
rect 16500 17524 16528 17632
rect 17402 17620 17408 17632
rect 17460 17620 17466 17672
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 17644 17632 19901 17660
rect 17644 17620 17650 17632
rect 19889 17629 19901 17632
rect 19935 17629 19947 17663
rect 19889 17623 19947 17629
rect 17034 17552 17040 17604
rect 17092 17592 17098 17604
rect 17497 17595 17555 17601
rect 17497 17592 17509 17595
rect 17092 17564 17509 17592
rect 17092 17552 17098 17564
rect 17497 17561 17509 17564
rect 17543 17561 17555 17595
rect 17497 17555 17555 17561
rect 17678 17552 17684 17604
rect 17736 17592 17742 17604
rect 18509 17595 18567 17601
rect 18509 17592 18521 17595
rect 17736 17564 18521 17592
rect 17736 17552 17742 17564
rect 18509 17561 18521 17564
rect 18555 17561 18567 17595
rect 18509 17555 18567 17561
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 18969 17595 19027 17601
rect 18969 17592 18981 17595
rect 18656 17564 18981 17592
rect 18656 17552 18662 17564
rect 18969 17561 18981 17564
rect 19015 17561 19027 17595
rect 18969 17555 19027 17561
rect 19797 17595 19855 17601
rect 19797 17561 19809 17595
rect 19843 17592 19855 17595
rect 19843 17564 20944 17592
rect 19843 17561 19855 17564
rect 19797 17555 19855 17561
rect 14555 17496 16528 17524
rect 16669 17527 16727 17533
rect 14277 17487 14335 17493
rect 16669 17493 16681 17527
rect 16715 17524 16727 17527
rect 17310 17524 17316 17536
rect 16715 17496 17316 17524
rect 16715 17493 16727 17496
rect 16669 17487 16727 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 17589 17527 17647 17533
rect 17589 17493 17601 17527
rect 17635 17524 17647 17527
rect 17770 17524 17776 17536
rect 17635 17496 17776 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 18230 17484 18236 17536
rect 18288 17524 18294 17536
rect 18874 17524 18880 17536
rect 18288 17496 18880 17524
rect 18288 17484 18294 17496
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19702 17524 19708 17536
rect 19475 17496 19708 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 20916 17524 20944 17564
rect 21634 17552 21640 17604
rect 21692 17552 21698 17604
rect 22664 17524 22692 17700
rect 22922 17688 22928 17740
rect 22980 17728 22986 17740
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 22980 17700 23029 17728
rect 22980 17688 22986 17700
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 23017 17691 23075 17697
rect 23566 17688 23572 17740
rect 23624 17728 23630 17740
rect 23845 17731 23903 17737
rect 23845 17728 23857 17731
rect 23624 17700 23857 17728
rect 23624 17688 23630 17700
rect 23845 17697 23857 17700
rect 23891 17697 23903 17731
rect 23845 17691 23903 17697
rect 25225 17731 25283 17737
rect 25225 17697 25237 17731
rect 25271 17728 25283 17731
rect 25590 17728 25596 17740
rect 25271 17700 25596 17728
rect 25271 17697 25283 17700
rect 25225 17691 25283 17697
rect 25590 17688 25596 17700
rect 25648 17688 25654 17740
rect 22830 17620 22836 17672
rect 22888 17660 22894 17672
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 22888 17632 23673 17660
rect 22888 17620 22894 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 23934 17660 23940 17672
rect 23799 17632 23940 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 23934 17620 23940 17632
rect 23992 17620 23998 17672
rect 22738 17552 22744 17604
rect 22796 17592 22802 17604
rect 25041 17595 25099 17601
rect 25041 17592 25053 17595
rect 22796 17564 25053 17592
rect 22796 17552 22802 17564
rect 25041 17561 25053 17564
rect 25087 17561 25099 17595
rect 25041 17555 25099 17561
rect 20916 17496 22692 17524
rect 22833 17527 22891 17533
rect 22833 17493 22845 17527
rect 22879 17524 22891 17527
rect 22922 17524 22928 17536
rect 22879 17496 22928 17524
rect 22879 17493 22891 17496
rect 22833 17487 22891 17493
rect 22922 17484 22928 17496
rect 22980 17484 22986 17536
rect 23750 17484 23756 17536
rect 23808 17524 23814 17536
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 23808 17496 24409 17524
rect 23808 17484 23814 17496
rect 24397 17493 24409 17496
rect 24443 17524 24455 17527
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24443 17496 24961 17524
rect 24443 17493 24455 17496
rect 24397 17487 24455 17493
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 1762 17320 1768 17332
rect 1627 17292 1768 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 2593 17323 2651 17329
rect 2593 17289 2605 17323
rect 2639 17320 2651 17323
rect 6546 17320 6552 17332
rect 2639 17292 6552 17320
rect 2639 17289 2651 17292
rect 2593 17283 2651 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 7193 17323 7251 17329
rect 7193 17289 7205 17323
rect 7239 17320 7251 17323
rect 7282 17320 7288 17332
rect 7239 17292 7288 17320
rect 7239 17289 7251 17292
rect 7193 17283 7251 17289
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7432 17292 7849 17320
rect 7432 17280 7438 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 8444 17292 15853 17320
rect 8444 17280 8450 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 15930 17280 15936 17332
rect 15988 17320 15994 17332
rect 17586 17320 17592 17332
rect 15988 17292 17592 17320
rect 15988 17280 15994 17292
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 17770 17280 17776 17332
rect 17828 17320 17834 17332
rect 17865 17323 17923 17329
rect 17865 17320 17877 17323
rect 17828 17292 17877 17320
rect 17828 17280 17834 17292
rect 17865 17289 17877 17292
rect 17911 17289 17923 17323
rect 17865 17283 17923 17289
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 20073 17323 20131 17329
rect 20073 17320 20085 17323
rect 19392 17292 20085 17320
rect 19392 17280 19398 17292
rect 20073 17289 20085 17292
rect 20119 17320 20131 17323
rect 20254 17320 20260 17332
rect 20119 17292 20260 17320
rect 20119 17289 20131 17292
rect 20073 17283 20131 17289
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 22278 17280 22284 17332
rect 22336 17280 22342 17332
rect 22370 17280 22376 17332
rect 22428 17320 22434 17332
rect 23014 17320 23020 17332
rect 22428 17292 23020 17320
rect 22428 17280 22434 17292
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 23658 17320 23664 17332
rect 23216 17292 23664 17320
rect 2317 17255 2375 17261
rect 2317 17221 2329 17255
rect 2363 17252 2375 17255
rect 3602 17252 3608 17264
rect 2363 17224 3608 17252
rect 2363 17221 2375 17224
rect 2317 17215 2375 17221
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2130 17184 2136 17196
rect 1811 17156 2136 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2792 17193 2820 17224
rect 3602 17212 3608 17224
rect 3660 17212 3666 17264
rect 7558 17252 7564 17264
rect 4816 17224 7564 17252
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 3237 17187 3295 17193
rect 2823 17156 2857 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 3237 17153 3249 17187
rect 3283 17184 3295 17187
rect 3326 17184 3332 17196
rect 3283 17156 3332 17184
rect 3283 17153 3295 17156
rect 3237 17147 3295 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17184 3571 17187
rect 4614 17184 4620 17196
rect 3559 17156 4620 17184
rect 3559 17153 3571 17156
rect 3513 17147 3571 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 4816 17193 4844 17224
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 7650 17212 7656 17264
rect 7708 17252 7714 17264
rect 8478 17252 8484 17264
rect 7708 17224 8484 17252
rect 7708 17212 7714 17224
rect 8478 17212 8484 17224
rect 8536 17212 8542 17264
rect 9493 17255 9551 17261
rect 9493 17221 9505 17255
rect 9539 17252 9551 17255
rect 9766 17252 9772 17264
rect 9539 17224 9772 17252
rect 9539 17221 9551 17224
rect 9493 17215 9551 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 10134 17212 10140 17264
rect 10192 17212 10198 17264
rect 12250 17252 12256 17264
rect 11256 17224 12256 17252
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17184 6055 17187
rect 6178 17184 6184 17196
rect 6043 17156 6184 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 6914 17184 6920 17196
rect 6779 17156 6920 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7374 17144 7380 17196
rect 7432 17144 7438 17196
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 7926 17184 7932 17196
rect 7800 17156 7932 17184
rect 7800 17144 7806 17156
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 4525 17119 4583 17125
rect 4525 17116 4537 17119
rect 4212 17088 4537 17116
rect 4212 17076 4218 17088
rect 4525 17085 4537 17088
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 8036 17116 8064 17147
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8996 17156 9229 17184
rect 8996 17144 9002 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11256 17193 11284 17224
rect 12250 17212 12256 17224
rect 12308 17252 12314 17264
rect 12308 17224 12466 17252
rect 12308 17212 12314 17224
rect 13446 17212 13452 17264
rect 13504 17252 13510 17264
rect 17678 17252 17684 17264
rect 13504 17224 17684 17252
rect 13504 17212 13510 17224
rect 17678 17212 17684 17224
rect 17736 17212 17742 17264
rect 18598 17212 18604 17264
rect 18656 17252 18662 17264
rect 18656 17224 19090 17252
rect 18656 17212 18662 17224
rect 22094 17212 22100 17264
rect 22152 17252 22158 17264
rect 22830 17252 22836 17264
rect 22152 17224 22836 17252
rect 22152 17212 22158 17224
rect 22830 17212 22836 17224
rect 22888 17212 22894 17264
rect 22922 17212 22928 17264
rect 22980 17252 22986 17264
rect 23216 17252 23244 17292
rect 23658 17280 23664 17292
rect 23716 17320 23722 17332
rect 23716 17292 23980 17320
rect 23716 17280 23722 17292
rect 22980 17224 23322 17252
rect 22980 17212 22986 17224
rect 11241 17187 11299 17193
rect 11241 17184 11253 17187
rect 11112 17156 11253 17184
rect 11112 17144 11118 17156
rect 11241 17153 11253 17156
rect 11287 17153 11299 17187
rect 11241 17147 11299 17153
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17184 14427 17187
rect 15286 17184 15292 17196
rect 14415 17156 15292 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 15286 17144 15292 17156
rect 15344 17184 15350 17196
rect 15344 17156 16896 17184
rect 15344 17144 15350 17156
rect 5592 17088 8064 17116
rect 5592 17076 5598 17088
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10100 17088 10977 17116
rect 10100 17076 10106 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 11977 17119 12035 17125
rect 11977 17085 11989 17119
rect 12023 17116 12035 17119
rect 12434 17116 12440 17128
rect 12023 17088 12440 17116
rect 12023 17085 12035 17088
rect 11977 17079 12035 17085
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 12676 17088 13461 17116
rect 12676 17076 12682 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14148 17088 15148 17116
rect 14148 17076 14154 17088
rect 5813 17051 5871 17057
rect 5813 17017 5825 17051
rect 5859 17048 5871 17051
rect 8294 17048 8300 17060
rect 5859 17020 8300 17048
rect 5859 17017 5871 17020
rect 5813 17011 5871 17017
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 8573 17051 8631 17057
rect 8573 17017 8585 17051
rect 8619 17048 8631 17051
rect 8662 17048 8668 17060
rect 8619 17020 8668 17048
rect 8619 17017 8631 17020
rect 8573 17011 8631 17017
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 11146 17008 11152 17060
rect 11204 17048 11210 17060
rect 15013 17051 15071 17057
rect 15013 17048 15025 17051
rect 11204 17020 11744 17048
rect 11204 17008 11210 17020
rect 6546 16940 6552 16992
rect 6604 16940 6610 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 11606 16980 11612 16992
rect 7432 16952 11612 16980
rect 7432 16940 7438 16952
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 11716 16980 11744 17020
rect 13004 17020 15025 17048
rect 13004 16980 13032 17020
rect 15013 17017 15025 17020
rect 15059 17017 15071 17051
rect 15120 17048 15148 17088
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 15528 17088 15945 17116
rect 15528 17076 15534 17088
rect 15933 17085 15945 17088
rect 15979 17085 15991 17119
rect 15933 17079 15991 17085
rect 16025 17119 16083 17125
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16868 17116 16896 17156
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17000 17156 17233 17184
rect 17000 17144 17006 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 17862 17184 17868 17196
rect 17359 17156 17868 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 20533 17187 20591 17193
rect 20533 17153 20545 17187
rect 20579 17184 20591 17187
rect 22278 17184 22284 17196
rect 20579 17156 22284 17184
rect 20579 17153 20591 17156
rect 20533 17147 20591 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 22554 17144 22560 17196
rect 22612 17144 22618 17196
rect 23952 17184 23980 17292
rect 24118 17280 24124 17332
rect 24176 17320 24182 17332
rect 24176 17292 24900 17320
rect 24176 17280 24182 17292
rect 24872 17261 24900 17292
rect 24857 17255 24915 17261
rect 24857 17221 24869 17255
rect 24903 17221 24915 17255
rect 24857 17215 24915 17221
rect 24210 17184 24216 17196
rect 23952 17170 24216 17184
rect 23966 17156 24216 17170
rect 24210 17144 24216 17156
rect 24268 17184 24274 17196
rect 25317 17187 25375 17193
rect 25317 17184 25329 17187
rect 24268 17156 25329 17184
rect 24268 17144 24274 17156
rect 25317 17153 25329 17156
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 16868 17088 16988 17116
rect 16025 17079 16083 17085
rect 16040 17048 16068 17079
rect 15120 17020 16068 17048
rect 15013 17011 15071 17017
rect 11716 16952 13032 16980
rect 13722 16940 13728 16992
rect 13780 16940 13786 16992
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16980 14151 16983
rect 14274 16980 14280 16992
rect 14139 16952 14280 16980
rect 14139 16949 14151 16952
rect 14093 16943 14151 16949
rect 14274 16940 14280 16952
rect 14332 16980 14338 16992
rect 14734 16980 14740 16992
rect 14332 16952 14740 16980
rect 14332 16940 14338 16952
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 15160 16952 15485 16980
rect 15160 16940 15166 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 16850 16940 16856 16992
rect 16908 16940 16914 16992
rect 16960 16980 16988 17088
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 18601 17119 18659 17125
rect 18601 17085 18613 17119
rect 18647 17116 18659 17119
rect 19150 17116 19156 17128
rect 18647 17088 19156 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 19610 17076 19616 17128
rect 19668 17116 19674 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 19668 17088 21189 17116
rect 19668 17076 19674 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21358 17076 21364 17128
rect 21416 17116 21422 17128
rect 21545 17119 21603 17125
rect 21545 17116 21557 17119
rect 21416 17088 21557 17116
rect 21416 17076 21422 17088
rect 21545 17085 21557 17088
rect 21591 17116 21603 17119
rect 21634 17116 21640 17128
rect 21591 17088 21640 17116
rect 21591 17085 21603 17088
rect 21545 17079 21603 17085
rect 21634 17076 21640 17088
rect 21692 17116 21698 17128
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21692 17088 21925 17116
rect 21692 17076 21698 17088
rect 21913 17085 21925 17088
rect 21959 17116 21971 17119
rect 22097 17119 22155 17125
rect 22097 17116 22109 17119
rect 21959 17088 22109 17116
rect 21959 17085 21971 17088
rect 21913 17079 21971 17085
rect 22097 17085 22109 17088
rect 22143 17116 22155 17119
rect 22922 17116 22928 17128
rect 22143 17088 22928 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 22922 17076 22928 17088
rect 22980 17076 22986 17128
rect 23566 17076 23572 17128
rect 23624 17116 23630 17128
rect 24305 17119 24363 17125
rect 24305 17116 24317 17119
rect 23624 17088 24317 17116
rect 23624 17076 23630 17088
rect 24305 17085 24317 17088
rect 24351 17085 24363 17119
rect 25682 17116 25688 17128
rect 24305 17079 24363 17085
rect 24964 17088 25688 17116
rect 20622 17048 20628 17060
rect 19996 17020 20628 17048
rect 19996 16980 20024 17020
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 24118 17008 24124 17060
rect 24176 17048 24182 17060
rect 24486 17048 24492 17060
rect 24176 17020 24492 17048
rect 24176 17008 24182 17020
rect 24486 17008 24492 17020
rect 24544 17008 24550 17060
rect 16960 16952 20024 16980
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20806 16980 20812 16992
rect 20220 16952 20812 16980
rect 20220 16940 20226 16952
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 22820 16983 22878 16989
rect 22820 16949 22832 16983
rect 22866 16980 22878 16983
rect 24964 16980 24992 17088
rect 25682 17076 25688 17088
rect 25740 17076 25746 17128
rect 25041 17051 25099 17057
rect 25041 17017 25053 17051
rect 25087 17048 25099 17051
rect 26510 17048 26516 17060
rect 25087 17020 26516 17048
rect 25087 17017 25099 17020
rect 25041 17011 25099 17017
rect 26510 17008 26516 17020
rect 26568 17008 26574 17060
rect 22866 16952 24992 16980
rect 22866 16949 22878 16952
rect 22820 16943 22878 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 5813 16779 5871 16785
rect 5813 16745 5825 16779
rect 5859 16776 5871 16779
rect 6638 16776 6644 16788
rect 5859 16748 6644 16776
rect 5859 16745 5871 16748
rect 5813 16739 5871 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 7282 16736 7288 16788
rect 7340 16736 7346 16788
rect 7745 16779 7803 16785
rect 7745 16745 7757 16779
rect 7791 16776 7803 16779
rect 7791 16748 7880 16776
rect 7791 16745 7803 16748
rect 7745 16739 7803 16745
rect 5902 16708 5908 16720
rect 4540 16680 5908 16708
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 2547 16612 2774 16640
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 2746 16584 2774 16612
rect 3878 16600 3884 16652
rect 3936 16600 3942 16652
rect 4540 16649 4568 16680
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 6549 16711 6607 16717
rect 6549 16677 6561 16711
rect 6595 16708 6607 16711
rect 7466 16708 7472 16720
rect 6595 16680 7472 16708
rect 6595 16677 6607 16680
rect 6549 16671 6607 16677
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 7650 16708 7656 16720
rect 7576 16680 7656 16708
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16609 4583 16643
rect 4525 16603 4583 16609
rect 4706 16600 4712 16652
rect 4764 16640 4770 16652
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4764 16612 4813 16640
rect 4764 16600 4770 16612
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 7576 16640 7604 16680
rect 7650 16668 7656 16680
rect 7708 16668 7714 16720
rect 7852 16708 7880 16748
rect 9030 16736 9036 16788
rect 9088 16736 9094 16788
rect 9217 16779 9275 16785
rect 9217 16745 9229 16779
rect 9263 16776 9275 16779
rect 9950 16776 9956 16788
rect 9263 16748 9956 16776
rect 9263 16745 9275 16748
rect 9217 16739 9275 16745
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 15102 16776 15108 16788
rect 10060 16748 11008 16776
rect 8294 16708 8300 16720
rect 7852 16680 8300 16708
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 8389 16711 8447 16717
rect 8389 16677 8401 16711
rect 8435 16677 8447 16711
rect 8389 16671 8447 16677
rect 7147 16612 7604 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 2746 16544 2780 16584
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 3896 16572 3924 16600
rect 8404 16584 8432 16671
rect 9490 16668 9496 16720
rect 9548 16668 9554 16720
rect 10060 16708 10088 16748
rect 10318 16708 10324 16720
rect 9600 16680 10088 16708
rect 10152 16680 10324 16708
rect 3467 16544 3924 16572
rect 5997 16575 6055 16581
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 5997 16541 6009 16575
rect 6043 16541 6055 16575
rect 5997 16535 6055 16541
rect 4154 16504 4160 16516
rect 2608 16476 4160 16504
rect 1946 16396 1952 16448
rect 2004 16396 2010 16448
rect 2608 16445 2636 16476
rect 4154 16464 4160 16476
rect 4212 16464 4218 16516
rect 6012 16504 6040 16535
rect 6730 16532 6736 16584
rect 6788 16532 6794 16584
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16572 7527 16575
rect 7558 16572 7564 16584
rect 7515 16544 7564 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 7926 16532 7932 16584
rect 7984 16532 7990 16584
rect 8386 16532 8392 16584
rect 8444 16532 8450 16584
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 8662 16572 8668 16584
rect 8619 16544 8668 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8662 16532 8668 16544
rect 8720 16532 8726 16584
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 9600 16572 9628 16680
rect 10152 16649 10180 16680
rect 10318 16668 10324 16680
rect 10376 16668 10382 16720
rect 10594 16668 10600 16720
rect 10652 16708 10658 16720
rect 10781 16711 10839 16717
rect 10781 16708 10793 16711
rect 10652 16680 10793 16708
rect 10652 16668 10658 16680
rect 10781 16677 10793 16680
rect 10827 16677 10839 16711
rect 10781 16671 10839 16677
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16609 10195 16643
rect 10980 16640 11008 16748
rect 11256 16748 15108 16776
rect 11256 16649 11284 16748
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 19518 16776 19524 16788
rect 16132 16748 19524 16776
rect 15654 16668 15660 16720
rect 15712 16708 15718 16720
rect 16132 16708 16160 16748
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 19692 16779 19750 16785
rect 19692 16745 19704 16779
rect 19738 16776 19750 16779
rect 20162 16776 20168 16788
rect 19738 16748 20168 16776
rect 19738 16745 19750 16748
rect 19692 16739 19750 16745
rect 20162 16736 20168 16748
rect 20220 16736 20226 16788
rect 20346 16736 20352 16788
rect 20404 16776 20410 16788
rect 21450 16776 21456 16788
rect 20404 16748 21456 16776
rect 20404 16736 20410 16748
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 15712 16680 16160 16708
rect 15712 16668 15718 16680
rect 11241 16643 11299 16649
rect 10980 16612 11100 16640
rect 10137 16603 10195 16609
rect 8904 16544 9628 16572
rect 9677 16575 9735 16581
rect 8904 16532 8910 16544
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 10962 16572 10968 16584
rect 9723 16544 10968 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11072 16572 11100 16612
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11425 16643 11483 16649
rect 11425 16609 11437 16643
rect 11471 16640 11483 16643
rect 11606 16640 11612 16652
rect 11471 16612 11612 16640
rect 11471 16609 11483 16612
rect 11425 16603 11483 16609
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 12710 16600 12716 16652
rect 12768 16640 12774 16652
rect 13722 16640 13728 16652
rect 12768 16612 13728 16640
rect 12768 16600 12774 16612
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14918 16640 14924 16652
rect 14323 16612 14924 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 17405 16643 17463 16649
rect 15804 16612 17080 16640
rect 15804 16600 15810 16612
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 11072 16544 11161 16572
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11756 16544 11989 16572
rect 11756 16532 11762 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 10594 16504 10600 16516
rect 6012 16476 10600 16504
rect 10594 16464 10600 16476
rect 10652 16464 10658 16516
rect 12253 16507 12311 16513
rect 12253 16473 12265 16507
rect 12299 16504 12311 16507
rect 12526 16504 12532 16516
rect 12299 16476 12532 16504
rect 12299 16473 12311 16476
rect 12253 16467 12311 16473
rect 12526 16464 12532 16476
rect 12584 16464 12590 16516
rect 12710 16464 12716 16516
rect 12768 16464 12774 16516
rect 14274 16464 14280 16516
rect 14332 16504 14338 16516
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 14332 16476 14565 16504
rect 14332 16464 14338 16476
rect 14553 16473 14565 16476
rect 14599 16473 14611 16507
rect 14553 16467 14611 16473
rect 15010 16464 15016 16516
rect 15068 16464 15074 16516
rect 17052 16504 17080 16612
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 19334 16640 19340 16652
rect 17451 16612 19340 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 22278 16640 22284 16652
rect 19475 16612 22284 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 22646 16640 22652 16652
rect 22603 16612 22652 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 17126 16532 17132 16584
rect 17184 16532 17190 16584
rect 21818 16532 21824 16584
rect 21876 16532 21882 16584
rect 23658 16532 23664 16584
rect 23716 16532 23722 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16572 24639 16575
rect 24854 16572 24860 16584
rect 24627 16544 24860 16572
rect 24627 16541 24639 16544
rect 24581 16535 24639 16541
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 25225 16575 25283 16581
rect 25225 16541 25237 16575
rect 25271 16572 25283 16575
rect 25498 16572 25504 16584
rect 25271 16544 25504 16572
rect 25271 16541 25283 16544
rect 25225 16535 25283 16541
rect 25498 16532 25504 16544
rect 25556 16532 25562 16584
rect 17310 16504 17316 16516
rect 17052 16476 17316 16504
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 17736 16476 17894 16504
rect 17736 16464 17742 16476
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19392 16476 20194 16504
rect 19392 16464 19398 16476
rect 2593 16439 2651 16445
rect 2593 16405 2605 16439
rect 2639 16405 2651 16439
rect 2593 16399 2651 16405
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 5166 16436 5172 16448
rect 3283 16408 5172 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 5626 16396 5632 16448
rect 5684 16436 5690 16448
rect 11974 16436 11980 16448
rect 5684 16408 11980 16436
rect 5684 16396 5690 16408
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12342 16396 12348 16448
rect 12400 16436 12406 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12400 16408 13737 16436
rect 12400 16396 12406 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 16485 16439 16543 16445
rect 16485 16436 16497 16439
rect 13872 16408 16497 16436
rect 13872 16396 13878 16408
rect 16485 16405 16497 16408
rect 16531 16405 16543 16439
rect 16485 16399 16543 16405
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 18877 16439 18935 16445
rect 18877 16436 18889 16439
rect 17276 16408 18889 16436
rect 17276 16396 17282 16408
rect 18877 16405 18889 16408
rect 18923 16405 18935 16439
rect 18877 16399 18935 16405
rect 19150 16396 19156 16448
rect 19208 16436 19214 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 19208 16408 21189 16436
rect 19208 16396 19214 16408
rect 21177 16405 21189 16408
rect 21223 16436 21235 16439
rect 21358 16436 21364 16448
rect 21223 16408 21364 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21358 16396 21364 16408
rect 21416 16396 21422 16448
rect 21637 16439 21695 16445
rect 21637 16405 21649 16439
rect 21683 16436 21695 16439
rect 21726 16436 21732 16448
rect 21683 16408 21732 16436
rect 21683 16405 21695 16408
rect 21637 16399 21695 16405
rect 21726 16396 21732 16408
rect 21784 16396 21790 16448
rect 23934 16396 23940 16448
rect 23992 16436 23998 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23992 16408 24041 16436
rect 23992 16396 23998 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3510 16232 3516 16244
rect 3283 16204 3516 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 3878 16192 3884 16244
rect 3936 16192 3942 16244
rect 4525 16235 4583 16241
rect 4525 16201 4537 16235
rect 4571 16232 4583 16235
rect 5626 16232 5632 16244
rect 4571 16204 5632 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 5626 16192 5632 16204
rect 5684 16192 5690 16244
rect 6270 16192 6276 16244
rect 6328 16232 6334 16244
rect 6328 16204 6684 16232
rect 6328 16192 6334 16204
rect 6454 16164 6460 16176
rect 4080 16136 6460 16164
rect 2130 16056 2136 16108
rect 2188 16056 2194 16108
rect 2777 16099 2835 16105
rect 2777 16065 2789 16099
rect 2823 16096 2835 16099
rect 3418 16096 3424 16108
rect 2823 16068 3424 16096
rect 2823 16065 2835 16068
rect 2777 16059 2835 16065
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 4080 16105 4108 16136
rect 6454 16124 6460 16136
rect 6512 16124 6518 16176
rect 6656 16164 6684 16204
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 6788 16204 9444 16232
rect 6788 16192 6794 16204
rect 6656 16136 8432 16164
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 5316 16068 5457 16096
rect 5316 16056 5322 16068
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 8018 16056 8024 16108
rect 8076 16056 8082 16108
rect 2222 15988 2228 16040
rect 2280 16028 2286 16040
rect 5169 16031 5227 16037
rect 2280 16000 3188 16028
rect 2280 15988 2286 16000
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 2866 15960 2872 15972
rect 1995 15932 2872 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 2866 15920 2872 15932
rect 2924 15920 2930 15972
rect 3160 15960 3188 16000
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5350 16028 5356 16040
rect 5215 16000 5356 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 6549 16031 6607 16037
rect 6549 15997 6561 16031
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 6564 15960 6592 15991
rect 6822 15988 6828 16040
rect 6880 15988 6886 16040
rect 7006 15988 7012 16040
rect 7064 16028 7070 16040
rect 8404 16028 8432 16136
rect 8478 16124 8484 16176
rect 8536 16164 8542 16176
rect 9416 16164 9444 16204
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 10376 16204 10793 16232
rect 10376 16192 10382 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 10781 16195 10839 16201
rect 10873 16235 10931 16241
rect 10873 16201 10885 16235
rect 10919 16232 10931 16235
rect 14369 16235 14427 16241
rect 10919 16204 13492 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 11882 16164 11888 16176
rect 8536 16136 9352 16164
rect 9416 16136 11888 16164
rect 8536 16124 8542 16136
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16096 8723 16099
rect 9030 16096 9036 16108
rect 8711 16068 9036 16096
rect 8711 16065 8723 16068
rect 8665 16059 8723 16065
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9324 16105 9352 16136
rect 11882 16124 11888 16136
rect 11940 16124 11946 16176
rect 12710 16124 12716 16176
rect 12768 16124 12774 16176
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 9950 16056 9956 16108
rect 10008 16056 10014 16108
rect 11514 16096 11520 16108
rect 10980 16068 11520 16096
rect 10980 16028 11008 16068
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 7064 16000 7972 16028
rect 8404 16000 11008 16028
rect 11057 16031 11115 16037
rect 7064 15988 7070 16000
rect 3160 15932 6592 15960
rect 7834 15920 7840 15972
rect 7892 15920 7898 15972
rect 7944 15960 7972 16000
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 9769 15963 9827 15969
rect 7944 15932 9260 15960
rect 2593 15895 2651 15901
rect 2593 15861 2605 15895
rect 2639 15892 2651 15895
rect 5534 15892 5540 15904
rect 2639 15864 5540 15892
rect 2639 15861 2651 15864
rect 2593 15855 2651 15861
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 8294 15892 8300 15904
rect 6144 15864 8300 15892
rect 6144 15852 6150 15864
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 8481 15895 8539 15901
rect 8481 15861 8493 15895
rect 8527 15892 8539 15895
rect 8754 15892 8760 15904
rect 8527 15864 8760 15892
rect 8527 15861 8539 15864
rect 8481 15855 8539 15861
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8996 15864 9137 15892
rect 8996 15852 9002 15864
rect 9125 15861 9137 15864
rect 9171 15861 9183 15895
rect 9232 15892 9260 15932
rect 9769 15929 9781 15963
rect 9815 15960 9827 15963
rect 10778 15960 10784 15972
rect 9815 15932 10784 15960
rect 9815 15929 9827 15932
rect 9769 15923 9827 15929
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 9232 15864 10425 15892
rect 9125 15855 9183 15861
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 11072 15892 11100 15991
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12342 16028 12348 16040
rect 12023 16000 12348 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 13464 16028 13492 16204
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 19337 16235 19395 16241
rect 19337 16232 19349 16235
rect 14415 16204 19349 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 19337 16201 19349 16204
rect 19383 16201 19395 16235
rect 19337 16195 19395 16201
rect 20901 16235 20959 16241
rect 20901 16201 20913 16235
rect 20947 16232 20959 16235
rect 20990 16232 20996 16244
rect 20947 16204 20996 16232
rect 20947 16201 20959 16204
rect 20901 16195 20959 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 21910 16192 21916 16244
rect 21968 16232 21974 16244
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 21968 16204 22477 16232
rect 21968 16192 21974 16204
rect 22465 16201 22477 16204
rect 22511 16201 22523 16235
rect 22465 16195 22523 16201
rect 22646 16192 22652 16244
rect 22704 16232 22710 16244
rect 23385 16235 23443 16241
rect 23385 16232 23397 16235
rect 22704 16204 23397 16232
rect 22704 16192 22710 16204
rect 23385 16201 23397 16204
rect 23431 16201 23443 16235
rect 23385 16195 23443 16201
rect 23842 16192 23848 16244
rect 23900 16192 23906 16244
rect 13722 16124 13728 16176
rect 13780 16164 13786 16176
rect 13780 16136 16068 16164
rect 13780 16124 13786 16136
rect 13538 16056 13544 16108
rect 13596 16096 13602 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13596 16068 14289 16096
rect 13596 16056 13602 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15194 16096 15200 16108
rect 15059 16068 15200 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15838 16056 15844 16108
rect 15896 16056 15902 16108
rect 13464 16000 14044 16028
rect 13909 15963 13967 15969
rect 13909 15960 13921 15963
rect 13188 15932 13921 15960
rect 11974 15892 11980 15904
rect 11072 15864 11980 15892
rect 10413 15855 10471 15861
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 13188 15892 13216 15932
rect 13909 15929 13921 15932
rect 13955 15929 13967 15963
rect 14016 15960 14044 16000
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 15212 16028 15240 16056
rect 16040 16037 16068 16136
rect 18782 16124 18788 16176
rect 18840 16164 18846 16176
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 18840 16136 19717 16164
rect 18840 16124 18846 16136
rect 19705 16133 19717 16136
rect 19751 16133 19763 16167
rect 19705 16127 19763 16133
rect 19797 16167 19855 16173
rect 19797 16133 19809 16167
rect 19843 16164 19855 16167
rect 19978 16164 19984 16176
rect 19843 16136 19984 16164
rect 19843 16133 19855 16136
rect 19797 16127 19855 16133
rect 19978 16124 19984 16136
rect 20036 16164 20042 16176
rect 21545 16167 21603 16173
rect 21545 16164 21557 16167
rect 20036 16136 21557 16164
rect 20036 16124 20042 16136
rect 21545 16133 21557 16136
rect 21591 16133 21603 16167
rect 24946 16164 24952 16176
rect 21545 16127 21603 16133
rect 22066 16136 24952 16164
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 19610 16096 19616 16108
rect 17175 16068 19616 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 19610 16056 19616 16068
rect 19668 16056 19674 16108
rect 21818 16096 21824 16108
rect 19720 16068 21824 16096
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15212 16000 15945 16028
rect 15933 15997 15945 16000
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 18874 15988 18880 16040
rect 18932 15988 18938 16040
rect 15473 15963 15531 15969
rect 15473 15960 15485 15963
rect 14016 15932 15485 15960
rect 13909 15923 13967 15929
rect 15473 15929 15485 15932
rect 15519 15929 15531 15963
rect 15473 15923 15531 15929
rect 16482 15920 16488 15972
rect 16540 15960 16546 15972
rect 19720 15960 19748 16068
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 19978 15988 19984 16040
rect 20036 15988 20042 16040
rect 20990 15988 20996 16040
rect 21048 15988 21054 16040
rect 21177 16031 21235 16037
rect 21177 15997 21189 16031
rect 21223 16028 21235 16031
rect 21266 16028 21272 16040
rect 21223 16000 21272 16028
rect 21223 15997 21235 16000
rect 21177 15991 21235 15997
rect 21266 15988 21272 16000
rect 21324 15988 21330 16040
rect 16540 15932 19748 15960
rect 20533 15963 20591 15969
rect 16540 15920 16546 15932
rect 20533 15929 20545 15963
rect 20579 15960 20591 15963
rect 22066 15960 22094 16136
rect 24946 16124 24952 16136
rect 25004 16124 25010 16176
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16096 22431 16099
rect 22738 16096 22744 16108
rect 22419 16068 22744 16096
rect 22419 16065 22431 16068
rect 22373 16059 22431 16065
rect 22738 16056 22744 16068
rect 22796 16056 22802 16108
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16096 23167 16099
rect 23198 16096 23204 16108
rect 23155 16068 23204 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22244 16000 22569 16028
rect 22244 15988 22250 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 20579 15932 22094 15960
rect 20579 15929 20591 15932
rect 20533 15923 20591 15929
rect 12400 15864 13216 15892
rect 12400 15852 12406 15864
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 13412 15864 13461 15892
rect 13412 15852 13418 15864
rect 13449 15861 13461 15864
rect 13495 15892 13507 15895
rect 14090 15892 14096 15904
rect 13495 15864 14096 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14642 15892 14648 15904
rect 14240 15864 14648 15892
rect 14240 15852 14246 15864
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15286 15892 15292 15904
rect 15243 15864 15292 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 16390 15892 16396 15904
rect 16264 15864 16396 15892
rect 16264 15852 16270 15864
rect 16390 15852 16396 15864
rect 16448 15892 16454 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16448 15864 16681 15892
rect 16448 15852 16454 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 19208 15864 22017 15892
rect 19208 15852 19214 15864
rect 22005 15861 22017 15864
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 23124 15892 23152 16059
rect 23198 16056 23204 16068
rect 23256 16056 23262 16108
rect 23753 16099 23811 16105
rect 23753 16096 23765 16099
rect 23308 16068 23765 16096
rect 23308 15904 23336 16068
rect 23753 16065 23765 16068
rect 23799 16065 23811 16099
rect 23753 16059 23811 16065
rect 24578 16056 24584 16108
rect 24636 16056 24642 16108
rect 23934 15988 23940 16040
rect 23992 15988 23998 16040
rect 22612 15864 23152 15892
rect 22612 15852 22618 15864
rect 23290 15852 23296 15904
rect 23348 15852 23354 15904
rect 25222 15852 25228 15904
rect 25280 15852 25286 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 2130 15648 2136 15700
rect 2188 15688 2194 15700
rect 2225 15691 2283 15697
rect 2225 15688 2237 15691
rect 2188 15660 2237 15688
rect 2188 15648 2194 15660
rect 2225 15657 2237 15660
rect 2271 15657 2283 15691
rect 2225 15651 2283 15657
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 3973 15691 4031 15697
rect 3973 15688 3985 15691
rect 2648 15660 3985 15688
rect 2648 15648 2654 15660
rect 3973 15657 3985 15660
rect 4019 15657 4031 15691
rect 3973 15651 4031 15657
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 6549 15691 6607 15697
rect 6549 15688 6561 15691
rect 4120 15660 6561 15688
rect 4120 15648 4126 15660
rect 6549 15657 6561 15660
rect 6595 15657 6607 15691
rect 6549 15651 6607 15657
rect 7742 15648 7748 15700
rect 7800 15648 7806 15700
rect 8018 15648 8024 15700
rect 8076 15648 8082 15700
rect 8297 15691 8355 15697
rect 8297 15657 8309 15691
rect 8343 15688 8355 15691
rect 8570 15688 8576 15700
rect 8343 15660 8576 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 2866 15580 2872 15632
rect 2924 15620 2930 15632
rect 5258 15620 5264 15632
rect 2924 15592 5264 15620
rect 2924 15580 2930 15592
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 7374 15580 7380 15632
rect 7432 15620 7438 15632
rect 7837 15623 7895 15629
rect 7837 15620 7849 15623
rect 7432 15592 7849 15620
rect 7432 15580 7438 15592
rect 7837 15589 7849 15592
rect 7883 15589 7895 15623
rect 7837 15583 7895 15589
rect 8404 15561 8432 15660
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 9217 15691 9275 15697
rect 9217 15657 9229 15691
rect 9263 15688 9275 15691
rect 9306 15688 9312 15700
rect 9263 15660 9312 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 16850 15688 16856 15700
rect 13188 15660 16856 15688
rect 9858 15620 9864 15632
rect 8496 15592 9864 15620
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15552 5411 15555
rect 8389 15555 8447 15561
rect 5399 15524 7880 15552
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4246 15484 4252 15496
rect 4203 15456 4252 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15484 4951 15487
rect 6733 15487 6791 15493
rect 4939 15456 5948 15484
rect 4939 15453 4951 15456
rect 4893 15447 4951 15453
rect 5920 15360 5948 15456
rect 6733 15453 6745 15487
rect 6779 15484 6791 15487
rect 6914 15484 6920 15496
rect 6779 15456 6920 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 6914 15444 6920 15456
rect 6972 15444 6978 15496
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 7742 15484 7748 15496
rect 7423 15456 7748 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 7852 15484 7880 15524
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 8496 15484 8524 15592
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 11882 15580 11888 15632
rect 11940 15620 11946 15632
rect 12713 15623 12771 15629
rect 12713 15620 12725 15623
rect 11940 15592 12725 15620
rect 11940 15580 11946 15592
rect 12713 15589 12725 15592
rect 12759 15589 12771 15623
rect 12713 15583 12771 15589
rect 13188 15561 13216 15660
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 17310 15648 17316 15700
rect 17368 15688 17374 15700
rect 17368 15660 18276 15688
rect 17368 15648 17374 15660
rect 15562 15580 15568 15632
rect 15620 15620 15626 15632
rect 16025 15623 16083 15629
rect 16025 15620 16037 15623
rect 15620 15592 16037 15620
rect 15620 15580 15626 15592
rect 16025 15589 16037 15592
rect 16071 15589 16083 15623
rect 16025 15583 16083 15589
rect 16390 15580 16396 15632
rect 16448 15580 16454 15632
rect 16574 15580 16580 15632
rect 16632 15580 16638 15632
rect 18248 15620 18276 15660
rect 18690 15648 18696 15700
rect 18748 15688 18754 15700
rect 19886 15688 19892 15700
rect 18748 15660 19892 15688
rect 18748 15648 18754 15660
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 19996 15660 23336 15688
rect 19996 15620 20024 15660
rect 18248 15592 20024 15620
rect 20717 15623 20775 15629
rect 20717 15589 20729 15623
rect 20763 15620 20775 15623
rect 22830 15620 22836 15632
rect 20763 15592 22836 15620
rect 20763 15589 20775 15592
rect 20717 15583 20775 15589
rect 22830 15580 22836 15592
rect 22888 15580 22894 15632
rect 23308 15620 23336 15660
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23937 15691 23995 15697
rect 23937 15688 23949 15691
rect 23440 15660 23949 15688
rect 23440 15648 23446 15660
rect 23937 15657 23949 15660
rect 23983 15657 23995 15691
rect 23937 15651 23995 15657
rect 24121 15623 24179 15629
rect 24121 15620 24133 15623
rect 23308 15592 24133 15620
rect 24121 15589 24133 15592
rect 24167 15620 24179 15623
rect 24578 15620 24584 15632
rect 24167 15592 24584 15620
rect 24167 15589 24179 15592
rect 24121 15583 24179 15589
rect 24578 15580 24584 15592
rect 24636 15580 24642 15632
rect 13173 15555 13231 15561
rect 9646 15524 12848 15552
rect 7852 15456 8524 15484
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15484 9459 15487
rect 9646 15484 9674 15524
rect 9447 15456 9674 15484
rect 9447 15453 9459 15456
rect 9401 15447 9459 15453
rect 10042 15444 10048 15496
rect 10100 15444 10106 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 9582 15416 9588 15428
rect 7208 15388 9588 15416
rect 4706 15308 4712 15360
rect 4764 15308 4770 15360
rect 5902 15308 5908 15360
rect 5960 15308 5966 15360
rect 7208 15357 7236 15388
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 10520 15416 10548 15447
rect 10686 15416 10692 15428
rect 10520 15388 10692 15416
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 10778 15376 10784 15428
rect 10836 15376 10842 15428
rect 12342 15416 12348 15428
rect 12006 15388 12348 15416
rect 12342 15376 12348 15388
rect 12400 15416 12406 15428
rect 12710 15416 12716 15428
rect 12400 15388 12716 15416
rect 12400 15376 12406 15388
rect 12710 15376 12716 15388
rect 12768 15376 12774 15428
rect 12820 15416 12848 15524
rect 13173 15521 13185 15555
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 14182 15552 14188 15564
rect 13403 15524 14188 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 16850 15552 16856 15564
rect 14332 15524 16856 15552
rect 14332 15512 14338 15524
rect 16850 15512 16856 15524
rect 16908 15552 16914 15564
rect 16945 15555 17003 15561
rect 16945 15552 16957 15555
rect 16908 15524 16957 15552
rect 16908 15512 16914 15524
rect 16945 15521 16957 15524
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 17218 15512 17224 15564
rect 17276 15552 17282 15564
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 17276 15524 20085 15552
rect 17276 15512 17282 15524
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20073 15515 20131 15521
rect 21174 15512 21180 15564
rect 21232 15512 21238 15564
rect 21358 15512 21364 15564
rect 21416 15512 21422 15564
rect 23290 15552 23296 15564
rect 21468 15524 23296 15552
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13814 15484 13820 15496
rect 13127 15456 13820 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 13906 15444 13912 15496
rect 13964 15444 13970 15496
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20530 15484 20536 15496
rect 20027 15456 20536 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 13924 15416 13952 15444
rect 12820 15388 13952 15416
rect 14553 15419 14611 15425
rect 14553 15385 14565 15419
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 7193 15351 7251 15357
rect 7193 15317 7205 15351
rect 7239 15317 7251 15351
rect 7193 15311 7251 15317
rect 9861 15351 9919 15357
rect 9861 15317 9873 15351
rect 9907 15348 9919 15351
rect 10594 15348 10600 15360
rect 9907 15320 10600 15348
rect 9907 15317 9919 15320
rect 9861 15311 9919 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 11606 15308 11612 15360
rect 11664 15348 11670 15360
rect 12253 15351 12311 15357
rect 12253 15348 12265 15351
rect 11664 15320 12265 15348
rect 11664 15308 11670 15320
rect 12253 15317 12265 15320
rect 12299 15317 12311 15351
rect 12253 15311 12311 15317
rect 13909 15351 13967 15357
rect 13909 15317 13921 15351
rect 13955 15348 13967 15351
rect 14090 15348 14096 15360
rect 13955 15320 14096 15348
rect 13955 15317 13967 15320
rect 13909 15311 13967 15317
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 14568 15348 14596 15379
rect 15010 15376 15016 15428
rect 15068 15376 15074 15428
rect 16666 15416 16672 15428
rect 15856 15388 16672 15416
rect 15856 15348 15884 15388
rect 16666 15376 16672 15388
rect 16724 15376 16730 15428
rect 17310 15376 17316 15428
rect 17368 15416 17374 15428
rect 17678 15416 17684 15428
rect 17368 15388 17684 15416
rect 17368 15376 17374 15388
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 18598 15376 18604 15428
rect 18656 15416 18662 15428
rect 18969 15419 19027 15425
rect 18969 15416 18981 15419
rect 18656 15388 18981 15416
rect 18656 15376 18662 15388
rect 18969 15385 18981 15388
rect 19015 15385 19027 15419
rect 18969 15379 19027 15385
rect 21174 15376 21180 15428
rect 21232 15416 21238 15428
rect 21468 15416 21496 15524
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15484 21971 15487
rect 22554 15484 22560 15496
rect 21959 15456 22560 15484
rect 21959 15453 21971 15456
rect 21913 15447 21971 15453
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 23017 15487 23075 15493
rect 23017 15453 23029 15487
rect 23063 15484 23075 15487
rect 23382 15484 23388 15496
rect 23063 15456 23388 15484
rect 23063 15453 23075 15456
rect 23017 15447 23075 15453
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 25406 15484 25412 15496
rect 24719 15456 25412 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 21232 15388 21496 15416
rect 21232 15376 21238 15388
rect 14568 15320 15884 15348
rect 16022 15308 16028 15360
rect 16080 15348 16086 15360
rect 19426 15348 19432 15360
rect 16080 15320 19432 15348
rect 16080 15308 16086 15320
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 19518 15308 19524 15360
rect 19576 15308 19582 15360
rect 19886 15308 19892 15360
rect 19944 15308 19950 15360
rect 20898 15308 20904 15360
rect 20956 15348 20962 15360
rect 21085 15351 21143 15357
rect 21085 15348 21097 15351
rect 20956 15320 21097 15348
rect 20956 15308 20962 15320
rect 21085 15317 21097 15320
rect 21131 15317 21143 15351
rect 21085 15311 21143 15317
rect 22186 15308 22192 15360
rect 22244 15348 22250 15360
rect 22370 15348 22376 15360
rect 22244 15320 22376 15348
rect 22244 15308 22250 15320
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 22554 15308 22560 15360
rect 22612 15308 22618 15360
rect 23566 15308 23572 15360
rect 23624 15348 23630 15360
rect 23661 15351 23719 15357
rect 23661 15348 23673 15351
rect 23624 15320 23673 15348
rect 23624 15308 23630 15320
rect 23661 15317 23673 15320
rect 23707 15317 23719 15351
rect 23661 15311 23719 15317
rect 25317 15351 25375 15357
rect 25317 15317 25329 15351
rect 25363 15348 25375 15351
rect 25958 15348 25964 15360
rect 25363 15320 25964 15348
rect 25363 15317 25375 15320
rect 25317 15311 25375 15317
rect 25958 15308 25964 15320
rect 26016 15308 26022 15360
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 4246 15104 4252 15156
rect 4304 15104 4310 15156
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 7006 15144 7012 15156
rect 4396 15116 7012 15144
rect 4396 15104 4402 15116
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 10042 15144 10048 15156
rect 9447 15116 10048 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 10321 15147 10379 15153
rect 10321 15113 10333 15147
rect 10367 15144 10379 15147
rect 10410 15144 10416 15156
rect 10367 15116 10416 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 13722 15144 13728 15156
rect 12676 15116 13728 15144
rect 12676 15104 12682 15116
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 16022 15144 16028 15156
rect 13872 15116 16028 15144
rect 13872 15104 13878 15116
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 18690 15144 18696 15156
rect 17144 15116 18696 15144
rect 6914 15036 6920 15088
rect 6972 15036 6978 15088
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 9732 15048 10640 15076
rect 9732 15036 9738 15048
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 9585 14875 9643 14881
rect 9585 14841 9597 14875
rect 9631 14872 9643 14875
rect 9674 14872 9680 14884
rect 9631 14844 9680 14872
rect 9631 14841 9643 14844
rect 9585 14835 9643 14841
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 10612 14804 10640 15048
rect 11882 15036 11888 15088
rect 11940 15076 11946 15088
rect 11977 15079 12035 15085
rect 11977 15076 11989 15079
rect 11940 15048 11989 15076
rect 11940 15036 11946 15048
rect 11977 15045 11989 15048
rect 12023 15045 12035 15079
rect 11977 15039 12035 15045
rect 12710 15036 12716 15088
rect 12768 15036 12774 15088
rect 16758 15076 16764 15088
rect 13924 15048 16764 15076
rect 11146 14968 11152 15020
rect 11204 14968 11210 15020
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13924 15008 13952 15048
rect 16758 15036 16764 15048
rect 16816 15036 16822 15088
rect 17144 15085 17172 15116
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 21542 15144 21548 15156
rect 18932 15116 21548 15144
rect 18932 15104 18938 15116
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 23934 15144 23940 15156
rect 23124 15116 23940 15144
rect 17129 15079 17187 15085
rect 17129 15045 17141 15079
rect 17175 15045 17187 15079
rect 17129 15039 17187 15045
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 19334 15076 19340 15088
rect 17276 15048 17618 15076
rect 18892 15048 19340 15076
rect 17276 15036 17282 15048
rect 13412 14980 13952 15008
rect 13412 14968 13418 14980
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 16574 15008 16580 15020
rect 15703 14980 16580 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11698 14940 11704 14952
rect 10744 14912 11704 14940
rect 10744 14900 10750 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11974 14900 11980 14952
rect 12032 14940 12038 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 12032 14912 13461 14940
rect 12032 14900 12038 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14940 14703 14943
rect 14734 14940 14740 14952
rect 14691 14912 14740 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14940 15255 14943
rect 16758 14940 16764 14952
rect 15243 14912 16764 14940
rect 15243 14909 15255 14912
rect 15197 14903 15255 14909
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 17126 14940 17132 14952
rect 16899 14912 17132 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 14458 14832 14464 14884
rect 14516 14872 14522 14884
rect 16301 14875 16359 14881
rect 16301 14872 16313 14875
rect 14516 14844 16313 14872
rect 14516 14832 14522 14844
rect 16301 14841 16313 14844
rect 16347 14841 16359 14875
rect 16301 14835 16359 14841
rect 16482 14832 16488 14884
rect 16540 14872 16546 14884
rect 16868 14872 16896 14903
rect 17126 14900 17132 14912
rect 17184 14900 17190 14952
rect 17678 14900 17684 14952
rect 17736 14940 17742 14952
rect 18598 14940 18604 14952
rect 17736 14912 18604 14940
rect 17736 14900 17742 14912
rect 18598 14900 18604 14912
rect 18656 14940 18662 14952
rect 18892 14949 18920 15048
rect 19334 15036 19340 15048
rect 19392 15076 19398 15088
rect 22097 15079 22155 15085
rect 19392 15048 20102 15076
rect 19392 15036 19398 15048
rect 22097 15045 22109 15079
rect 22143 15076 22155 15079
rect 22370 15076 22376 15088
rect 22143 15048 22376 15076
rect 22143 15045 22155 15048
rect 22097 15039 22155 15045
rect 22370 15036 22376 15048
rect 22428 15036 22434 15088
rect 23124 15085 23152 15116
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24581 15147 24639 15153
rect 24581 15113 24593 15147
rect 24627 15144 24639 15147
rect 24762 15144 24768 15156
rect 24627 15116 24768 15144
rect 24627 15113 24639 15116
rect 24581 15107 24639 15113
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 23109 15079 23167 15085
rect 23109 15045 23121 15079
rect 23155 15045 23167 15079
rect 23109 15039 23167 15045
rect 23750 15036 23756 15088
rect 23808 15036 23814 15088
rect 25130 15036 25136 15088
rect 25188 15036 25194 15088
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18656 14912 18889 14940
rect 18656 14900 18662 14912
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 19334 14900 19340 14952
rect 19392 14900 19398 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 20622 14940 20628 14952
rect 19659 14912 20628 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 20806 14900 20812 14952
rect 20864 14940 20870 14952
rect 21085 14943 21143 14949
rect 21085 14940 21097 14943
rect 20864 14912 21097 14940
rect 20864 14900 20870 14912
rect 21085 14909 21097 14912
rect 21131 14909 21143 14943
rect 21085 14903 21143 14909
rect 22278 14900 22284 14952
rect 22336 14940 22342 14952
rect 22833 14943 22891 14949
rect 22833 14940 22845 14943
rect 22336 14912 22845 14940
rect 22336 14900 22342 14912
rect 22833 14909 22845 14912
rect 22879 14909 22891 14943
rect 22833 14903 22891 14909
rect 19352 14872 19380 14900
rect 16540 14844 16896 14872
rect 16540 14832 16546 14844
rect 13814 14804 13820 14816
rect 10612 14776 13820 14804
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 13909 14807 13967 14813
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 15102 14804 15108 14816
rect 13955 14776 15108 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 16868 14804 16896 14844
rect 18156 14844 19380 14872
rect 25317 14875 25375 14881
rect 18156 14804 18184 14844
rect 25317 14841 25329 14875
rect 25363 14872 25375 14875
rect 25590 14872 25596 14884
rect 25363 14844 25596 14872
rect 25363 14841 25375 14844
rect 25317 14835 25375 14841
rect 25590 14832 25596 14844
rect 25648 14832 25654 14884
rect 16868 14776 18184 14804
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 18601 14807 18659 14813
rect 18601 14804 18613 14807
rect 18380 14776 18613 14804
rect 18380 14764 18386 14776
rect 18601 14773 18613 14776
rect 18647 14773 18659 14807
rect 18601 14767 18659 14773
rect 18690 14764 18696 14816
rect 18748 14804 18754 14816
rect 20714 14804 20720 14816
rect 18748 14776 20720 14804
rect 18748 14764 18754 14776
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 21358 14764 21364 14816
rect 21416 14764 21422 14816
rect 22189 14807 22247 14813
rect 22189 14773 22201 14807
rect 22235 14804 22247 14807
rect 25498 14804 25504 14816
rect 22235 14776 25504 14804
rect 22235 14773 22247 14776
rect 22189 14767 22247 14773
rect 25498 14764 25504 14776
rect 25556 14764 25562 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10091 14572 12020 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 11992 14532 12020 14572
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 18690 14600 18696 14612
rect 12492 14572 18696 14600
rect 12492 14560 12498 14572
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 19426 14560 19432 14612
rect 19484 14560 19490 14612
rect 19610 14560 19616 14612
rect 19668 14600 19674 14612
rect 20254 14600 20260 14612
rect 19668 14572 20260 14600
rect 19668 14560 19674 14572
rect 20254 14560 20260 14572
rect 20312 14600 20318 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 20312 14572 20453 14600
rect 20312 14560 20318 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 22094 14600 22100 14612
rect 20441 14563 20499 14569
rect 20548 14572 22100 14600
rect 13814 14532 13820 14544
rect 11992 14504 13820 14532
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 18233 14535 18291 14541
rect 18233 14501 18245 14535
rect 18279 14532 18291 14535
rect 18506 14532 18512 14544
rect 18279 14504 18512 14532
rect 18279 14501 18291 14504
rect 18233 14495 18291 14501
rect 18506 14492 18512 14504
rect 18564 14492 18570 14544
rect 18598 14492 18604 14544
rect 18656 14532 18662 14544
rect 20548 14532 20576 14572
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 22278 14560 22284 14612
rect 22336 14560 22342 14612
rect 18656 14504 20576 14532
rect 18656 14492 18662 14504
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 22554 14532 22560 14544
rect 20772 14504 22560 14532
rect 20772 14492 20778 14504
rect 22554 14492 22560 14504
rect 22612 14492 22618 14544
rect 2682 14424 2688 14476
rect 2740 14464 2746 14476
rect 5534 14464 5540 14476
rect 2740 14436 5540 14464
rect 2740 14424 2746 14436
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11606 14464 11612 14476
rect 11011 14436 11612 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12618 14464 12624 14476
rect 12483 14436 12624 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14550 14424 14556 14476
rect 14608 14424 14614 14476
rect 15102 14424 15108 14476
rect 15160 14464 15166 14476
rect 16761 14467 16819 14473
rect 15160 14436 16436 14464
rect 15160 14424 15166 14436
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14396 10287 14399
rect 10410 14396 10416 14408
rect 10275 14368 10416 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 10410 14356 10416 14368
rect 10468 14356 10474 14408
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 12342 14396 12348 14408
rect 12098 14368 12348 14396
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 12710 14356 12716 14408
rect 12768 14396 12774 14408
rect 13446 14396 13452 14408
rect 12768 14368 13452 14396
rect 12768 14356 12774 14368
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 12250 14288 12256 14340
rect 12308 14328 12314 14340
rect 14458 14328 14464 14340
rect 12308 14300 14464 14328
rect 12308 14288 12314 14300
rect 14458 14288 14464 14300
rect 14516 14288 14522 14340
rect 15010 14288 15016 14340
rect 15068 14288 15074 14340
rect 16408 14328 16436 14436
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 18322 14464 18328 14476
rect 16807 14436 18328 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 18708 14436 19993 14464
rect 16482 14356 16488 14408
rect 16540 14356 16546 14408
rect 18340 14396 18368 14424
rect 18708 14396 18736 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 22002 14464 22008 14476
rect 19981 14427 20039 14433
rect 20732 14436 22008 14464
rect 20732 14408 20760 14436
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 22738 14424 22744 14476
rect 22796 14424 22802 14476
rect 23474 14424 23480 14476
rect 23532 14464 23538 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23532 14436 23765 14464
rect 23532 14424 23538 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 23753 14427 23811 14433
rect 23937 14467 23995 14473
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24302 14464 24308 14476
rect 23983 14436 24308 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24302 14424 24308 14436
rect 24360 14424 24366 14476
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 18340 14368 18736 14396
rect 19306 14368 19809 14396
rect 16408 14300 17172 14328
rect 12897 14263 12955 14269
rect 12897 14229 12909 14263
rect 12943 14260 12955 14263
rect 13722 14260 13728 14272
rect 12943 14232 13728 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14918 14260 14924 14272
rect 13872 14232 14924 14260
rect 13872 14220 13878 14232
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 16666 14260 16672 14272
rect 16071 14232 16672 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 17144 14260 17172 14300
rect 17218 14288 17224 14340
rect 17276 14288 17282 14340
rect 18046 14288 18052 14340
rect 18104 14328 18110 14340
rect 19306 14328 19334 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 20714 14356 20720 14408
rect 20772 14356 20778 14408
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21542 14396 21548 14408
rect 20864 14368 21548 14396
rect 20864 14356 20870 14368
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 18104 14300 19334 14328
rect 18104 14288 18110 14300
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 19484 14300 21588 14328
rect 19484 14288 19490 14300
rect 21560 14272 21588 14300
rect 22756 14272 22784 14424
rect 24486 14356 24492 14408
rect 24544 14396 24550 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24544 14368 24593 14396
rect 24544 14356 24550 14368
rect 24581 14365 24593 14368
rect 24627 14396 24639 14399
rect 24854 14396 24860 14408
rect 24627 14368 24860 14396
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 22925 14331 22983 14337
rect 22925 14297 22937 14331
rect 22971 14328 22983 14331
rect 23750 14328 23756 14340
rect 22971 14300 23756 14328
rect 22971 14297 22983 14300
rect 22925 14291 22983 14297
rect 23750 14288 23756 14300
rect 23808 14288 23814 14340
rect 17770 14260 17776 14272
rect 17144 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18656 14232 18705 14260
rect 18656 14220 18662 14232
rect 18693 14229 18705 14232
rect 18739 14229 18751 14263
rect 18693 14223 18751 14229
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19300 14232 19901 14260
rect 19300 14220 19306 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 19889 14223 19947 14229
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 21082 14260 21088 14272
rect 20220 14232 21088 14260
rect 20220 14220 20226 14232
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 21542 14220 21548 14272
rect 21600 14220 21606 14272
rect 22738 14220 22744 14272
rect 22796 14220 22802 14272
rect 23290 14220 23296 14272
rect 23348 14220 23354 14272
rect 23658 14220 23664 14272
rect 23716 14220 23722 14272
rect 23842 14220 23848 14272
rect 23900 14260 23906 14272
rect 25225 14263 25283 14269
rect 25225 14260 25237 14263
rect 23900 14232 25237 14260
rect 23900 14220 23906 14232
rect 25225 14229 25237 14232
rect 25271 14229 25283 14263
rect 25225 14223 25283 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10560 14028 10609 14056
rect 10560 14016 10566 14028
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 10597 14019 10655 14025
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14025 11023 14059
rect 10965 14019 11023 14025
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 10980 13988 11008 14019
rect 11606 14016 11612 14068
rect 11664 14016 11670 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12710 14056 12716 14068
rect 12299 14028 12716 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 12897 14059 12955 14065
rect 12897 14025 12909 14059
rect 12943 14056 12955 14059
rect 13354 14056 13360 14068
rect 12943 14028 13360 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 17037 14059 17095 14065
rect 13648 14028 16160 14056
rect 10284 13960 11008 13988
rect 10284 13948 10290 13960
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 11149 13923 11207 13929
rect 9456 13892 11100 13920
rect 9456 13880 9462 13892
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 11072 13852 11100 13892
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11624 13920 11652 14016
rect 13648 13988 13676 14028
rect 14274 13988 14280 14000
rect 11195 13892 11652 13920
rect 11716 13960 13676 13988
rect 13740 13960 14280 13988
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11716 13852 11744 13960
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13920 11851 13923
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11839 13892 11989 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 11977 13889 11989 13892
rect 12023 13920 12035 13923
rect 12342 13920 12348 13932
rect 12023 13892 12348 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 13740 13929 13768 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14458 13948 14464 14000
rect 14516 13948 14522 14000
rect 16132 13997 16160 14028
rect 17037 14025 17049 14059
rect 17083 14025 17095 14059
rect 17037 14019 17095 14025
rect 16117 13991 16175 13997
rect 16117 13957 16129 13991
rect 16163 13957 16175 13991
rect 17052 13988 17080 14019
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19392 14028 19533 14056
rect 19392 14016 19398 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20349 14059 20407 14065
rect 20349 14025 20361 14059
rect 20395 14056 20407 14059
rect 20806 14056 20812 14068
rect 20395 14028 20812 14056
rect 20395 14025 20407 14028
rect 20349 14019 20407 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21048 14028 21833 14056
rect 21048 14016 21054 14028
rect 21821 14025 21833 14028
rect 21867 14056 21879 14059
rect 22189 14059 22247 14065
rect 21867 14028 22140 14056
rect 21867 14025 21879 14028
rect 21821 14019 21879 14025
rect 17678 13988 17684 14000
rect 17052 13960 17684 13988
rect 16117 13951 16175 13957
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 17770 13948 17776 14000
rect 17828 13988 17834 14000
rect 18233 13991 18291 13997
rect 17828 13960 18184 13988
rect 17828 13948 17834 13960
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 11072 13824 11744 13852
rect 9582 13744 9588 13796
rect 9640 13784 9646 13796
rect 12360 13784 12388 13880
rect 13096 13852 13124 13883
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 15068 13892 16681 13920
rect 15068 13880 15074 13892
rect 16669 13889 16681 13892
rect 16715 13920 16727 13923
rect 17218 13920 17224 13932
rect 16715 13892 17224 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 17862 13920 17868 13932
rect 17451 13892 17868 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 18156 13920 18184 13960
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18874 13988 18880 14000
rect 18279 13960 18880 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18874 13948 18880 13960
rect 18932 13948 18938 14000
rect 20438 13948 20444 14000
rect 20496 13988 20502 14000
rect 22112 13997 22140 14028
rect 22189 14025 22201 14059
rect 22235 14056 22247 14059
rect 22462 14056 22468 14068
rect 22235 14028 22468 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 24762 14056 24768 14068
rect 23492 14028 24768 14056
rect 21177 13991 21235 13997
rect 21177 13988 21189 13991
rect 20496 13960 21189 13988
rect 20496 13948 20502 13960
rect 21177 13957 21189 13960
rect 21223 13957 21235 13991
rect 21177 13951 21235 13957
rect 22097 13991 22155 13997
rect 22097 13957 22109 13991
rect 22143 13957 22155 13991
rect 22097 13951 22155 13957
rect 23109 13991 23167 13997
rect 23109 13957 23121 13991
rect 23155 13988 23167 13991
rect 23492 13988 23520 14028
rect 24762 14016 24768 14028
rect 24820 14016 24826 14068
rect 23155 13960 23520 13988
rect 23155 13957 23167 13960
rect 23109 13951 23167 13957
rect 23750 13948 23756 14000
rect 23808 13948 23814 14000
rect 20714 13920 20720 13932
rect 18156 13892 20720 13920
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13920 21143 13923
rect 21818 13920 21824 13932
rect 21131 13892 21824 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22336 13892 22845 13920
rect 22336 13880 22342 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 25130 13880 25136 13932
rect 25188 13920 25194 13932
rect 25406 13920 25412 13932
rect 25188 13892 25412 13920
rect 25188 13880 25194 13892
rect 25406 13880 25412 13892
rect 25464 13880 25470 13932
rect 13096 13824 13860 13852
rect 12710 13784 12716 13796
rect 9640 13756 11100 13784
rect 12360 13756 12716 13784
rect 9640 13744 9646 13756
rect 11072 13716 11100 13756
rect 12710 13744 12716 13756
rect 12768 13784 12774 13796
rect 13449 13787 13507 13793
rect 13449 13784 13461 13787
rect 12768 13756 13461 13784
rect 12768 13744 12774 13756
rect 13449 13753 13461 13756
rect 13495 13784 13507 13787
rect 13722 13784 13728 13796
rect 13495 13756 13728 13784
rect 13495 13753 13507 13756
rect 13449 13747 13507 13753
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 13832 13728 13860 13824
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 14608 13824 15485 13852
rect 14608 13812 14614 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16390 13852 16396 13864
rect 16347 13824 16396 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 17696 13784 17724 13815
rect 19242 13812 19248 13864
rect 19300 13852 19306 13864
rect 21174 13852 21180 13864
rect 19300 13824 21180 13852
rect 19300 13812 19306 13824
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13821 21327 13855
rect 21269 13815 21327 13821
rect 17644 13756 17724 13784
rect 17644 13744 17650 13756
rect 20622 13744 20628 13796
rect 20680 13784 20686 13796
rect 21284 13784 21312 13815
rect 20680 13756 21312 13784
rect 20680 13744 20686 13756
rect 22204 13728 22232 13880
rect 24302 13812 24308 13864
rect 24360 13852 24366 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 24360 13824 24593 13852
rect 24360 13812 24366 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 25038 13812 25044 13864
rect 25096 13852 25102 13864
rect 25317 13855 25375 13861
rect 25317 13852 25329 13855
rect 25096 13824 25329 13852
rect 25096 13812 25102 13824
rect 25317 13821 25329 13824
rect 25363 13821 25375 13855
rect 25317 13815 25375 13821
rect 24210 13744 24216 13796
rect 24268 13784 24274 13796
rect 24670 13784 24676 13796
rect 24268 13756 24676 13784
rect 24268 13744 24274 13756
rect 24670 13744 24676 13756
rect 24728 13744 24734 13796
rect 13354 13716 13360 13728
rect 11072 13688 13360 13716
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 13814 13676 13820 13728
rect 13872 13676 13878 13728
rect 13988 13719 14046 13725
rect 13988 13685 14000 13719
rect 14034 13716 14046 13719
rect 16022 13716 16028 13728
rect 14034 13688 16028 13716
rect 14034 13685 14046 13688
rect 13988 13679 14046 13685
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 17402 13716 17408 13728
rect 16816 13688 17408 13716
rect 16816 13676 16822 13688
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 19610 13676 19616 13728
rect 19668 13716 19674 13728
rect 19978 13716 19984 13728
rect 19668 13688 19984 13716
rect 19668 13676 19674 13688
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 20714 13676 20720 13728
rect 20772 13676 20778 13728
rect 22186 13676 22192 13728
rect 22244 13676 22250 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 13906 13472 13912 13524
rect 13964 13472 13970 13524
rect 15930 13512 15936 13524
rect 14016 13484 15936 13512
rect 13354 13404 13360 13456
rect 13412 13444 13418 13456
rect 14016 13444 14044 13484
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 19610 13512 19616 13524
rect 16080 13484 19616 13512
rect 16080 13472 16086 13484
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 19968 13515 20026 13521
rect 19968 13481 19980 13515
rect 20014 13512 20026 13515
rect 20162 13512 20168 13524
rect 20014 13484 20168 13512
rect 20014 13481 20026 13484
rect 19968 13475 20026 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 20622 13472 20628 13524
rect 20680 13512 20686 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 20680 13484 21465 13512
rect 20680 13472 20686 13484
rect 21453 13481 21465 13484
rect 21499 13481 21511 13515
rect 23661 13515 23719 13521
rect 23661 13512 23673 13515
rect 21453 13475 21511 13481
rect 21560 13484 23673 13512
rect 13412 13416 14044 13444
rect 13412 13404 13418 13416
rect 17770 13404 17776 13456
rect 17828 13444 17834 13456
rect 17828 13416 19380 13444
rect 17828 13404 17834 13416
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 15010 13376 15016 13388
rect 14608 13348 15016 13376
rect 14608 13336 14614 13348
rect 15010 13336 15016 13348
rect 15068 13336 15074 13388
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 16298 13376 16304 13388
rect 15160 13348 16304 13376
rect 15160 13336 15166 13348
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 18506 13376 18512 13388
rect 16807 13348 18512 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 11238 13240 11244 13252
rect 9631 13212 11244 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 11238 13200 11244 13212
rect 11296 13200 11302 13252
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10686 13172 10692 13184
rect 10100 13144 10692 13172
rect 10100 13132 10106 13144
rect 10686 13132 10692 13144
rect 10744 13172 10750 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10744 13144 10885 13172
rect 10744 13132 10750 13144
rect 10873 13141 10885 13144
rect 10919 13172 10931 13175
rect 11808 13172 11836 13271
rect 18046 13268 18052 13320
rect 18104 13308 18110 13320
rect 18693 13311 18751 13317
rect 18693 13308 18705 13311
rect 18104 13280 18705 13308
rect 18104 13268 18110 13280
rect 18693 13277 18705 13280
rect 18739 13277 18751 13311
rect 18693 13271 18751 13277
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 12069 13243 12127 13249
rect 12069 13240 12081 13243
rect 12032 13212 12081 13240
rect 12032 13200 12038 13212
rect 12069 13209 12081 13212
rect 12115 13209 12127 13243
rect 12069 13203 12127 13209
rect 12710 13200 12716 13252
rect 12768 13200 12774 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14550 13240 14556 13252
rect 14240 13212 14556 13240
rect 14240 13200 14246 13212
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 15010 13200 15016 13252
rect 15068 13200 15074 13252
rect 16758 13240 16764 13252
rect 15856 13212 16764 13240
rect 10919 13144 11836 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13412 13144 13553 13172
rect 13412 13132 13418 13144
rect 13541 13141 13553 13144
rect 13587 13172 13599 13175
rect 15856 13172 15884 13212
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 17218 13200 17224 13252
rect 17276 13200 17282 13252
rect 19352 13249 19380 13416
rect 21082 13404 21088 13456
rect 21140 13444 21146 13456
rect 21560 13444 21588 13484
rect 23661 13481 23673 13484
rect 23707 13481 23719 13515
rect 23661 13475 23719 13481
rect 26050 13444 26056 13456
rect 21140 13416 21588 13444
rect 25056 13416 26056 13444
rect 21140 13404 21146 13416
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13376 19763 13379
rect 19978 13376 19984 13388
rect 19751 13348 19984 13376
rect 19751 13345 19763 13348
rect 19705 13339 19763 13345
rect 19978 13336 19984 13348
rect 20036 13376 20042 13388
rect 25056 13385 25084 13416
rect 26050 13404 26056 13416
rect 26108 13404 26114 13456
rect 25041 13379 25099 13385
rect 20036 13348 21956 13376
rect 20036 13336 20042 13348
rect 21928 13317 21956 13348
rect 25041 13345 25053 13379
rect 25087 13345 25099 13379
rect 25041 13339 25099 13345
rect 25130 13336 25136 13388
rect 25188 13336 25194 13388
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13277 21971 13311
rect 21913 13271 21971 13277
rect 19337 13243 19395 13249
rect 19337 13209 19349 13243
rect 19383 13240 19395 13243
rect 21928 13240 21956 13271
rect 22094 13240 22100 13252
rect 19383 13212 20470 13240
rect 21928 13212 22100 13240
rect 19383 13209 19395 13212
rect 19337 13203 19395 13209
rect 22094 13200 22100 13212
rect 22152 13200 22158 13252
rect 22186 13200 22192 13252
rect 22244 13200 22250 13252
rect 24949 13243 25007 13249
rect 23414 13212 23520 13240
rect 23492 13184 23520 13212
rect 24949 13209 24961 13243
rect 24995 13240 25007 13243
rect 26050 13240 26056 13252
rect 24995 13212 26056 13240
rect 24995 13209 25007 13212
rect 24949 13203 25007 13209
rect 26050 13200 26056 13212
rect 26108 13200 26114 13252
rect 13587 13144 15884 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 17586 13172 17592 13184
rect 16356 13144 17592 13172
rect 16356 13132 16362 13144
rect 17586 13132 17592 13144
rect 17644 13172 17650 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 17644 13144 18245 13172
rect 17644 13132 17650 13144
rect 18233 13141 18245 13144
rect 18279 13141 18291 13175
rect 18233 13135 18291 13141
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19058 13172 19064 13184
rect 18932 13144 19064 13172
rect 18932 13132 18938 13144
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 23474 13132 23480 13184
rect 23532 13172 23538 13184
rect 23750 13172 23756 13184
rect 23532 13144 23756 13172
rect 23532 13132 23538 13144
rect 23750 13132 23756 13144
rect 23808 13172 23814 13184
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 23808 13144 23949 13172
rect 23808 13132 23814 13144
rect 23937 13141 23949 13144
rect 23983 13172 23995 13175
rect 24121 13175 24179 13181
rect 24121 13172 24133 13175
rect 23983 13144 24133 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 24121 13141 24133 13144
rect 24167 13141 24179 13175
rect 24121 13135 24179 13141
rect 24394 13132 24400 13184
rect 24452 13172 24458 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24452 13144 24593 13172
rect 24452 13132 24458 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11296 12940 11345 12968
rect 11296 12928 11302 12940
rect 11333 12937 11345 12940
rect 11379 12968 11391 12971
rect 11790 12968 11796 12980
rect 11379 12940 11796 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12710 12928 12716 12980
rect 12768 12928 12774 12980
rect 14274 12928 14280 12980
rect 14332 12928 14338 12980
rect 17770 12968 17776 12980
rect 17512 12940 17776 12968
rect 11808 12900 11836 12928
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 11808 12872 13001 12900
rect 12989 12869 13001 12872
rect 13035 12900 13047 12903
rect 15013 12903 15071 12909
rect 15013 12900 15025 12903
rect 13035 12872 15025 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 15013 12869 15025 12872
rect 15059 12869 15071 12903
rect 15013 12863 15071 12869
rect 17218 12860 17224 12912
rect 17276 12900 17282 12912
rect 17512 12900 17540 12940
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 19521 12971 19579 12977
rect 19521 12968 19533 12971
rect 18932 12940 19533 12968
rect 18932 12928 18938 12940
rect 19521 12937 19533 12940
rect 19567 12937 19579 12971
rect 19521 12931 19579 12937
rect 19794 12928 19800 12980
rect 19852 12968 19858 12980
rect 20717 12971 20775 12977
rect 20717 12968 20729 12971
rect 19852 12940 20729 12968
rect 19852 12928 19858 12940
rect 20717 12937 20729 12940
rect 20763 12937 20775 12971
rect 20717 12931 20775 12937
rect 22094 12928 22100 12980
rect 22152 12928 22158 12980
rect 22186 12928 22192 12980
rect 22244 12968 22250 12980
rect 23753 12971 23811 12977
rect 23753 12968 23765 12971
rect 22244 12940 23765 12968
rect 22244 12928 22250 12940
rect 23753 12937 23765 12940
rect 23799 12968 23811 12971
rect 25130 12968 25136 12980
rect 23799 12940 25136 12968
rect 23799 12937 23811 12940
rect 23753 12931 23811 12937
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 25222 12928 25228 12980
rect 25280 12968 25286 12980
rect 25317 12971 25375 12977
rect 25317 12968 25329 12971
rect 25280 12940 25329 12968
rect 25280 12928 25286 12940
rect 25317 12937 25329 12940
rect 25363 12937 25375 12971
rect 25317 12931 25375 12937
rect 19150 12900 19156 12912
rect 17276 12872 17618 12900
rect 18524 12872 19156 12900
rect 17276 12860 17282 12872
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12832 12035 12835
rect 12342 12832 12348 12844
rect 12023 12804 12348 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 14366 12792 14372 12844
rect 14424 12832 14430 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 14424 12804 15485 12832
rect 14424 12792 14430 12804
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16758 12832 16764 12844
rect 16347 12804 16764 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17494 12764 17500 12776
rect 17175 12736 17500 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 17494 12724 17500 12736
rect 17552 12764 17558 12776
rect 18322 12764 18328 12776
rect 17552 12736 18328 12764
rect 17552 12724 17558 12736
rect 18322 12724 18328 12736
rect 18380 12724 18386 12776
rect 18524 12708 18552 12872
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 19429 12903 19487 12909
rect 19429 12869 19441 12903
rect 19475 12900 19487 12903
rect 19610 12900 19616 12912
rect 19475 12872 19616 12900
rect 19475 12869 19487 12872
rect 19429 12863 19487 12869
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 22112 12900 22140 12928
rect 19720 12872 20944 12900
rect 19720 12832 19748 12872
rect 18984 12804 19748 12832
rect 18984 12776 19012 12804
rect 20530 12792 20536 12844
rect 20588 12832 20594 12844
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20588 12804 20637 12832
rect 20588 12792 20594 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 18966 12724 18972 12776
rect 19024 12724 19030 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 20809 12767 20867 12773
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 20916 12764 20944 12872
rect 22020 12872 22140 12900
rect 22281 12903 22339 12909
rect 22020 12841 22048 12872
rect 22281 12869 22293 12903
rect 22327 12900 22339 12903
rect 22370 12900 22376 12912
rect 22327 12872 22376 12900
rect 22327 12869 22339 12872
rect 22281 12863 22339 12869
rect 22370 12860 22376 12872
rect 22428 12900 22434 12912
rect 22554 12900 22560 12912
rect 22428 12872 22560 12900
rect 22428 12860 22434 12872
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 23382 12792 23388 12844
rect 23440 12792 23446 12844
rect 24210 12792 24216 12844
rect 24268 12792 24274 12844
rect 20916 12736 22094 12764
rect 20809 12727 20867 12733
rect 7282 12656 7288 12708
rect 7340 12696 7346 12708
rect 16117 12699 16175 12705
rect 16117 12696 16129 12699
rect 7340 12668 16129 12696
rect 7340 12656 7346 12668
rect 16117 12665 16129 12668
rect 16163 12665 16175 12699
rect 16117 12659 16175 12665
rect 18506 12656 18512 12708
rect 18564 12656 18570 12708
rect 18598 12656 18604 12708
rect 18656 12696 18662 12708
rect 19628 12696 19656 12727
rect 18656 12668 19656 12696
rect 18656 12656 18662 12668
rect 20622 12656 20628 12708
rect 20680 12696 20686 12708
rect 20824 12696 20852 12727
rect 20680 12668 20852 12696
rect 20680 12656 20686 12668
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11793 12631 11851 12637
rect 11793 12628 11805 12631
rect 11388 12600 11805 12628
rect 11388 12588 11394 12600
rect 11793 12597 11805 12600
rect 11839 12597 11851 12631
rect 11793 12591 11851 12597
rect 19058 12588 19064 12640
rect 19116 12588 19122 12640
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19978 12628 19984 12640
rect 19484 12600 19984 12628
rect 19484 12588 19490 12600
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20257 12631 20315 12637
rect 20257 12597 20269 12631
rect 20303 12628 20315 12631
rect 20346 12628 20352 12640
rect 20303 12600 20352 12628
rect 20303 12597 20315 12600
rect 20257 12591 20315 12597
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 20864 12600 21281 12628
rect 20864 12588 20870 12600
rect 21269 12597 21281 12600
rect 21315 12628 21327 12631
rect 21358 12628 21364 12640
rect 21315 12600 21364 12628
rect 21315 12597 21327 12600
rect 21269 12591 21327 12597
rect 21358 12588 21364 12600
rect 21416 12628 21422 12640
rect 21453 12631 21511 12637
rect 21453 12628 21465 12631
rect 21416 12600 21465 12628
rect 21416 12588 21422 12600
rect 21453 12597 21465 12600
rect 21499 12597 21511 12631
rect 22066 12628 22094 12736
rect 24857 12699 24915 12705
rect 24857 12696 24869 12699
rect 23308 12668 24869 12696
rect 23308 12628 23336 12668
rect 24857 12665 24869 12668
rect 24903 12665 24915 12699
rect 24857 12659 24915 12665
rect 22066 12600 23336 12628
rect 21453 12591 21511 12597
rect 24946 12588 24952 12640
rect 25004 12628 25010 12640
rect 25133 12631 25191 12637
rect 25133 12628 25145 12631
rect 25004 12600 25145 12628
rect 25004 12588 25010 12600
rect 25133 12597 25145 12600
rect 25179 12597 25191 12631
rect 25133 12591 25191 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 14185 12427 14243 12433
rect 14185 12393 14197 12427
rect 14231 12424 14243 12427
rect 14458 12424 14464 12436
rect 14231 12396 14464 12424
rect 14231 12393 14243 12396
rect 14185 12387 14243 12393
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 14752 12396 17448 12424
rect 14752 12297 14780 12396
rect 17420 12356 17448 12396
rect 17494 12384 17500 12436
rect 17552 12384 17558 12436
rect 22094 12424 22100 12436
rect 17880 12396 22100 12424
rect 17880 12356 17908 12396
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 22370 12384 22376 12436
rect 22428 12424 22434 12436
rect 24029 12427 24087 12433
rect 24029 12424 24041 12427
rect 22428 12396 24041 12424
rect 22428 12384 22434 12396
rect 24029 12393 24041 12396
rect 24075 12393 24087 12427
rect 24029 12387 24087 12393
rect 17420 12328 17908 12356
rect 17957 12359 18015 12365
rect 17957 12325 17969 12359
rect 18003 12325 18015 12359
rect 17957 12319 18015 12325
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16758 12288 16764 12300
rect 15795 12260 16764 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 17218 12288 17224 12300
rect 17092 12260 17224 12288
rect 17092 12248 17098 12260
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 17972 12288 18000 12319
rect 20990 12288 20996 12300
rect 17972 12260 20996 12288
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 22186 12288 22192 12300
rect 21416 12260 22192 12288
rect 21416 12248 21422 12260
rect 22186 12248 22192 12260
rect 22244 12288 22250 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 22244 12260 22293 12288
rect 22244 12248 22250 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 24302 12288 24308 12300
rect 22603 12260 24308 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 24302 12248 24308 12260
rect 24360 12248 24366 12300
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 5500 12192 12909 12220
rect 5500 12180 5506 12192
rect 12897 12189 12909 12192
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 14366 12220 14372 12232
rect 13219 12192 14372 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 15654 12220 15660 12232
rect 14507 12192 15660 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 16025 12155 16083 12161
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 16298 12152 16304 12164
rect 16071 12124 16304 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 16298 12112 16304 12124
rect 16356 12112 16362 12164
rect 16482 12112 16488 12164
rect 16540 12112 16546 12164
rect 17034 12044 17040 12096
rect 17092 12084 17098 12096
rect 18156 12084 18184 12183
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19392 12192 19441 12220
rect 19392 12180 19398 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 20806 12180 20812 12232
rect 20864 12220 20870 12232
rect 20864 12192 21404 12220
rect 20864 12180 20870 12192
rect 18690 12112 18696 12164
rect 18748 12112 18754 12164
rect 18874 12112 18880 12164
rect 18932 12112 18938 12164
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 19978 12152 19984 12164
rect 19760 12124 19984 12152
rect 19760 12112 19766 12124
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 21376 12152 21404 12192
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21637 12223 21695 12229
rect 21637 12220 21649 12223
rect 21508 12192 21649 12220
rect 21508 12180 21514 12192
rect 21637 12189 21649 12192
rect 21683 12189 21695 12223
rect 21637 12183 21695 12189
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 21376 12124 23046 12152
rect 17092 12056 18184 12084
rect 17092 12044 17098 12056
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 20622 12084 20628 12096
rect 19852 12056 20628 12084
rect 19852 12044 19858 12056
rect 20622 12044 20628 12056
rect 20680 12084 20686 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 20680 12056 21189 12084
rect 20680 12044 20686 12056
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 22940 12084 22968 12124
rect 23382 12084 23388 12096
rect 22940 12056 23388 12084
rect 21177 12047 21235 12053
rect 23382 12044 23388 12056
rect 23440 12084 23446 12096
rect 24946 12084 24952 12096
rect 23440 12056 24952 12084
rect 23440 12044 23446 12056
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 25222 12044 25228 12096
rect 25280 12044 25286 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 14090 11880 14096 11892
rect 12820 11852 14096 11880
rect 5810 11772 5816 11824
rect 5868 11812 5874 11824
rect 12710 11812 12716 11824
rect 5868 11784 12716 11812
rect 5868 11772 5874 11784
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 12820 11753 12848 11852
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14550 11840 14556 11892
rect 14608 11840 14614 11892
rect 15102 11840 15108 11892
rect 15160 11840 15166 11892
rect 15565 11883 15623 11889
rect 15565 11880 15577 11883
rect 15212 11852 15577 11880
rect 13081 11815 13139 11821
rect 13081 11781 13093 11815
rect 13127 11812 13139 11815
rect 13354 11812 13360 11824
rect 13127 11784 13360 11812
rect 13127 11781 13139 11784
rect 13081 11775 13139 11781
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 14458 11812 14464 11824
rect 14306 11798 14464 11812
rect 14292 11784 14464 11798
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14292 11676 14320 11784
rect 14458 11772 14464 11784
rect 14516 11812 14522 11824
rect 15212 11812 15240 11852
rect 15565 11849 15577 11852
rect 15611 11880 15623 11883
rect 16482 11880 16488 11892
rect 15611 11852 16488 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 16482 11840 16488 11852
rect 16540 11880 16546 11892
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 16540 11852 16681 11880
rect 16540 11840 16546 11852
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 19334 11880 19340 11892
rect 16669 11843 16727 11849
rect 17144 11852 19340 11880
rect 15838 11812 15844 11824
rect 14516 11784 15240 11812
rect 15304 11784 15844 11812
rect 14516 11772 14522 11784
rect 15304 11753 15332 11784
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 17144 11753 17172 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 22186 11880 22192 11892
rect 21600 11852 22192 11880
rect 21600 11840 21606 11852
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 22278 11840 22284 11892
rect 22336 11840 22342 11892
rect 17310 11772 17316 11824
rect 17368 11812 17374 11824
rect 19705 11815 19763 11821
rect 17368 11784 17894 11812
rect 17368 11772 17374 11784
rect 19705 11781 19717 11815
rect 19751 11812 19763 11815
rect 19794 11812 19800 11824
rect 19751 11784 19800 11812
rect 19751 11781 19763 11784
rect 19705 11775 19763 11781
rect 19794 11772 19800 11784
rect 19852 11772 19858 11824
rect 20990 11772 20996 11824
rect 21048 11812 21054 11824
rect 22296 11812 22324 11840
rect 21048 11784 22324 11812
rect 23293 11815 23351 11821
rect 21048 11772 21054 11784
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 13872 11648 14320 11676
rect 16316 11676 16344 11707
rect 19426 11704 19432 11756
rect 19484 11704 19490 11756
rect 20806 11704 20812 11756
rect 20864 11744 20870 11756
rect 21542 11744 21548 11756
rect 20864 11716 21548 11744
rect 20864 11704 20870 11716
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 22278 11704 22284 11756
rect 22336 11704 22342 11756
rect 23934 11704 23940 11756
rect 23992 11704 23998 11756
rect 17405 11679 17463 11685
rect 16316 11648 17264 11676
rect 13872 11636 13878 11648
rect 16117 11611 16175 11617
rect 16117 11608 16129 11611
rect 14476 11580 16129 11608
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 14476 11540 14504 11580
rect 16117 11577 16129 11580
rect 16163 11577 16175 11611
rect 16117 11571 16175 11577
rect 12860 11512 14504 11540
rect 17236 11540 17264 11648
rect 17405 11645 17417 11679
rect 17451 11676 17463 11679
rect 18598 11676 18604 11688
rect 17451 11648 18604 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 18708 11648 22094 11676
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 18708 11608 18736 11648
rect 19150 11608 19156 11620
rect 18564 11580 18736 11608
rect 18800 11580 19156 11608
rect 18564 11568 18570 11580
rect 18800 11540 18828 11580
rect 19150 11568 19156 11580
rect 19208 11568 19214 11620
rect 22066 11608 22094 11648
rect 22738 11608 22744 11620
rect 22066 11580 22744 11608
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 17236 11512 18828 11540
rect 18877 11543 18935 11549
rect 12860 11500 12866 11512
rect 18877 11509 18889 11543
rect 18923 11540 18935 11543
rect 19702 11540 19708 11552
rect 18923 11512 19708 11540
rect 18923 11509 18935 11512
rect 18877 11503 18935 11509
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 19886 11500 19892 11552
rect 19944 11540 19950 11552
rect 20346 11540 20352 11552
rect 19944 11512 20352 11540
rect 19944 11500 19950 11512
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 21174 11500 21180 11552
rect 21232 11500 21238 11552
rect 21542 11500 21548 11552
rect 21600 11500 21606 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 14884 11308 15485 11336
rect 14884 11296 14890 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16942 11336 16948 11348
rect 16807 11308 16948 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17402 11296 17408 11348
rect 17460 11296 17466 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 18782 11336 18788 11348
rect 18739 11308 18788 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 19426 11336 19432 11348
rect 18892 11308 19432 11336
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 18506 11268 18512 11280
rect 9180 11240 12434 11268
rect 9180 11228 9186 11240
rect 12406 11064 12434 11240
rect 14844 11240 18512 11268
rect 14844 11209 14872 11240
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17920 11172 18061 11200
rect 17920 11160 17926 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 15194 11132 15200 11144
rect 13587 11104 15200 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 15746 11132 15752 11144
rect 15703 11104 15752 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16666 11132 16672 11144
rect 16347 11104 16672 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11132 17003 11135
rect 17126 11132 17132 11144
rect 16991 11104 17132 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 18892 11141 18920 11308
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19628 11308 19840 11336
rect 19150 11228 19156 11280
rect 19208 11268 19214 11280
rect 19628 11268 19656 11308
rect 19208 11240 19656 11268
rect 19812 11268 19840 11308
rect 22097 11271 22155 11277
rect 22097 11268 22109 11271
rect 19812 11240 22109 11268
rect 19208 11228 19214 11240
rect 22097 11237 22109 11240
rect 22143 11237 22155 11271
rect 22097 11231 22155 11237
rect 19334 11200 19340 11212
rect 18984 11172 19340 11200
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11101 17647 11135
rect 17589 11095 17647 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 17034 11064 17040 11076
rect 12406 11036 17040 11064
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 17604 11064 17632 11095
rect 17954 11064 17960 11076
rect 17604 11036 17960 11064
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 18138 11024 18144 11076
rect 18196 11064 18202 11076
rect 18984 11064 19012 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19794 11200 19800 11212
rect 19444 11172 19800 11200
rect 19444 11064 19472 11172
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 19886 11160 19892 11212
rect 19944 11160 19950 11212
rect 20806 11200 20812 11212
rect 20088 11172 20812 11200
rect 20088 11132 20116 11172
rect 20806 11160 20812 11172
rect 20864 11160 20870 11212
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 24854 11200 24860 11212
rect 23891 11172 24860 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 25130 11160 25136 11212
rect 25188 11200 25194 11212
rect 25406 11200 25412 11212
rect 25188 11172 25412 11200
rect 25188 11160 25194 11172
rect 25406 11160 25412 11172
rect 25464 11160 25470 11212
rect 18196 11036 19012 11064
rect 19260 11036 19472 11064
rect 19628 11104 20116 11132
rect 18196 11024 18202 11036
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 19260 10996 19288 11036
rect 14792 10968 19288 10996
rect 19337 10999 19395 11005
rect 14792 10956 14798 10968
rect 19337 10965 19349 10999
rect 19383 10996 19395 10999
rect 19628 10996 19656 11104
rect 20162 11092 20168 11144
rect 20220 11132 20226 11144
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 20220 11104 20361 11132
rect 20220 11092 20226 11104
rect 20349 11101 20361 11104
rect 20395 11132 20407 11135
rect 20622 11132 20628 11144
rect 20395 11104 20628 11132
rect 20395 11101 20407 11104
rect 20349 11095 20407 11101
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21453 11135 21511 11141
rect 21453 11132 21465 11135
rect 21048 11104 21465 11132
rect 21048 11092 21054 11104
rect 21453 11101 21465 11104
rect 21499 11132 21511 11135
rect 22002 11132 22008 11144
rect 21499 11104 22008 11132
rect 21499 11101 21511 11104
rect 21453 11095 21511 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 24670 11132 24676 11144
rect 24627 11104 24676 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 24670 11092 24676 11104
rect 24728 11132 24734 11144
rect 25314 11132 25320 11144
rect 24728 11104 25320 11132
rect 24728 11092 24734 11104
rect 25314 11092 25320 11104
rect 25372 11092 25378 11144
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20070 11064 20076 11076
rect 19751 11036 20076 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 25225 11067 25283 11073
rect 25225 11033 25237 11067
rect 25271 11064 25283 11067
rect 25406 11064 25412 11076
rect 25271 11036 25412 11064
rect 25271 11033 25283 11036
rect 25225 11027 25283 11033
rect 25406 11024 25412 11036
rect 25464 11024 25470 11076
rect 19383 10968 19656 10996
rect 19383 10965 19395 10968
rect 19337 10959 19395 10965
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 20993 10999 21051 11005
rect 20993 10996 21005 10999
rect 19852 10968 21005 10996
rect 19852 10956 19858 10968
rect 20993 10965 21005 10968
rect 21039 10965 21051 10999
rect 20993 10959 21051 10965
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 8812 10764 12434 10792
rect 8812 10752 8818 10764
rect 12406 10724 12434 10764
rect 15746 10752 15752 10804
rect 15804 10752 15810 10804
rect 16666 10752 16672 10804
rect 16724 10752 16730 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17126 10792 17132 10804
rect 16991 10764 17132 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 17313 10795 17371 10801
rect 17313 10761 17325 10795
rect 17359 10792 17371 10795
rect 17405 10795 17463 10801
rect 17405 10792 17417 10795
rect 17359 10764 17417 10792
rect 17359 10761 17371 10764
rect 17313 10755 17371 10761
rect 17405 10761 17417 10764
rect 17451 10792 17463 10795
rect 17586 10792 17592 10804
rect 17451 10764 17592 10792
rect 17451 10761 17463 10764
rect 17405 10755 17463 10761
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 18693 10795 18751 10801
rect 18693 10792 18705 10795
rect 17920 10764 18705 10792
rect 17920 10752 17926 10764
rect 18693 10761 18705 10764
rect 18739 10761 18751 10795
rect 18693 10755 18751 10761
rect 19426 10752 19432 10804
rect 19484 10792 19490 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19484 10764 19809 10792
rect 19484 10752 19490 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 20070 10752 20076 10804
rect 20128 10752 20134 10804
rect 20162 10752 20168 10804
rect 20220 10752 20226 10804
rect 20346 10752 20352 10804
rect 20404 10792 20410 10804
rect 20533 10795 20591 10801
rect 20533 10792 20545 10795
rect 20404 10764 20545 10792
rect 20404 10752 20410 10764
rect 20533 10761 20545 10764
rect 20579 10761 20591 10795
rect 20533 10755 20591 10761
rect 18230 10724 18236 10736
rect 12406 10696 18236 10724
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 23293 10727 23351 10733
rect 18340 10696 22232 10724
rect 16298 10616 16304 10668
rect 16356 10616 16362 10668
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 18340 10656 18368 10696
rect 17972 10628 18368 10656
rect 18877 10659 18935 10665
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 17972 10588 18000 10628
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 19150 10656 19156 10668
rect 18923 10628 19156 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10656 19579 10659
rect 19567 10628 20852 10656
rect 19567 10625 19579 10628
rect 19521 10619 19579 10625
rect 14424 10560 18000 10588
rect 18049 10591 18107 10597
rect 14424 10548 14430 10560
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 19702 10588 19708 10600
rect 18095 10560 19708 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 20824 10588 20852 10628
rect 21266 10616 21272 10668
rect 21324 10616 21330 10668
rect 22094 10616 22100 10668
rect 22152 10616 22158 10668
rect 22204 10656 22232 10696
rect 23293 10693 23305 10727
rect 23339 10724 23351 10727
rect 24854 10724 24860 10736
rect 23339 10696 24860 10724
rect 23339 10693 23351 10696
rect 23293 10687 23351 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 22204 10628 23949 10656
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 24394 10588 24400 10600
rect 20824 10560 24400 10588
rect 24394 10548 24400 10560
rect 24452 10548 24458 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 13630 10480 13636 10532
rect 13688 10520 13694 10532
rect 16117 10523 16175 10529
rect 16117 10520 16129 10523
rect 13688 10492 16129 10520
rect 13688 10480 13694 10492
rect 16117 10489 16129 10492
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 19337 10523 19395 10529
rect 19337 10489 19349 10523
rect 19383 10520 19395 10523
rect 20806 10520 20812 10532
rect 19383 10492 20812 10520
rect 19383 10489 19395 10492
rect 19337 10483 19395 10489
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 21453 10523 21511 10529
rect 21453 10489 21465 10523
rect 21499 10520 21511 10523
rect 21910 10520 21916 10532
rect 21499 10492 21916 10520
rect 21499 10489 21511 10492
rect 21453 10483 21511 10489
rect 21910 10480 21916 10492
rect 21968 10480 21974 10532
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 15654 10208 15660 10260
rect 15712 10248 15718 10260
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 15712 10220 16773 10248
rect 15712 10208 15718 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 19978 10248 19984 10260
rect 16761 10211 16819 10217
rect 17788 10220 19984 10248
rect 15010 10140 15016 10192
rect 15068 10180 15074 10192
rect 16485 10183 16543 10189
rect 16485 10180 16497 10183
rect 15068 10152 16497 10180
rect 15068 10140 15074 10152
rect 16485 10149 16497 10152
rect 16531 10180 16543 10183
rect 17788 10180 17816 10220
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 22646 10248 22652 10260
rect 20088 10220 22652 10248
rect 16531 10152 17816 10180
rect 18049 10183 18107 10189
rect 16531 10149 16543 10152
rect 16485 10143 16543 10149
rect 18049 10149 18061 10183
rect 18095 10180 18107 10183
rect 20088 10180 20116 10220
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 18095 10152 20116 10180
rect 20180 10152 21496 10180
rect 18095 10149 18107 10152
rect 18049 10143 18107 10149
rect 18414 10112 18420 10124
rect 17604 10084 18420 10112
rect 17604 10053 17632 10084
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 19886 10112 19892 10124
rect 18892 10084 19892 10112
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 16960 9976 16988 10007
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 18892 10053 18920 10084
rect 19886 10072 19892 10084
rect 19944 10072 19950 10124
rect 18877 10047 18935 10053
rect 18524 10016 18828 10044
rect 18322 9976 18328 9988
rect 16960 9948 18328 9976
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 17405 9911 17463 9917
rect 17405 9877 17417 9911
rect 17451 9908 17463 9911
rect 18524 9908 18552 10016
rect 18598 9936 18604 9988
rect 18656 9976 18662 9988
rect 18656 9948 18736 9976
rect 18656 9936 18662 9948
rect 18708 9917 18736 9948
rect 17451 9880 18552 9908
rect 18693 9911 18751 9917
rect 17451 9877 17463 9880
rect 17405 9871 17463 9877
rect 18693 9877 18705 9911
rect 18739 9877 18751 9911
rect 18800 9908 18828 10016
rect 18877 10013 18889 10047
rect 18923 10013 18935 10047
rect 18877 10007 18935 10013
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10044 19671 10047
rect 20070 10044 20076 10056
rect 19659 10016 20076 10044
rect 19659 10013 19671 10016
rect 19613 10007 19671 10013
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20180 10044 20208 10152
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10112 20775 10115
rect 20898 10112 20904 10124
rect 20763 10084 20904 10112
rect 20763 10081 20775 10084
rect 20717 10075 20775 10081
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 21358 10072 21364 10124
rect 21416 10072 21422 10124
rect 21468 10112 21496 10152
rect 22738 10140 22744 10192
rect 22796 10180 22802 10192
rect 24581 10183 24639 10189
rect 24581 10180 24593 10183
rect 22796 10152 24593 10180
rect 22796 10140 22802 10152
rect 24581 10149 24593 10152
rect 24627 10149 24639 10183
rect 24581 10143 24639 10149
rect 23290 10112 23296 10124
rect 21468 10084 23296 10112
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 25133 10115 25191 10121
rect 25133 10112 25145 10115
rect 23440 10084 25145 10112
rect 23440 10072 23446 10084
rect 25133 10081 25145 10084
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 20180 10016 20269 10044
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 23474 10044 23480 10056
rect 22770 10016 23480 10044
rect 20257 10007 20315 10013
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 24946 10004 24952 10056
rect 25004 10044 25010 10056
rect 25041 10047 25099 10053
rect 25041 10044 25053 10047
rect 25004 10016 25053 10044
rect 25004 10004 25010 10016
rect 25041 10013 25053 10016
rect 25087 10013 25099 10047
rect 25041 10007 25099 10013
rect 19150 9936 19156 9988
rect 19208 9976 19214 9988
rect 20898 9976 20904 9988
rect 19208 9948 20904 9976
rect 19208 9936 19214 9948
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21174 9936 21180 9988
rect 21232 9976 21238 9988
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 21232 9948 21649 9976
rect 21232 9936 21238 9948
rect 21637 9945 21649 9948
rect 21683 9945 21695 9979
rect 23845 9979 23903 9985
rect 23845 9976 23857 9979
rect 21637 9939 21695 9945
rect 22940 9948 23857 9976
rect 19334 9908 19340 9920
rect 18800 9880 19340 9908
rect 18693 9871 18751 9877
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 19426 9868 19432 9920
rect 19484 9868 19490 9920
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 20073 9911 20131 9917
rect 20073 9908 20085 9911
rect 19944 9880 20085 9908
rect 19944 9868 19950 9880
rect 20073 9877 20085 9880
rect 20119 9877 20131 9911
rect 20073 9871 20131 9877
rect 20162 9868 20168 9920
rect 20220 9908 20226 9920
rect 22940 9908 22968 9948
rect 23845 9945 23857 9948
rect 23891 9945 23903 9979
rect 23845 9939 23903 9945
rect 24026 9936 24032 9988
rect 24084 9936 24090 9988
rect 20220 9880 22968 9908
rect 23109 9911 23167 9917
rect 20220 9868 20226 9880
rect 23109 9877 23121 9911
rect 23155 9908 23167 9911
rect 23382 9908 23388 9920
rect 23155 9880 23388 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 23382 9868 23388 9880
rect 23440 9868 23446 9920
rect 24946 9868 24952 9920
rect 25004 9868 25010 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 19426 9664 19432 9716
rect 19484 9704 19490 9716
rect 19484 9676 20668 9704
rect 19484 9664 19490 9676
rect 20162 9636 20168 9648
rect 19628 9608 20168 9636
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16632 9540 17049 9568
rect 16632 9528 16638 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17586 9528 17592 9580
rect 17644 9528 17650 9580
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 17828 9540 18245 9568
rect 17828 9528 17834 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 19150 9568 19156 9580
rect 18923 9540 19156 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 19628 9577 19656 9608
rect 20162 9596 20168 9608
rect 20220 9636 20226 9648
rect 20640 9636 20668 9676
rect 20220 9608 20576 9636
rect 20640 9608 22140 9636
rect 20220 9596 20226 9608
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 20257 9572 20315 9577
rect 20257 9571 20392 9572
rect 20257 9537 20269 9571
rect 20303 9544 20392 9571
rect 20303 9537 20315 9544
rect 20257 9531 20315 9537
rect 20364 9500 20392 9544
rect 17420 9472 20392 9500
rect 20548 9500 20576 9608
rect 20622 9528 20628 9580
rect 20680 9528 20686 9580
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9568 20867 9571
rect 20898 9568 20904 9580
rect 20855 9540 20904 9568
rect 20855 9537 20867 9540
rect 20809 9531 20867 9537
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9568 21051 9571
rect 21082 9568 21088 9580
rect 21039 9540 21088 9568
rect 21039 9537 21051 9540
rect 20993 9531 21051 9537
rect 21082 9528 21088 9540
rect 21140 9528 21146 9580
rect 21450 9528 21456 9580
rect 21508 9528 21514 9580
rect 22112 9577 22140 9608
rect 23290 9596 23296 9648
rect 23348 9596 23354 9648
rect 26142 9636 26148 9648
rect 23400 9608 26148 9636
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 23400 9500 23428 9608
rect 26142 9596 26148 9608
rect 26200 9596 26206 9648
rect 23937 9571 23995 9577
rect 23937 9537 23949 9571
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 20548 9472 23428 9500
rect 17420 9441 17448 9472
rect 17405 9435 17463 9441
rect 17405 9401 17417 9435
rect 17451 9401 17463 9435
rect 18693 9435 18751 9441
rect 18693 9432 18705 9435
rect 17405 9395 17463 9401
rect 17512 9404 18705 9432
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 17512 9364 17540 9404
rect 18693 9401 18705 9404
rect 18739 9401 18751 9435
rect 18693 9395 18751 9401
rect 19429 9435 19487 9441
rect 19429 9401 19441 9435
rect 19475 9432 19487 9435
rect 19610 9432 19616 9444
rect 19475 9404 19616 9432
rect 19475 9401 19487 9404
rect 19429 9395 19487 9401
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 20073 9435 20131 9441
rect 20073 9401 20085 9435
rect 20119 9432 20131 9435
rect 23952 9432 23980 9531
rect 24670 9460 24676 9512
rect 24728 9460 24734 9512
rect 20119 9404 23980 9432
rect 20119 9401 20131 9404
rect 20073 9395 20131 9401
rect 16080 9336 17540 9364
rect 18049 9367 18107 9373
rect 16080 9324 16086 9336
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 19702 9364 19708 9376
rect 18095 9336 19708 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 21266 9324 21272 9376
rect 21324 9324 21330 9376
rect 21450 9324 21456 9376
rect 21508 9364 21514 9376
rect 26418 9364 26424 9376
rect 21508 9336 26424 9364
rect 21508 9324 21514 9336
rect 26418 9324 26424 9336
rect 26476 9324 26482 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 14458 9160 14464 9172
rect 11839 9132 14464 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 17681 9163 17739 9169
rect 17681 9160 17693 9163
rect 17644 9132 17693 9160
rect 17644 9120 17650 9132
rect 17681 9129 17693 9132
rect 17727 9129 17739 9163
rect 17681 9123 17739 9129
rect 19426 9120 19432 9172
rect 19484 9120 19490 9172
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 20990 9160 20996 9172
rect 20947 9132 20996 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 21085 9163 21143 9169
rect 21085 9129 21097 9163
rect 21131 9160 21143 9163
rect 21542 9160 21548 9172
rect 21131 9132 21548 9160
rect 21131 9129 21143 9132
rect 21085 9123 21143 9129
rect 21542 9120 21548 9132
rect 21600 9160 21606 9172
rect 23474 9160 23480 9172
rect 21600 9132 23480 9160
rect 21600 9120 21606 9132
rect 23474 9120 23480 9132
rect 23532 9120 23538 9172
rect 24578 9120 24584 9172
rect 24636 9120 24642 9172
rect 25041 9163 25099 9169
rect 25041 9129 25053 9163
rect 25087 9160 25099 9163
rect 25130 9160 25136 9172
rect 25087 9132 25136 9160
rect 25087 9129 25099 9132
rect 25041 9123 25099 9129
rect 25130 9120 25136 9132
rect 25188 9120 25194 9172
rect 24946 9092 24952 9104
rect 20088 9064 24952 9092
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 18049 9027 18107 9033
rect 18049 8993 18061 9027
rect 18095 9024 18107 9027
rect 19702 9024 19708 9036
rect 18095 8996 19708 9024
rect 18095 8993 18107 8996
rect 18049 8987 18107 8993
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 20088 9033 20116 9064
rect 24946 9052 24952 9064
rect 25004 9052 25010 9104
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 8993 20131 9027
rect 21450 9024 21456 9036
rect 20073 8987 20131 8993
rect 20180 8996 21456 9024
rect 18322 8916 18328 8968
rect 18380 8916 18386 8968
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8956 19671 8959
rect 19978 8956 19984 8968
rect 19659 8928 19984 8956
rect 19659 8925 19671 8928
rect 19613 8919 19671 8925
rect 19978 8916 19984 8928
rect 20036 8956 20042 8968
rect 20180 8956 20208 8996
rect 21450 8984 21456 8996
rect 21508 8984 21514 9036
rect 21637 9027 21695 9033
rect 21637 8993 21649 9027
rect 21683 9024 21695 9027
rect 22002 9024 22008 9036
rect 21683 8996 22008 9024
rect 21683 8993 21695 8996
rect 21637 8987 21695 8993
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 9024 23903 9027
rect 24854 9024 24860 9036
rect 23891 8996 24860 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 20036 8928 20208 8956
rect 20717 8959 20775 8965
rect 20036 8916 20042 8928
rect 20717 8925 20729 8959
rect 20763 8956 20775 8959
rect 21082 8956 21088 8968
rect 20763 8928 21088 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 21082 8916 21088 8928
rect 21140 8916 21146 8968
rect 21358 8916 21364 8968
rect 21416 8916 21422 8968
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 21600 8928 22661 8956
rect 21600 8916 21606 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 9364 8860 10333 8888
rect 9364 8848 9370 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 12161 8891 12219 8897
rect 12161 8888 12173 8891
rect 11546 8860 12173 8888
rect 10321 8851 10379 8857
rect 12161 8857 12173 8860
rect 12207 8888 12219 8891
rect 13814 8888 13820 8900
rect 12207 8860 13820 8888
rect 12207 8857 12219 8860
rect 12161 8851 12219 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 21376 8888 21404 8916
rect 24118 8888 24124 8900
rect 21376 8860 24124 8888
rect 24118 8848 24124 8860
rect 24176 8848 24182 8900
rect 21542 8780 21548 8832
rect 21600 8820 21606 8832
rect 22186 8820 22192 8832
rect 21600 8792 22192 8820
rect 21600 8780 21606 8792
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 24489 8823 24547 8829
rect 24489 8820 24501 8823
rect 23532 8792 24501 8820
rect 23532 8780 23538 8792
rect 24489 8789 24501 8792
rect 24535 8820 24547 8823
rect 24857 8823 24915 8829
rect 24857 8820 24869 8823
rect 24535 8792 24869 8820
rect 24535 8789 24547 8792
rect 24489 8783 24547 8789
rect 24857 8789 24869 8792
rect 24903 8820 24915 8823
rect 25225 8823 25283 8829
rect 25225 8820 25237 8823
rect 24903 8792 25237 8820
rect 24903 8789 24915 8792
rect 24857 8783 24915 8789
rect 25225 8789 25237 8792
rect 25271 8820 25283 8823
rect 25409 8823 25467 8829
rect 25409 8820 25421 8823
rect 25271 8792 25421 8820
rect 25271 8789 25283 8792
rect 25225 8783 25283 8789
rect 25409 8789 25421 8792
rect 25455 8820 25467 8823
rect 26142 8820 26148 8832
rect 25455 8792 26148 8820
rect 25455 8789 25467 8792
rect 25409 8783 25467 8789
rect 26142 8780 26148 8792
rect 26200 8780 26206 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 19429 8619 19487 8625
rect 19429 8585 19441 8619
rect 19475 8616 19487 8619
rect 26510 8616 26516 8628
rect 19475 8588 22048 8616
rect 19475 8585 19487 8588
rect 19429 8579 19487 8585
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 14056 8520 19656 8548
rect 14056 8508 14062 8520
rect 18969 8483 19027 8489
rect 18969 8449 18981 8483
rect 19015 8480 19027 8483
rect 19518 8480 19524 8492
rect 19015 8452 19524 8480
rect 19015 8449 19027 8452
rect 18969 8443 19027 8449
rect 19518 8440 19524 8452
rect 19576 8440 19582 8492
rect 19628 8489 19656 8520
rect 19978 8508 19984 8560
rect 20036 8508 20042 8560
rect 20162 8508 20168 8560
rect 20220 8508 20226 8560
rect 20530 8508 20536 8560
rect 20588 8548 20594 8560
rect 21269 8551 21327 8557
rect 21269 8548 21281 8551
rect 20588 8520 21281 8548
rect 20588 8508 20594 8520
rect 21269 8517 21281 8520
rect 21315 8517 21327 8551
rect 21269 8511 21327 8517
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 20714 8440 20720 8492
rect 20772 8480 20778 8492
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20772 8452 20821 8480
rect 20772 8440 20778 8452
rect 20809 8449 20821 8452
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 20349 8415 20407 8421
rect 20349 8412 20361 8415
rect 19208 8384 20361 8412
rect 19208 8372 19214 8384
rect 20349 8381 20361 8384
rect 20395 8412 20407 8415
rect 21634 8412 21640 8424
rect 20395 8384 21640 8412
rect 20395 8381 20407 8384
rect 20349 8375 20407 8381
rect 21634 8372 21640 8384
rect 21692 8372 21698 8424
rect 22020 8412 22048 8588
rect 22112 8588 26516 8616
rect 22112 8489 22140 8588
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 23293 8551 23351 8557
rect 23293 8517 23305 8551
rect 23339 8548 23351 8551
rect 24854 8548 24860 8560
rect 23339 8520 24860 8548
rect 23339 8517 23351 8520
rect 23293 8511 23351 8517
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 22244 8452 23949 8480
rect 22244 8440 22250 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 22278 8412 22284 8424
rect 22020 8384 22284 8412
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 24762 8372 24768 8424
rect 24820 8372 24826 8424
rect 18785 8347 18843 8353
rect 18785 8313 18797 8347
rect 18831 8344 18843 8347
rect 18831 8316 20576 8344
rect 18831 8313 18843 8316
rect 18785 8307 18843 8313
rect 20548 8276 20576 8316
rect 20622 8304 20628 8356
rect 20680 8304 20686 8356
rect 20898 8304 20904 8356
rect 20956 8344 20962 8356
rect 25222 8344 25228 8356
rect 20956 8316 25228 8344
rect 20956 8304 20962 8316
rect 25222 8304 25228 8316
rect 25280 8304 25286 8356
rect 21634 8276 21640 8288
rect 20548 8248 21640 8276
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 15436 8044 18705 8072
rect 15436 8032 15442 8044
rect 18693 8041 18705 8044
rect 18739 8041 18751 8075
rect 18693 8035 18751 8041
rect 19981 8075 20039 8081
rect 19981 8041 19993 8075
rect 20027 8072 20039 8075
rect 22186 8072 22192 8084
rect 20027 8044 22192 8072
rect 20027 8041 20039 8044
rect 19981 8035 20039 8041
rect 22186 8032 22192 8044
rect 22244 8032 22250 8084
rect 24210 8032 24216 8084
rect 24268 8072 24274 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 24268 8044 24685 8072
rect 24268 8032 24274 8044
rect 24673 8041 24685 8044
rect 24719 8041 24731 8075
rect 24673 8035 24731 8041
rect 19705 8007 19763 8013
rect 19705 7973 19717 8007
rect 19751 8004 19763 8007
rect 21358 8004 21364 8016
rect 19751 7976 21364 8004
rect 19751 7973 19763 7976
rect 19705 7967 19763 7973
rect 21358 7964 21364 7976
rect 21416 7964 21422 8016
rect 22066 7976 22692 8004
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 22066 7936 22094 7976
rect 16448 7908 22094 7936
rect 16448 7896 16454 7908
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 18966 7868 18972 7880
rect 18923 7840 18972 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 19392 7840 20177 7868
rect 19392 7828 19398 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20898 7828 20904 7880
rect 20956 7828 20962 7880
rect 21542 7828 21548 7880
rect 21600 7828 21606 7880
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 22664 7877 22692 7976
rect 24486 7964 24492 8016
rect 24544 7964 24550 8016
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24854 7936 24860 7948
rect 23891 7908 24860 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24854 7896 24860 7908
rect 24912 7896 24918 7948
rect 22189 7871 22247 7877
rect 22189 7868 22201 7871
rect 21692 7840 22201 7868
rect 21692 7828 21698 7840
rect 22189 7837 22201 7840
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22649 7871 22707 7877
rect 22649 7837 22661 7871
rect 22695 7837 22707 7871
rect 22649 7831 22707 7837
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 25133 7871 25191 7877
rect 25133 7868 25145 7871
rect 24728 7840 25145 7868
rect 24728 7828 24734 7840
rect 25133 7837 25145 7840
rect 25179 7837 25191 7871
rect 25133 7831 25191 7837
rect 19058 7760 19064 7812
rect 19116 7800 19122 7812
rect 24946 7800 24952 7812
rect 19116 7772 20944 7800
rect 19116 7760 19122 7772
rect 20916 7744 20944 7772
rect 21376 7772 24952 7800
rect 20346 7692 20352 7744
rect 20404 7732 20410 7744
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 20404 7704 20729 7732
rect 20404 7692 20410 7704
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 20717 7695 20775 7701
rect 20898 7692 20904 7744
rect 20956 7692 20962 7744
rect 21376 7741 21404 7772
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 25317 7803 25375 7809
rect 25317 7769 25329 7803
rect 25363 7800 25375 7803
rect 25958 7800 25964 7812
rect 25363 7772 25964 7800
rect 25363 7769 25375 7772
rect 25317 7763 25375 7769
rect 25958 7760 25964 7772
rect 26016 7760 26022 7812
rect 21361 7735 21419 7741
rect 21361 7701 21373 7735
rect 21407 7701 21419 7735
rect 21361 7695 21419 7701
rect 22002 7692 22008 7744
rect 22060 7692 22066 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 6880 7488 6914 7528
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 19300 7500 19993 7528
rect 19300 7488 19306 7500
rect 19981 7497 19993 7500
rect 20027 7497 20039 7531
rect 25406 7528 25412 7540
rect 19981 7491 20039 7497
rect 20732 7500 25412 7528
rect 6886 7324 6914 7488
rect 20165 7395 20223 7401
rect 20165 7361 20177 7395
rect 20211 7392 20223 7395
rect 20732 7392 20760 7500
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 23293 7463 23351 7469
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24854 7460 24860 7472
rect 23339 7432 24860 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 20211 7364 20760 7392
rect 20809 7395 20867 7401
rect 20211 7361 20223 7364
rect 20165 7355 20223 7361
rect 20809 7361 20821 7395
rect 20855 7392 20867 7395
rect 20898 7392 20904 7404
rect 20855 7364 20904 7392
rect 20855 7361 20867 7364
rect 20809 7355 20867 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 21726 7392 21732 7404
rect 21499 7364 21732 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 21910 7352 21916 7404
rect 21968 7392 21974 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 21968 7364 22109 7392
rect 21968 7352 21974 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 6886 7296 21496 7324
rect 20625 7259 20683 7265
rect 20625 7225 20637 7259
rect 20671 7256 20683 7259
rect 21174 7256 21180 7268
rect 20671 7228 21180 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 21468 7256 21496 7296
rect 21542 7284 21548 7336
rect 21600 7324 21606 7336
rect 23952 7324 23980 7355
rect 25406 7352 25412 7404
rect 25464 7392 25470 7404
rect 26142 7392 26148 7404
rect 25464 7364 26148 7392
rect 25464 7352 25470 7364
rect 26142 7352 26148 7364
rect 26200 7352 26206 7404
rect 21600 7296 23980 7324
rect 21600 7284 21606 7296
rect 24670 7256 24676 7268
rect 21468 7228 24676 7256
rect 24670 7216 24676 7228
rect 24728 7256 24734 7268
rect 25130 7256 25136 7268
rect 24728 7228 25136 7256
rect 24728 7216 24734 7228
rect 25130 7216 25136 7228
rect 25188 7216 25194 7268
rect 20070 7148 20076 7200
rect 20128 7188 20134 7200
rect 21269 7191 21327 7197
rect 21269 7188 21281 7191
rect 20128 7160 21281 7188
rect 20128 7148 20134 7160
rect 21269 7157 21281 7160
rect 21315 7157 21327 7191
rect 21269 7151 21327 7157
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 20625 6987 20683 6993
rect 20625 6953 20637 6987
rect 20671 6984 20683 6987
rect 21542 6984 21548 6996
rect 20671 6956 21548 6984
rect 20671 6953 20683 6956
rect 20625 6947 20683 6953
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 24578 6876 24584 6928
rect 24636 6916 24642 6928
rect 25038 6916 25044 6928
rect 24636 6888 25044 6916
rect 24636 6876 24642 6888
rect 25038 6876 25044 6888
rect 25096 6876 25102 6928
rect 21266 6808 21272 6860
rect 21324 6808 21330 6860
rect 21545 6851 21603 6857
rect 21545 6817 21557 6851
rect 21591 6848 21603 6851
rect 23845 6851 23903 6857
rect 21591 6820 23796 6848
rect 21591 6817 21603 6820
rect 21545 6811 21603 6817
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 20180 6712 20208 6743
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 22646 6740 22652 6792
rect 22704 6740 22710 6792
rect 22830 6740 22836 6792
rect 22888 6740 22894 6792
rect 23768 6780 23796 6820
rect 23845 6817 23857 6851
rect 23891 6848 23903 6851
rect 24946 6848 24952 6860
rect 23891 6820 24952 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 25225 6851 25283 6857
rect 25225 6817 25237 6851
rect 25271 6848 25283 6851
rect 25406 6848 25412 6860
rect 25271 6820 25412 6848
rect 25271 6817 25283 6820
rect 25225 6811 25283 6817
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 23934 6780 23940 6792
rect 23768 6752 23940 6780
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 24854 6740 24860 6792
rect 24912 6740 24918 6792
rect 20346 6712 20352 6724
rect 20180 6684 20352 6712
rect 20346 6672 20352 6684
rect 20404 6712 20410 6724
rect 22848 6712 22876 6740
rect 20404 6684 22876 6712
rect 20404 6672 20410 6684
rect 23290 6672 23296 6724
rect 23348 6712 23354 6724
rect 24578 6712 24584 6724
rect 23348 6684 24584 6712
rect 23348 6672 23354 6684
rect 24578 6672 24584 6684
rect 24636 6672 24642 6724
rect 25409 6715 25467 6721
rect 25409 6681 25421 6715
rect 25455 6712 25467 6715
rect 25682 6712 25688 6724
rect 25455 6684 25688 6712
rect 25455 6681 25467 6684
rect 25409 6675 25467 6681
rect 25682 6672 25688 6684
rect 25740 6672 25746 6724
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 19981 6647 20039 6653
rect 19981 6644 19993 6647
rect 17276 6616 19993 6644
rect 17276 6604 17282 6616
rect 19981 6613 19993 6616
rect 20027 6613 20039 6647
rect 19981 6607 20039 6613
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 24673 6647 24731 6653
rect 24673 6644 24685 6647
rect 22888 6616 24685 6644
rect 22888 6604 22894 6616
rect 24673 6613 24685 6616
rect 24719 6613 24731 6647
rect 24673 6607 24731 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 20346 6400 20352 6452
rect 20404 6400 20410 6452
rect 21269 6443 21327 6449
rect 21269 6409 21281 6443
rect 21315 6440 21327 6443
rect 23658 6440 23664 6452
rect 21315 6412 23664 6440
rect 21315 6409 21327 6412
rect 21269 6403 21327 6409
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 24854 6372 24860 6384
rect 23339 6344 24860 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20496 6276 20821 6304
rect 20496 6264 20502 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 22002 6264 22008 6316
rect 22060 6304 22066 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 22060 6276 22109 6304
rect 22060 6264 22066 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6304 24179 6307
rect 25866 6304 25872 6316
rect 24167 6276 25872 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 25866 6264 25872 6276
rect 25924 6264 25930 6316
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 20625 6103 20683 6109
rect 20625 6069 20637 6103
rect 20671 6100 20683 6103
rect 23474 6100 23480 6112
rect 20671 6072 23480 6100
rect 20671 6069 20683 6072
rect 20625 6063 20683 6069
rect 23474 6060 23480 6072
rect 23532 6060 23538 6112
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 20625 5899 20683 5905
rect 20625 5865 20637 5899
rect 20671 5896 20683 5899
rect 22646 5896 22652 5908
rect 20671 5868 22652 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 22646 5856 22652 5868
rect 22704 5856 22710 5908
rect 25314 5856 25320 5908
rect 25372 5856 25378 5908
rect 19702 5788 19708 5840
rect 19760 5828 19766 5840
rect 21269 5831 21327 5837
rect 21269 5828 21281 5831
rect 19760 5800 21281 5828
rect 19760 5788 19766 5800
rect 21269 5797 21281 5800
rect 21315 5797 21327 5831
rect 21269 5791 21327 5797
rect 25225 5831 25283 5837
rect 25225 5797 25237 5831
rect 25271 5828 25283 5831
rect 25774 5828 25780 5840
rect 25271 5800 25780 5828
rect 25271 5797 25283 5800
rect 25225 5791 25283 5797
rect 25774 5788 25780 5800
rect 25832 5788 25838 5840
rect 21818 5720 21824 5772
rect 21876 5760 21882 5772
rect 22005 5763 22063 5769
rect 22005 5760 22017 5763
rect 21876 5732 22017 5760
rect 21876 5720 21882 5732
rect 22005 5729 22017 5732
rect 22051 5729 22063 5763
rect 22005 5723 22063 5729
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 20809 5695 20867 5701
rect 20809 5692 20821 5695
rect 20680 5664 20821 5692
rect 20680 5652 20686 5664
rect 20809 5661 20821 5664
rect 20855 5661 20867 5695
rect 20809 5655 20867 5661
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5692 21511 5695
rect 22554 5692 22560 5704
rect 21499 5664 22560 5692
rect 21499 5661 21511 5664
rect 21453 5655 21511 5661
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 22830 5652 22836 5704
rect 22888 5652 22894 5704
rect 23845 5695 23903 5701
rect 23845 5661 23857 5695
rect 23891 5692 23903 5695
rect 24946 5692 24952 5704
rect 23891 5664 24952 5692
rect 23891 5661 23903 5664
rect 23845 5655 23903 5661
rect 24946 5652 24952 5664
rect 25004 5652 25010 5704
rect 19610 5584 19616 5636
rect 19668 5624 19674 5636
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 19668 5596 24685 5624
rect 19668 5584 19674 5596
rect 24673 5593 24685 5596
rect 24719 5593 24731 5627
rect 24673 5587 24731 5593
rect 24857 5627 24915 5633
rect 24857 5593 24869 5627
rect 24903 5624 24915 5627
rect 25038 5624 25044 5636
rect 24903 5596 25044 5624
rect 24903 5593 24915 5596
rect 24857 5587 24915 5593
rect 25038 5584 25044 5596
rect 25096 5584 25102 5636
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 21269 5355 21327 5361
rect 21269 5321 21281 5355
rect 21315 5352 21327 5355
rect 21450 5352 21456 5364
rect 21315 5324 21456 5352
rect 21315 5321 21327 5324
rect 21269 5315 21327 5321
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 18322 5244 18328 5296
rect 18380 5284 18386 5296
rect 23293 5287 23351 5293
rect 18380 5256 22600 5284
rect 18380 5244 18386 5256
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 21453 5219 21511 5225
rect 21453 5216 21465 5219
rect 19944 5188 21465 5216
rect 19944 5176 19950 5188
rect 21453 5185 21465 5188
rect 21499 5185 21511 5219
rect 21453 5179 21511 5185
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22462 5216 22468 5228
rect 22327 5188 22468 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22572 5216 22600 5256
rect 23293 5253 23305 5287
rect 23339 5284 23351 5287
rect 24854 5284 24860 5296
rect 23339 5256 24860 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 22572 5188 23949 5216
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24670 5108 24676 5160
rect 24728 5108 24734 5160
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 8662 4808 8668 4820
rect 8619 4780 8668 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 25130 4768 25136 4820
rect 25188 4768 25194 4820
rect 21361 4743 21419 4749
rect 21361 4709 21373 4743
rect 21407 4740 21419 4743
rect 24578 4740 24584 4752
rect 21407 4712 24584 4740
rect 21407 4709 21419 4712
rect 21361 4703 21419 4709
rect 24578 4700 24584 4712
rect 24636 4700 24642 4752
rect 24670 4700 24676 4752
rect 24728 4700 24734 4752
rect 22738 4672 22744 4684
rect 22066 4644 22744 4672
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7064 4576 7941 4604
rect 7064 4564 7070 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 22066 4604 22094 4644
rect 22738 4632 22744 4644
rect 22796 4632 22802 4684
rect 25590 4672 25596 4684
rect 22848 4644 25596 4672
rect 22848 4613 22876 4644
rect 25590 4632 25596 4644
rect 25648 4632 25654 4684
rect 21591 4576 22094 4604
rect 22833 4607 22891 4613
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 22833 4573 22845 4607
rect 22879 4573 22891 4607
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 22833 4567 22891 4573
rect 22940 4576 24869 4604
rect 21174 4496 21180 4548
rect 21232 4536 21238 4548
rect 22940 4536 22968 4576
rect 24857 4573 24869 4576
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 21232 4508 22968 4536
rect 23845 4539 23903 4545
rect 21232 4496 21238 4508
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 24946 4536 24952 4548
rect 23891 4508 24952 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 22005 4471 22063 4477
rect 22005 4437 22017 4471
rect 22051 4468 22063 4471
rect 26050 4468 26056 4480
rect 22051 4440 26056 4468
rect 22051 4437 22063 4440
rect 22005 4431 22063 4437
rect 26050 4428 26056 4440
rect 26108 4428 26114 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 23952 4168 25176 4196
rect 23952 4137 23980 4168
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 22281 4131 22339 4137
rect 20303 4100 22232 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 22094 4060 22100 4072
rect 21315 4032 22100 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 22204 4060 22232 4100
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 23937 4131 23995 4137
rect 22327 4100 23428 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 23198 4060 23204 4072
rect 22204 4032 23204 4060
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23400 4060 23428 4100
rect 23937 4097 23949 4131
rect 23983 4097 23995 4131
rect 25038 4128 25044 4140
rect 23937 4091 23995 4097
rect 24044 4100 25044 4128
rect 24044 4060 24072 4100
rect 25038 4088 25044 4100
rect 25096 4088 25102 4140
rect 25148 4128 25176 4168
rect 25498 4128 25504 4140
rect 25148 4100 25504 4128
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 23400 4032 24072 4060
rect 23293 4023 23351 4029
rect 23308 3992 23336 4023
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 24946 3992 24952 4004
rect 23308 3964 24952 3992
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 23532 3556 24900 3584
rect 23532 3544 23538 3556
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7466 3516 7472 3528
rect 6871 3488 7472 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 19794 3476 19800 3528
rect 19852 3516 19858 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 19852 3488 20821 3516
rect 19852 3476 19858 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 24670 3516 24676 3528
rect 22879 3488 24676 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24872 3525 24900 3556
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 23845 3451 23903 3457
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24946 3448 24952 3460
rect 23891 3420 24952 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 24946 3408 24952 3420
rect 25004 3408 25010 3460
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 7248 3352 7481 3380
rect 7248 3340 7254 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 22278 3340 22284 3392
rect 22336 3380 22342 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 22336 3352 24685 3380
rect 22336 3340 22342 3352
rect 24673 3349 24685 3352
rect 24719 3349 24731 3383
rect 24673 3343 24731 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 7466 3136 7472 3188
rect 7524 3136 7530 3188
rect 25958 3176 25964 3188
rect 22066 3148 25964 3176
rect 22066 3108 22094 3148
rect 25958 3136 25964 3148
rect 26016 3136 26022 3188
rect 18432 3080 22094 3108
rect 23293 3111 23351 3117
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 18432 3049 18460 3080
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24854 3108 24860 3120
rect 23339 3080 24860 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 25130 3068 25136 3120
rect 25188 3068 25194 3120
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 18932 3012 20085 3040
rect 18932 3000 18938 3012
rect 20073 3009 20085 3012
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 22278 3000 22284 3052
rect 22336 3000 22342 3052
rect 24026 3000 24032 3052
rect 24084 3000 24090 3052
rect 19334 2932 19340 2984
rect 19392 2932 19398 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 25038 2972 25044 2984
rect 21315 2944 25044 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 6549 2839 6607 2845
rect 6549 2805 6561 2839
rect 6595 2836 6607 2839
rect 6730 2836 6736 2848
rect 6595 2808 6736 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 7006 2632 7012 2644
rect 6595 2604 7012 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 22830 2632 22836 2644
rect 19392 2604 22836 2632
rect 19392 2592 19398 2604
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 23382 2592 23388 2644
rect 23440 2592 23446 2644
rect 23400 2564 23428 2592
rect 21192 2536 23428 2564
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 6886 2468 7849 2496
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 6886 2428 6914 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 6779 2400 6914 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2428 20315 2431
rect 21192 2428 21220 2536
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2496 21327 2499
rect 23382 2496 23388 2508
rect 21315 2468 23388 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 20303 2400 21220 2428
rect 22833 2431 22891 2437
rect 20303 2397 20315 2400
rect 20257 2391 20315 2397
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 22848 2292 22876 2391
rect 24578 2388 24584 2440
rect 24636 2428 24642 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24636 2400 24777 2428
rect 24636 2388 24642 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 22848 2264 24593 2292
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 3056 26392 3108 26444
rect 3424 26392 3476 26444
rect 1952 26324 2004 26376
rect 18696 26324 18748 26376
rect 12808 24964 12860 25016
rect 14924 24964 14976 25016
rect 15476 24964 15528 25016
rect 20076 24964 20128 25016
rect 11612 24896 11664 24948
rect 13084 24896 13136 24948
rect 16212 24896 16264 24948
rect 18236 24896 18288 24948
rect 3700 24828 3752 24880
rect 18420 24828 18472 24880
rect 11888 24760 11940 24812
rect 12072 24760 12124 24812
rect 13544 24760 13596 24812
rect 18604 24760 18656 24812
rect 7472 24692 7524 24744
rect 20536 24692 20588 24744
rect 4160 24624 4212 24676
rect 13728 24624 13780 24676
rect 15016 24624 15068 24676
rect 21456 24624 21508 24676
rect 5816 24556 5868 24608
rect 12256 24556 12308 24608
rect 14096 24556 14148 24608
rect 17224 24556 17276 24608
rect 17592 24556 17644 24608
rect 24124 24556 24176 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 6736 24352 6788 24404
rect 4712 24284 4764 24336
rect 5356 24284 5408 24336
rect 11796 24352 11848 24404
rect 9772 24284 9824 24336
rect 6460 24216 6512 24268
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 5264 24148 5316 24200
rect 6736 24191 6788 24200
rect 6736 24157 6745 24191
rect 6745 24157 6779 24191
rect 6779 24157 6788 24191
rect 6736 24148 6788 24157
rect 9680 24216 9732 24268
rect 11244 24216 11296 24268
rect 7748 24148 7800 24200
rect 14096 24352 14148 24404
rect 16856 24352 16908 24404
rect 16948 24395 17000 24404
rect 16948 24361 16957 24395
rect 16957 24361 16991 24395
rect 16991 24361 17000 24395
rect 16948 24352 17000 24361
rect 13636 24284 13688 24336
rect 15476 24284 15528 24336
rect 15568 24327 15620 24336
rect 15568 24293 15577 24327
rect 15577 24293 15611 24327
rect 15611 24293 15620 24327
rect 15568 24284 15620 24293
rect 12348 24216 12400 24268
rect 14004 24216 14056 24268
rect 14556 24216 14608 24268
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 16212 24259 16264 24268
rect 16212 24225 16221 24259
rect 16221 24225 16255 24259
rect 16255 24225 16264 24259
rect 16212 24216 16264 24225
rect 19892 24352 19944 24404
rect 16488 24148 16540 24200
rect 17960 24216 18012 24268
rect 18236 24284 18288 24336
rect 23756 24352 23808 24404
rect 18328 24216 18380 24268
rect 5632 24080 5684 24132
rect 8392 24080 8444 24132
rect 8576 24080 8628 24132
rect 12164 24080 12216 24132
rect 12256 24080 12308 24132
rect 13820 24080 13872 24132
rect 4988 24012 5040 24064
rect 6552 24055 6604 24064
rect 6552 24021 6561 24055
rect 6561 24021 6595 24055
rect 6595 24021 6604 24055
rect 6552 24012 6604 24021
rect 10968 24012 11020 24064
rect 11796 24012 11848 24064
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 22652 24216 22704 24268
rect 25228 24259 25280 24268
rect 25228 24225 25237 24259
rect 25237 24225 25271 24259
rect 25271 24225 25280 24259
rect 25228 24216 25280 24225
rect 20168 24191 20220 24200
rect 20168 24157 20177 24191
rect 20177 24157 20211 24191
rect 20211 24157 20220 24191
rect 20168 24148 20220 24157
rect 20536 24191 20588 24200
rect 20536 24157 20545 24191
rect 20545 24157 20579 24191
rect 20579 24157 20588 24191
rect 20536 24148 20588 24157
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 22284 24191 22336 24200
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 25044 24148 25096 24200
rect 14740 24055 14792 24064
rect 14740 24021 14749 24055
rect 14749 24021 14783 24055
rect 14783 24021 14792 24055
rect 14740 24012 14792 24021
rect 14832 24055 14884 24064
rect 14832 24021 14841 24055
rect 14841 24021 14875 24055
rect 14875 24021 14884 24055
rect 14832 24012 14884 24021
rect 15568 24012 15620 24064
rect 17316 24055 17368 24064
rect 17316 24021 17325 24055
rect 17325 24021 17359 24055
rect 17359 24021 17368 24055
rect 17316 24012 17368 24021
rect 22468 24080 22520 24132
rect 18696 24012 18748 24064
rect 19524 24012 19576 24064
rect 21272 24055 21324 24064
rect 21272 24021 21281 24055
rect 21281 24021 21315 24055
rect 21315 24021 21324 24055
rect 21272 24012 21324 24021
rect 23020 24080 23072 24132
rect 23848 24012 23900 24064
rect 24124 24012 24176 24064
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 24676 24012 24728 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 3792 23808 3844 23860
rect 5172 23740 5224 23792
rect 7380 23740 7432 23792
rect 1860 23672 1912 23724
rect 4160 23672 4212 23724
rect 5632 23672 5684 23724
rect 7564 23672 7616 23724
rect 9312 23604 9364 23656
rect 5172 23536 5224 23588
rect 10692 23808 10744 23860
rect 10876 23783 10928 23792
rect 10876 23749 10885 23783
rect 10885 23749 10919 23783
rect 10919 23749 10928 23783
rect 10876 23740 10928 23749
rect 10140 23604 10192 23656
rect 11428 23604 11480 23656
rect 14740 23740 14792 23792
rect 15568 23740 15620 23792
rect 16120 23740 16172 23792
rect 24676 23808 24728 23860
rect 20260 23740 20312 23792
rect 11888 23672 11940 23724
rect 12164 23672 12216 23724
rect 11980 23604 12032 23656
rect 13820 23604 13872 23656
rect 13636 23536 13688 23588
rect 14740 23647 14792 23656
rect 14740 23613 14749 23647
rect 14749 23613 14783 23647
rect 14783 23613 14792 23647
rect 14740 23604 14792 23613
rect 17040 23672 17092 23724
rect 2228 23468 2280 23520
rect 6920 23468 6972 23520
rect 11796 23468 11848 23520
rect 11980 23468 12032 23520
rect 12440 23468 12492 23520
rect 14924 23468 14976 23520
rect 15384 23468 15436 23520
rect 16396 23468 16448 23520
rect 17592 23604 17644 23656
rect 17868 23468 17920 23520
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 18328 23647 18380 23656
rect 18328 23613 18337 23647
rect 18337 23613 18371 23647
rect 18371 23613 18380 23647
rect 18328 23604 18380 23613
rect 18696 23604 18748 23656
rect 21824 23604 21876 23656
rect 23020 23740 23072 23792
rect 24032 23740 24084 23792
rect 24400 23740 24452 23792
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 25780 23740 25832 23792
rect 23848 23672 23900 23724
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 25320 23672 25372 23724
rect 18512 23468 18564 23520
rect 18788 23468 18840 23520
rect 21916 23536 21968 23588
rect 19800 23511 19852 23520
rect 19800 23477 19809 23511
rect 19809 23477 19843 23511
rect 19843 23477 19852 23511
rect 19800 23468 19852 23477
rect 22192 23536 22244 23588
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 1768 23307 1820 23316
rect 1768 23273 1777 23307
rect 1777 23273 1811 23307
rect 1811 23273 1820 23307
rect 1768 23264 1820 23273
rect 9312 23307 9364 23316
rect 9312 23273 9321 23307
rect 9321 23273 9355 23307
rect 9355 23273 9364 23307
rect 9312 23264 9364 23273
rect 11336 23264 11388 23316
rect 13360 23264 13412 23316
rect 8484 23196 8536 23248
rect 2320 23060 2372 23112
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 5448 23103 5500 23112
rect 5448 23069 5457 23103
rect 5457 23069 5491 23103
rect 5491 23069 5500 23103
rect 5448 23060 5500 23069
rect 4620 22992 4672 23044
rect 4896 22992 4948 23044
rect 9404 23060 9456 23112
rect 9496 23060 9548 23112
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 11060 23196 11112 23248
rect 14188 23264 14240 23316
rect 14924 23264 14976 23316
rect 16304 23264 16356 23316
rect 16948 23264 17000 23316
rect 18052 23264 18104 23316
rect 18328 23264 18380 23316
rect 21272 23264 21324 23316
rect 22376 23264 22428 23316
rect 22560 23264 22612 23316
rect 24308 23264 24360 23316
rect 14648 23196 14700 23248
rect 16764 23196 16816 23248
rect 18696 23196 18748 23248
rect 23940 23196 23992 23248
rect 12072 23128 12124 23180
rect 13912 23128 13964 23180
rect 17776 23171 17828 23180
rect 17776 23137 17785 23171
rect 17785 23137 17819 23171
rect 17819 23137 17828 23171
rect 17776 23128 17828 23137
rect 17960 23128 18012 23180
rect 18972 23128 19024 23180
rect 19248 23128 19300 23180
rect 7656 22992 7708 23044
rect 8392 22992 8444 23044
rect 9312 22992 9364 23044
rect 14188 23060 14240 23112
rect 16672 23060 16724 23112
rect 16856 23060 16908 23112
rect 18052 23060 18104 23112
rect 21180 23128 21232 23180
rect 22284 23128 22336 23180
rect 23296 23128 23348 23180
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 25504 23060 25556 23112
rect 9404 22924 9456 22976
rect 15384 22924 15436 22976
rect 15476 22924 15528 22976
rect 17132 22992 17184 23044
rect 18328 22992 18380 23044
rect 18788 22992 18840 23044
rect 16764 22967 16816 22976
rect 16764 22933 16773 22967
rect 16773 22933 16807 22967
rect 16807 22933 16816 22967
rect 16764 22924 16816 22933
rect 17408 22924 17460 22976
rect 17684 22967 17736 22976
rect 17684 22933 17693 22967
rect 17693 22933 17727 22967
rect 17727 22933 17736 22967
rect 17684 22924 17736 22933
rect 18420 22924 18472 22976
rect 18696 22924 18748 22976
rect 19156 22924 19208 22976
rect 20260 22992 20312 23044
rect 21640 22992 21692 23044
rect 22192 22992 22244 23044
rect 23664 22992 23716 23044
rect 20996 22924 21048 22976
rect 22928 22924 22980 22976
rect 24124 22924 24176 22976
rect 24308 22924 24360 22976
rect 25596 22924 25648 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 4252 22652 4304 22704
rect 1400 22584 1452 22636
rect 1952 22584 2004 22636
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2780 22584 2832 22593
rect 9404 22720 9456 22772
rect 5724 22695 5776 22704
rect 5724 22661 5733 22695
rect 5733 22661 5767 22695
rect 5767 22661 5776 22695
rect 5724 22652 5776 22661
rect 6920 22695 6972 22704
rect 6920 22661 6929 22695
rect 6929 22661 6963 22695
rect 6963 22661 6972 22695
rect 6920 22652 6972 22661
rect 7104 22652 7156 22704
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 12348 22720 12400 22772
rect 14740 22720 14792 22772
rect 16304 22720 16356 22772
rect 16672 22720 16724 22772
rect 4160 22516 4212 22568
rect 4620 22448 4672 22500
rect 7656 22584 7708 22636
rect 11704 22652 11756 22704
rect 12164 22652 12216 22704
rect 13544 22652 13596 22704
rect 9036 22516 9088 22568
rect 12072 22516 12124 22568
rect 12256 22559 12308 22568
rect 12256 22525 12265 22559
rect 12265 22525 12299 22559
rect 12299 22525 12308 22559
rect 12256 22516 12308 22525
rect 2688 22380 2740 22432
rect 6000 22380 6052 22432
rect 9404 22380 9456 22432
rect 9680 22380 9732 22432
rect 11244 22380 11296 22432
rect 11520 22380 11572 22432
rect 13360 22584 13412 22636
rect 14188 22652 14240 22704
rect 14924 22652 14976 22704
rect 15660 22652 15712 22704
rect 16488 22652 16540 22704
rect 17224 22652 17276 22704
rect 19616 22720 19668 22772
rect 20260 22720 20312 22772
rect 21088 22763 21140 22772
rect 21088 22729 21097 22763
rect 21097 22729 21131 22763
rect 21131 22729 21140 22763
rect 21088 22720 21140 22729
rect 21640 22720 21692 22772
rect 22376 22720 22428 22772
rect 18604 22652 18656 22704
rect 22928 22652 22980 22704
rect 24308 22720 24360 22772
rect 24860 22720 24912 22772
rect 25228 22720 25280 22772
rect 23848 22652 23900 22704
rect 16764 22584 16816 22636
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 19432 22584 19484 22636
rect 22652 22584 22704 22636
rect 14556 22516 14608 22568
rect 14648 22516 14700 22568
rect 17776 22516 17828 22568
rect 19616 22516 19668 22568
rect 21364 22516 21416 22568
rect 14924 22448 14976 22500
rect 16488 22491 16540 22500
rect 16488 22457 16497 22491
rect 16497 22457 16531 22491
rect 16531 22457 16540 22491
rect 16488 22448 16540 22457
rect 16856 22448 16908 22500
rect 12716 22380 12768 22432
rect 13544 22380 13596 22432
rect 17132 22380 17184 22432
rect 17592 22380 17644 22432
rect 19708 22448 19760 22500
rect 22284 22559 22336 22568
rect 22284 22525 22293 22559
rect 22293 22525 22327 22559
rect 22327 22525 22336 22559
rect 22284 22516 22336 22525
rect 23296 22559 23348 22568
rect 23296 22525 23305 22559
rect 23305 22525 23339 22559
rect 23339 22525 23348 22559
rect 23296 22516 23348 22525
rect 24952 22516 25004 22568
rect 25228 22448 25280 22500
rect 19432 22380 19484 22432
rect 21456 22423 21508 22432
rect 21456 22389 21465 22423
rect 21465 22389 21499 22423
rect 21499 22389 21508 22423
rect 21456 22380 21508 22389
rect 22836 22380 22888 22432
rect 25412 22380 25464 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 2412 22176 2464 22228
rect 2964 22176 3016 22228
rect 13544 22176 13596 22228
rect 14740 22176 14792 22228
rect 14924 22176 14976 22228
rect 16212 22176 16264 22228
rect 2320 22108 2372 22160
rect 9772 22108 9824 22160
rect 12072 22108 12124 22160
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 3884 22040 3936 22092
rect 1768 21947 1820 21956
rect 1768 21913 1777 21947
rect 1777 21913 1811 21947
rect 1811 21913 1820 21947
rect 1768 21904 1820 21913
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 4528 21904 4580 21956
rect 6092 22083 6144 22092
rect 6092 22049 6101 22083
rect 6101 22049 6135 22083
rect 6135 22049 6144 22083
rect 6092 22040 6144 22049
rect 8300 22083 8352 22092
rect 8300 22049 8309 22083
rect 8309 22049 8343 22083
rect 8343 22049 8352 22083
rect 8300 22040 8352 22049
rect 9036 22040 9088 22092
rect 11060 22040 11112 22092
rect 12256 22040 12308 22092
rect 12716 22108 12768 22160
rect 13912 22108 13964 22160
rect 17224 22176 17276 22228
rect 18604 22176 18656 22228
rect 18972 22176 19024 22228
rect 20444 22176 20496 22228
rect 21180 22176 21232 22228
rect 7840 21972 7892 22024
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 9404 21904 9456 21956
rect 12900 21972 12952 22024
rect 13084 22015 13136 22024
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 13636 21972 13688 22024
rect 14188 21972 14240 22024
rect 9772 21904 9824 21956
rect 1952 21836 2004 21888
rect 4436 21836 4488 21888
rect 5540 21836 5592 21888
rect 6736 21836 6788 21888
rect 8392 21836 8444 21888
rect 9864 21836 9916 21888
rect 9956 21836 10008 21888
rect 11888 21836 11940 21888
rect 12900 21836 12952 21888
rect 13176 21904 13228 21956
rect 15844 21904 15896 21956
rect 13820 21836 13872 21888
rect 14096 21836 14148 21888
rect 17132 22083 17184 22092
rect 17132 22049 17141 22083
rect 17141 22049 17175 22083
rect 17175 22049 17184 22083
rect 17132 22040 17184 22049
rect 18144 22040 18196 22092
rect 19800 22108 19852 22160
rect 16764 21904 16816 21956
rect 17500 21972 17552 22024
rect 20720 22040 20772 22092
rect 19340 21972 19392 22024
rect 22652 22015 22704 22024
rect 22652 21981 22661 22015
rect 22661 21981 22695 22015
rect 22695 21981 22704 22015
rect 22652 21972 22704 21981
rect 24952 22015 25004 22024
rect 24952 21981 24961 22015
rect 24961 21981 24995 22015
rect 24995 21981 25004 22015
rect 24952 21972 25004 21981
rect 17132 21904 17184 21956
rect 16856 21879 16908 21888
rect 16856 21845 16865 21879
rect 16865 21845 16899 21879
rect 16899 21845 16908 21879
rect 16856 21836 16908 21845
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 17776 21836 17828 21888
rect 19156 21904 19208 21956
rect 19616 21904 19668 21956
rect 19708 21947 19760 21956
rect 19708 21913 19717 21947
rect 19717 21913 19751 21947
rect 19751 21913 19760 21947
rect 19708 21904 19760 21913
rect 21088 21904 21140 21956
rect 22192 21904 22244 21956
rect 23480 21904 23532 21956
rect 23848 21904 23900 21956
rect 24124 21904 24176 21956
rect 25228 21904 25280 21956
rect 18236 21836 18288 21888
rect 18972 21836 19024 21888
rect 20720 21836 20772 21888
rect 21272 21836 21324 21888
rect 21916 21836 21968 21888
rect 22376 21836 22428 21888
rect 22560 21836 22612 21888
rect 25412 21836 25464 21888
rect 26148 21836 26200 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 1584 21564 1636 21616
rect 9404 21564 9456 21616
rect 10324 21564 10376 21616
rect 3332 21496 3384 21548
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 10968 21632 11020 21684
rect 12716 21675 12768 21684
rect 12716 21641 12725 21675
rect 12725 21641 12759 21675
rect 12759 21641 12768 21675
rect 12716 21632 12768 21641
rect 13728 21632 13780 21684
rect 13912 21632 13964 21684
rect 16672 21632 16724 21684
rect 18512 21632 18564 21684
rect 20536 21632 20588 21684
rect 11152 21607 11204 21616
rect 11152 21573 11161 21607
rect 11161 21573 11195 21607
rect 11195 21573 11204 21607
rect 11152 21564 11204 21573
rect 13084 21564 13136 21616
rect 17684 21564 17736 21616
rect 20628 21564 20680 21616
rect 11888 21496 11940 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 7288 21428 7340 21480
rect 11244 21428 11296 21480
rect 11336 21428 11388 21480
rect 4068 21360 4120 21412
rect 4252 21360 4304 21412
rect 7012 21292 7064 21344
rect 10508 21292 10560 21344
rect 11704 21428 11756 21480
rect 12072 21428 12124 21480
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 12440 21360 12492 21412
rect 13176 21496 13228 21548
rect 15108 21496 15160 21548
rect 15200 21496 15252 21548
rect 13452 21428 13504 21480
rect 15568 21496 15620 21548
rect 15844 21496 15896 21548
rect 16304 21496 16356 21548
rect 17040 21496 17092 21548
rect 13912 21360 13964 21412
rect 15660 21471 15712 21480
rect 15660 21437 15669 21471
rect 15669 21437 15703 21471
rect 15703 21437 15712 21471
rect 15660 21428 15712 21437
rect 16488 21428 16540 21480
rect 16028 21360 16080 21412
rect 16304 21403 16356 21412
rect 16304 21369 16313 21403
rect 16313 21369 16347 21403
rect 16347 21369 16356 21403
rect 16304 21360 16356 21369
rect 16764 21403 16816 21412
rect 16764 21369 16773 21403
rect 16773 21369 16807 21403
rect 16807 21369 16816 21403
rect 16764 21360 16816 21369
rect 17132 21360 17184 21412
rect 17500 21539 17552 21548
rect 17500 21505 17509 21539
rect 17509 21505 17543 21539
rect 17543 21505 17552 21539
rect 17500 21496 17552 21505
rect 17316 21428 17368 21480
rect 17868 21360 17920 21412
rect 18972 21496 19024 21548
rect 18328 21428 18380 21480
rect 20904 21607 20956 21616
rect 20904 21573 20913 21607
rect 20913 21573 20947 21607
rect 20947 21573 20956 21607
rect 20904 21564 20956 21573
rect 21456 21564 21508 21616
rect 21732 21564 21784 21616
rect 23664 21632 23716 21684
rect 23848 21632 23900 21684
rect 24124 21564 24176 21616
rect 23296 21496 23348 21548
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 21732 21428 21784 21480
rect 21548 21403 21600 21412
rect 21548 21369 21557 21403
rect 21557 21369 21591 21403
rect 21591 21369 21600 21403
rect 21548 21360 21600 21369
rect 12532 21292 12584 21344
rect 12900 21292 12952 21344
rect 14740 21292 14792 21344
rect 14924 21292 14976 21344
rect 16212 21292 16264 21344
rect 17040 21335 17092 21344
rect 17040 21301 17049 21335
rect 17049 21301 17083 21335
rect 17083 21301 17092 21335
rect 17040 21292 17092 21301
rect 17500 21292 17552 21344
rect 19340 21292 19392 21344
rect 20260 21292 20312 21344
rect 24860 21428 24912 21480
rect 22836 21292 22888 21344
rect 23756 21292 23808 21344
rect 25412 21335 25464 21344
rect 25412 21301 25421 21335
rect 25421 21301 25455 21335
rect 25455 21301 25464 21335
rect 25412 21292 25464 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 2872 20995 2924 21004
rect 2872 20961 2881 20995
rect 2881 20961 2915 20995
rect 2915 20961 2924 20995
rect 2872 20952 2924 20961
rect 3332 21088 3384 21140
rect 8484 21020 8536 21072
rect 13544 21088 13596 21140
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 15200 21088 15252 21140
rect 16212 21088 16264 21140
rect 16672 21131 16724 21140
rect 16672 21097 16681 21131
rect 16681 21097 16715 21131
rect 16715 21097 16724 21131
rect 16672 21088 16724 21097
rect 17224 21088 17276 21140
rect 18420 21088 18472 21140
rect 18972 21131 19024 21140
rect 18972 21097 18981 21131
rect 18981 21097 19015 21131
rect 19015 21097 19024 21131
rect 18972 21088 19024 21097
rect 19524 21088 19576 21140
rect 21180 21131 21232 21140
rect 21180 21097 21189 21131
rect 21189 21097 21223 21131
rect 21223 21097 21232 21131
rect 21180 21088 21232 21097
rect 21364 21088 21416 21140
rect 4252 20952 4304 21004
rect 4344 20952 4396 21004
rect 6920 20952 6972 21004
rect 8760 20995 8812 21004
rect 8760 20961 8769 20995
rect 8769 20961 8803 20995
rect 8803 20961 8812 20995
rect 8760 20952 8812 20961
rect 18328 21020 18380 21072
rect 10508 20995 10560 21004
rect 10508 20961 10517 20995
rect 10517 20961 10551 20995
rect 10551 20961 10560 20995
rect 10508 20952 10560 20961
rect 11060 20952 11112 21004
rect 12072 20952 12124 21004
rect 12808 20952 12860 21004
rect 12900 20952 12952 21004
rect 16212 20952 16264 21004
rect 16396 20952 16448 21004
rect 4160 20927 4212 20936
rect 4160 20893 4169 20927
rect 4169 20893 4203 20927
rect 4203 20893 4212 20927
rect 4160 20884 4212 20893
rect 7012 20884 7064 20936
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 12532 20884 12584 20936
rect 12716 20884 12768 20936
rect 1952 20748 2004 20800
rect 2412 20748 2464 20800
rect 3056 20748 3108 20800
rect 5632 20748 5684 20800
rect 6460 20791 6512 20800
rect 6460 20757 6469 20791
rect 6469 20757 6503 20791
rect 6503 20757 6512 20791
rect 6460 20748 6512 20757
rect 6644 20816 6696 20868
rect 14004 20884 14056 20936
rect 14280 20884 14332 20936
rect 16304 20884 16356 20936
rect 17132 20884 17184 20936
rect 17408 20884 17460 20936
rect 21456 21020 21508 21072
rect 18696 20952 18748 21004
rect 21640 20952 21692 21004
rect 23480 20952 23532 21004
rect 24676 21020 24728 21072
rect 19340 20884 19392 20936
rect 24032 20884 24084 20936
rect 8300 20748 8352 20800
rect 9772 20748 9824 20800
rect 9956 20748 10008 20800
rect 10416 20748 10468 20800
rect 11244 20748 11296 20800
rect 12900 20748 12952 20800
rect 13176 20748 13228 20800
rect 15200 20816 15252 20868
rect 16764 20816 16816 20868
rect 17684 20816 17736 20868
rect 19984 20816 20036 20868
rect 21088 20816 21140 20868
rect 21272 20816 21324 20868
rect 23204 20859 23256 20868
rect 23204 20825 23213 20859
rect 23213 20825 23247 20859
rect 23247 20825 23256 20859
rect 23204 20816 23256 20825
rect 24584 20816 24636 20868
rect 14004 20748 14056 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 16028 20748 16080 20800
rect 21180 20748 21232 20800
rect 21456 20748 21508 20800
rect 21916 20748 21968 20800
rect 22008 20791 22060 20800
rect 22008 20757 22017 20791
rect 22017 20757 22051 20791
rect 22051 20757 22060 20791
rect 22008 20748 22060 20757
rect 23664 20748 23716 20800
rect 23848 20748 23900 20800
rect 24124 20748 24176 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 26056 20680 26108 20732
rect 26424 20680 26476 20732
rect 1676 20519 1728 20528
rect 1676 20485 1685 20519
rect 1685 20485 1719 20519
rect 1719 20485 1728 20519
rect 1676 20476 1728 20485
rect 7472 20544 7524 20596
rect 11520 20587 11572 20596
rect 3608 20476 3660 20528
rect 3056 20451 3108 20460
rect 3056 20417 3065 20451
rect 3065 20417 3099 20451
rect 3099 20417 3108 20451
rect 3056 20408 3108 20417
rect 8392 20476 8444 20528
rect 11520 20553 11529 20587
rect 11529 20553 11563 20587
rect 11563 20553 11572 20587
rect 11520 20544 11572 20553
rect 11704 20587 11756 20596
rect 11704 20553 11713 20587
rect 11713 20553 11747 20587
rect 11747 20553 11756 20587
rect 11704 20544 11756 20553
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 13176 20587 13228 20596
rect 9312 20476 9364 20528
rect 10600 20476 10652 20528
rect 11612 20476 11664 20528
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 10324 20408 10376 20460
rect 11888 20476 11940 20528
rect 13176 20553 13185 20587
rect 13185 20553 13219 20587
rect 13219 20553 13228 20587
rect 13176 20544 13228 20553
rect 13912 20544 13964 20596
rect 14740 20544 14792 20596
rect 14096 20476 14148 20528
rect 15476 20544 15528 20596
rect 17960 20544 18012 20596
rect 15200 20476 15252 20528
rect 16764 20476 16816 20528
rect 2596 20383 2648 20392
rect 2596 20349 2605 20383
rect 2605 20349 2639 20383
rect 2639 20349 2648 20383
rect 2596 20340 2648 20349
rect 3424 20383 3476 20392
rect 3424 20349 3433 20383
rect 3433 20349 3467 20383
rect 3467 20349 3476 20383
rect 3424 20340 3476 20349
rect 8944 20340 8996 20392
rect 10508 20340 10560 20392
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 20444 20544 20496 20596
rect 21088 20544 21140 20596
rect 21824 20544 21876 20596
rect 22008 20544 22060 20596
rect 23204 20544 23256 20596
rect 23388 20544 23440 20596
rect 23480 20544 23532 20596
rect 18604 20476 18656 20528
rect 19984 20476 20036 20528
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 4068 20204 4120 20256
rect 5356 20204 5408 20256
rect 6920 20204 6972 20256
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 11888 20204 11940 20256
rect 12440 20272 12492 20324
rect 13452 20340 13504 20392
rect 16028 20204 16080 20256
rect 16212 20247 16264 20256
rect 16212 20213 16221 20247
rect 16221 20213 16255 20247
rect 16255 20213 16264 20247
rect 16212 20204 16264 20213
rect 18328 20408 18380 20460
rect 23756 20519 23808 20528
rect 23756 20485 23765 20519
rect 23765 20485 23799 20519
rect 23799 20485 23808 20519
rect 23756 20476 23808 20485
rect 24032 20476 24084 20528
rect 23296 20408 23348 20460
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 17224 20340 17276 20349
rect 18236 20204 18288 20256
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 19892 20340 19944 20392
rect 19984 20340 20036 20392
rect 20720 20340 20772 20392
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 22652 20383 22704 20392
rect 22652 20349 22661 20383
rect 22661 20349 22695 20383
rect 22695 20349 22704 20383
rect 22652 20340 22704 20349
rect 21364 20272 21416 20324
rect 23848 20204 23900 20256
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 1400 20000 1452 20052
rect 1676 20043 1728 20052
rect 1676 20009 1685 20043
rect 1685 20009 1719 20043
rect 1719 20009 1728 20043
rect 1676 20000 1728 20009
rect 4160 20000 4212 20052
rect 6644 20043 6696 20052
rect 6644 20009 6653 20043
rect 6653 20009 6687 20043
rect 6687 20009 6696 20043
rect 6644 20000 6696 20009
rect 7288 20043 7340 20052
rect 7288 20009 7297 20043
rect 7297 20009 7331 20043
rect 7331 20009 7340 20043
rect 7288 20000 7340 20009
rect 9220 20000 9272 20052
rect 9312 20000 9364 20052
rect 10784 20000 10836 20052
rect 11152 20000 11204 20052
rect 16028 20000 16080 20052
rect 6828 19932 6880 19984
rect 8852 19932 8904 19984
rect 10600 19932 10652 19984
rect 4436 19864 4488 19916
rect 6092 19864 6144 19916
rect 4252 19839 4304 19848
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 6552 19796 6604 19848
rect 8944 19864 8996 19916
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 8760 19796 8812 19848
rect 9220 19796 9272 19848
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 12900 19932 12952 19984
rect 13728 19932 13780 19984
rect 14096 19932 14148 19984
rect 14464 19932 14516 19984
rect 16396 19932 16448 19984
rect 16672 19932 16724 19984
rect 18052 19932 18104 19984
rect 18788 19932 18840 19984
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 13544 19796 13596 19848
rect 13912 19796 13964 19848
rect 14648 19796 14700 19848
rect 15200 19796 15252 19848
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 17500 19864 17552 19916
rect 17592 19864 17644 19916
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 18696 19864 18748 19916
rect 19340 19864 19392 19916
rect 20720 20000 20772 20052
rect 23572 20000 23624 20052
rect 24216 20000 24268 20052
rect 22376 19932 22428 19984
rect 23296 19864 23348 19916
rect 24768 19864 24820 19916
rect 25044 19907 25096 19916
rect 25044 19873 25053 19907
rect 25053 19873 25087 19907
rect 25087 19873 25096 19907
rect 25044 19864 25096 19873
rect 20076 19796 20128 19848
rect 23388 19796 23440 19848
rect 2044 19728 2096 19780
rect 9496 19728 9548 19780
rect 11152 19728 11204 19780
rect 4436 19660 4488 19712
rect 6276 19660 6328 19712
rect 9128 19660 9180 19712
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10416 19660 10468 19669
rect 14464 19728 14516 19780
rect 14924 19728 14976 19780
rect 13912 19660 13964 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 15476 19728 15528 19780
rect 16672 19660 16724 19712
rect 16764 19660 16816 19712
rect 17960 19660 18012 19712
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 18236 19660 18288 19712
rect 18972 19660 19024 19712
rect 19340 19703 19392 19712
rect 19340 19669 19349 19703
rect 19349 19669 19383 19703
rect 19383 19669 19392 19703
rect 19340 19660 19392 19669
rect 20720 19728 20772 19780
rect 21364 19728 21416 19780
rect 20352 19660 20404 19712
rect 21640 19660 21692 19712
rect 23480 19660 23532 19712
rect 24124 19660 24176 19712
rect 24400 19660 24452 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 4528 19499 4580 19508
rect 4528 19465 4537 19499
rect 4537 19465 4571 19499
rect 4571 19465 4580 19499
rect 4528 19456 4580 19465
rect 6552 19499 6604 19508
rect 6552 19465 6561 19499
rect 6561 19465 6595 19499
rect 6595 19465 6604 19499
rect 6552 19456 6604 19465
rect 6736 19456 6788 19508
rect 9220 19456 9272 19508
rect 10968 19456 11020 19508
rect 11612 19456 11664 19508
rect 1584 19252 1636 19304
rect 1860 19252 1912 19304
rect 4160 19320 4212 19372
rect 3700 19252 3752 19304
rect 5172 19295 5224 19304
rect 5172 19261 5181 19295
rect 5181 19261 5215 19295
rect 5215 19261 5224 19295
rect 5172 19252 5224 19261
rect 7748 19388 7800 19440
rect 2780 19184 2832 19236
rect 4988 19184 5040 19236
rect 6552 19252 6604 19304
rect 6828 19252 6880 19304
rect 6276 19184 6328 19236
rect 8760 19388 8812 19440
rect 9312 19431 9364 19440
rect 9312 19397 9321 19431
rect 9321 19397 9355 19431
rect 9355 19397 9364 19431
rect 9312 19388 9364 19397
rect 8852 19320 8904 19372
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 11704 19320 11756 19372
rect 12164 19320 12216 19372
rect 13820 19456 13872 19508
rect 14464 19499 14516 19508
rect 14464 19465 14473 19499
rect 14473 19465 14507 19499
rect 14507 19465 14516 19499
rect 14464 19456 14516 19465
rect 14556 19456 14608 19508
rect 15476 19456 15528 19508
rect 16212 19456 16264 19508
rect 16764 19456 16816 19508
rect 17040 19456 17092 19508
rect 14280 19388 14332 19440
rect 18328 19388 18380 19440
rect 14096 19320 14148 19372
rect 14740 19320 14792 19372
rect 15108 19320 15160 19372
rect 16856 19320 16908 19372
rect 19524 19456 19576 19508
rect 20996 19456 21048 19508
rect 21180 19456 21232 19508
rect 23388 19456 23440 19508
rect 25136 19456 25188 19508
rect 25688 19456 25740 19508
rect 19892 19388 19944 19440
rect 20076 19388 20128 19440
rect 24032 19388 24084 19440
rect 19984 19320 20036 19372
rect 21088 19320 21140 19372
rect 22100 19320 22152 19372
rect 22192 19320 22244 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 7472 19252 7524 19304
rect 8392 19252 8444 19304
rect 10968 19252 11020 19304
rect 12532 19252 12584 19304
rect 13452 19252 13504 19304
rect 16028 19252 16080 19304
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 7288 19184 7340 19236
rect 3424 19116 3476 19168
rect 8852 19116 8904 19168
rect 10416 19184 10468 19236
rect 9864 19116 9916 19168
rect 10324 19116 10376 19168
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 12072 19159 12124 19168
rect 12072 19125 12081 19159
rect 12081 19125 12115 19159
rect 12115 19125 12124 19159
rect 12072 19116 12124 19125
rect 14096 19184 14148 19236
rect 14740 19184 14792 19236
rect 14924 19184 14976 19236
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 21364 19252 21416 19304
rect 22008 19252 22060 19304
rect 20168 19184 20220 19236
rect 13728 19116 13780 19168
rect 15660 19116 15712 19168
rect 18328 19116 18380 19168
rect 19248 19116 19300 19168
rect 19432 19116 19484 19168
rect 19984 19116 20036 19168
rect 20812 19184 20864 19236
rect 25228 19252 25280 19304
rect 21824 19116 21876 19168
rect 22008 19116 22060 19168
rect 25136 19116 25188 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 3884 18912 3936 18964
rect 2412 18844 2464 18896
rect 3792 18776 3844 18828
rect 7288 18912 7340 18964
rect 4988 18844 5040 18896
rect 5356 18844 5408 18896
rect 7840 18844 7892 18896
rect 10968 18844 11020 18896
rect 4896 18776 4948 18828
rect 5908 18776 5960 18828
rect 1492 18708 1544 18760
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 6552 18776 6604 18828
rect 9404 18776 9456 18828
rect 9588 18776 9640 18828
rect 14096 18912 14148 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 15568 18912 15620 18964
rect 16764 18912 16816 18964
rect 14740 18844 14792 18896
rect 2688 18640 2740 18692
rect 4344 18640 4396 18692
rect 10232 18708 10284 18760
rect 11704 18708 11756 18760
rect 14464 18776 14516 18828
rect 17224 18887 17276 18896
rect 17224 18853 17233 18887
rect 17233 18853 17267 18887
rect 17267 18853 17276 18887
rect 17224 18844 17276 18853
rect 17592 18887 17644 18896
rect 17592 18853 17601 18887
rect 17601 18853 17635 18887
rect 17635 18853 17644 18887
rect 17592 18844 17644 18853
rect 19064 18844 19116 18896
rect 19156 18844 19208 18896
rect 16948 18776 17000 18828
rect 18604 18819 18656 18828
rect 18604 18785 18613 18819
rect 18613 18785 18647 18819
rect 18647 18785 18656 18819
rect 18604 18776 18656 18785
rect 21824 18912 21876 18964
rect 22836 18912 22888 18964
rect 24676 18912 24728 18964
rect 23388 18844 23440 18896
rect 19800 18776 19852 18828
rect 21640 18776 21692 18828
rect 22468 18776 22520 18828
rect 8300 18640 8352 18692
rect 9496 18640 9548 18692
rect 13820 18708 13872 18760
rect 14924 18708 14976 18760
rect 19248 18708 19300 18760
rect 26056 18844 26108 18896
rect 25044 18776 25096 18828
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 13912 18640 13964 18692
rect 14556 18640 14608 18692
rect 15200 18640 15252 18692
rect 15660 18640 15712 18692
rect 16028 18640 16080 18692
rect 16212 18640 16264 18692
rect 17224 18640 17276 18692
rect 19156 18640 19208 18692
rect 19524 18683 19576 18692
rect 19524 18649 19533 18683
rect 19533 18649 19567 18683
rect 19567 18649 19576 18683
rect 19524 18640 19576 18649
rect 2136 18572 2188 18624
rect 5356 18572 5408 18624
rect 5816 18615 5868 18624
rect 5816 18581 5825 18615
rect 5825 18581 5859 18615
rect 5859 18581 5868 18615
rect 5816 18572 5868 18581
rect 5908 18572 5960 18624
rect 8392 18615 8444 18624
rect 8392 18581 8401 18615
rect 8401 18581 8435 18615
rect 8435 18581 8444 18615
rect 8392 18572 8444 18581
rect 8852 18572 8904 18624
rect 9864 18572 9916 18624
rect 10140 18572 10192 18624
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 12256 18572 12308 18624
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 15108 18572 15160 18624
rect 17776 18572 17828 18624
rect 20720 18640 20772 18692
rect 21364 18640 21416 18692
rect 19984 18572 20036 18624
rect 20996 18572 21048 18624
rect 21640 18572 21692 18624
rect 22192 18572 22244 18624
rect 22836 18640 22888 18692
rect 23204 18640 23256 18692
rect 25136 18708 25188 18760
rect 22744 18572 22796 18624
rect 24400 18615 24452 18624
rect 24400 18581 24409 18615
rect 24409 18581 24443 18615
rect 24443 18581 24452 18615
rect 24400 18572 24452 18581
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 24676 18572 24728 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 2872 18368 2924 18420
rect 5632 18368 5684 18420
rect 6184 18368 6236 18420
rect 7012 18368 7064 18420
rect 8300 18411 8352 18420
rect 8300 18377 8309 18411
rect 8309 18377 8343 18411
rect 8343 18377 8352 18411
rect 8300 18368 8352 18377
rect 8392 18368 8444 18420
rect 12532 18368 12584 18420
rect 13360 18368 13412 18420
rect 13820 18368 13872 18420
rect 14464 18368 14516 18420
rect 15476 18368 15528 18420
rect 4160 18300 4212 18352
rect 9220 18343 9272 18352
rect 9220 18309 9229 18343
rect 9229 18309 9263 18343
rect 9263 18309 9272 18343
rect 9220 18300 9272 18309
rect 10876 18300 10928 18352
rect 2044 18232 2096 18284
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 2780 18275 2832 18284
rect 2780 18241 2789 18275
rect 2789 18241 2823 18275
rect 2823 18241 2832 18275
rect 2780 18232 2832 18241
rect 4068 18275 4120 18284
rect 4068 18241 4077 18275
rect 4077 18241 4111 18275
rect 4111 18241 4120 18275
rect 4068 18232 4120 18241
rect 4344 18232 4396 18284
rect 4436 18164 4488 18216
rect 6368 18164 6420 18216
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8484 18275 8536 18284
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 10324 18232 10376 18284
rect 11060 18275 11112 18284
rect 11060 18241 11069 18275
rect 11069 18241 11103 18275
rect 11103 18241 11112 18275
rect 11060 18232 11112 18241
rect 11796 18232 11848 18284
rect 9772 18164 9824 18216
rect 9864 18164 9916 18216
rect 10508 18164 10560 18216
rect 10968 18164 11020 18216
rect 7196 18096 7248 18148
rect 7656 18139 7708 18148
rect 7656 18105 7665 18139
rect 7665 18105 7699 18139
rect 7699 18105 7708 18139
rect 7656 18096 7708 18105
rect 10232 18096 10284 18148
rect 3332 18028 3384 18080
rect 5816 18071 5868 18080
rect 5816 18037 5825 18071
rect 5825 18037 5859 18071
rect 5859 18037 5868 18071
rect 5816 18028 5868 18037
rect 9404 18028 9456 18080
rect 9772 18028 9824 18080
rect 10876 18028 10928 18080
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 14004 18232 14056 18284
rect 15660 18275 15712 18284
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 13084 18164 13136 18216
rect 15476 18164 15528 18216
rect 15844 18300 15896 18352
rect 18880 18300 18932 18352
rect 16212 18232 16264 18284
rect 16764 18232 16816 18284
rect 17500 18232 17552 18284
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 17960 18232 18012 18284
rect 12808 18028 12860 18080
rect 18236 18096 18288 18148
rect 17500 18028 17552 18080
rect 18512 18096 18564 18148
rect 19248 18071 19300 18080
rect 19248 18037 19257 18071
rect 19257 18037 19291 18071
rect 19291 18037 19300 18071
rect 19248 18028 19300 18037
rect 19984 18232 20036 18284
rect 19708 18207 19760 18216
rect 19708 18173 19717 18207
rect 19717 18173 19751 18207
rect 19751 18173 19760 18207
rect 19708 18164 19760 18173
rect 19892 18207 19944 18216
rect 19892 18173 19901 18207
rect 19901 18173 19935 18207
rect 19935 18173 19944 18207
rect 19892 18164 19944 18173
rect 20904 18207 20956 18216
rect 20904 18173 20913 18207
rect 20913 18173 20947 18207
rect 20947 18173 20956 18207
rect 20904 18164 20956 18173
rect 21088 18207 21140 18216
rect 21088 18173 21097 18207
rect 21097 18173 21131 18207
rect 21131 18173 21140 18207
rect 21088 18164 21140 18173
rect 21548 18411 21600 18420
rect 21548 18377 21557 18411
rect 21557 18377 21591 18411
rect 21591 18377 21600 18411
rect 21548 18368 21600 18377
rect 21640 18368 21692 18420
rect 22744 18368 22796 18420
rect 23296 18411 23348 18420
rect 22560 18300 22612 18352
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 23664 18368 23716 18420
rect 22928 18300 22980 18352
rect 23388 18232 23440 18284
rect 24400 18164 24452 18216
rect 25320 18164 25372 18216
rect 19984 18028 20036 18080
rect 20444 18071 20496 18080
rect 20444 18037 20453 18071
rect 20453 18037 20487 18071
rect 20487 18037 20496 18071
rect 20444 18028 20496 18037
rect 20720 18096 20772 18148
rect 21456 18028 21508 18080
rect 23388 18028 23440 18080
rect 23756 18028 23808 18080
rect 24032 18071 24084 18080
rect 24032 18037 24041 18071
rect 24041 18037 24075 18071
rect 24075 18037 24084 18071
rect 24032 18028 24084 18037
rect 24216 18071 24268 18080
rect 24216 18037 24225 18071
rect 24225 18037 24259 18071
rect 24259 18037 24268 18071
rect 24216 18028 24268 18037
rect 25044 18028 25096 18080
rect 25872 18028 25924 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 4068 17824 4120 17876
rect 4436 17824 4488 17876
rect 5540 17824 5592 17876
rect 7104 17824 7156 17876
rect 8392 17824 8444 17876
rect 8576 17824 8628 17876
rect 8668 17824 8720 17876
rect 14004 17824 14056 17876
rect 5356 17756 5408 17808
rect 13452 17756 13504 17808
rect 17592 17824 17644 17876
rect 17868 17824 17920 17876
rect 22192 17824 22244 17876
rect 22652 17824 22704 17876
rect 23020 17824 23072 17876
rect 24952 17824 25004 17876
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 5080 17688 5132 17740
rect 5448 17731 5500 17740
rect 5448 17697 5457 17731
rect 5457 17697 5491 17731
rect 5491 17697 5500 17731
rect 5448 17688 5500 17697
rect 8944 17688 8996 17740
rect 11704 17688 11756 17740
rect 12624 17688 12676 17740
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 15568 17688 15620 17740
rect 15936 17688 15988 17740
rect 16672 17688 16724 17740
rect 20076 17731 20128 17740
rect 20076 17697 20085 17731
rect 20085 17697 20119 17731
rect 20119 17697 20128 17731
rect 20076 17688 20128 17697
rect 22560 17688 22612 17740
rect 24124 17756 24176 17808
rect 4804 17620 4856 17672
rect 4988 17620 5040 17672
rect 6644 17663 6696 17672
rect 6644 17629 6653 17663
rect 6653 17629 6687 17663
rect 6687 17629 6696 17663
rect 6644 17620 6696 17629
rect 7012 17620 7064 17672
rect 7472 17620 7524 17672
rect 6736 17552 6788 17604
rect 2688 17484 2740 17536
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 5448 17484 5500 17536
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 9680 17620 9732 17672
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 9588 17552 9640 17604
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 10140 17552 10192 17604
rect 10324 17552 10376 17604
rect 12256 17552 12308 17604
rect 12716 17552 12768 17604
rect 11336 17484 11388 17536
rect 12440 17484 12492 17536
rect 12532 17484 12584 17536
rect 14004 17484 14056 17536
rect 15108 17552 15160 17604
rect 15476 17552 15528 17604
rect 15660 17552 15712 17604
rect 17408 17620 17460 17672
rect 17592 17620 17644 17672
rect 17040 17552 17092 17604
rect 17684 17552 17736 17604
rect 18604 17552 18656 17604
rect 17316 17484 17368 17536
rect 17776 17484 17828 17536
rect 18236 17484 18288 17536
rect 18880 17484 18932 17536
rect 19708 17484 19760 17536
rect 21640 17552 21692 17604
rect 22928 17688 22980 17740
rect 23572 17688 23624 17740
rect 25596 17688 25648 17740
rect 22836 17620 22888 17672
rect 23940 17620 23992 17672
rect 22744 17552 22796 17604
rect 22928 17484 22980 17536
rect 23756 17484 23808 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 1768 17280 1820 17332
rect 6552 17280 6604 17332
rect 7288 17280 7340 17332
rect 7380 17280 7432 17332
rect 8392 17280 8444 17332
rect 15936 17280 15988 17332
rect 17592 17280 17644 17332
rect 17776 17280 17828 17332
rect 19340 17280 19392 17332
rect 20260 17280 20312 17332
rect 22284 17323 22336 17332
rect 22284 17289 22293 17323
rect 22293 17289 22327 17323
rect 22327 17289 22336 17323
rect 22284 17280 22336 17289
rect 22376 17280 22428 17332
rect 23020 17280 23072 17332
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 3608 17212 3660 17264
rect 3332 17144 3384 17196
rect 4620 17144 4672 17196
rect 7564 17212 7616 17264
rect 7656 17212 7708 17264
rect 8484 17212 8536 17264
rect 9772 17212 9824 17264
rect 10140 17212 10192 17264
rect 6184 17144 6236 17196
rect 6920 17144 6972 17196
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 7748 17144 7800 17196
rect 7932 17144 7984 17196
rect 4160 17076 4212 17128
rect 5540 17076 5592 17128
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 8944 17144 8996 17196
rect 11060 17144 11112 17196
rect 12256 17212 12308 17264
rect 13452 17212 13504 17264
rect 17684 17212 17736 17264
rect 18604 17212 18656 17264
rect 22100 17212 22152 17264
rect 22836 17212 22888 17264
rect 22928 17212 22980 17264
rect 23664 17280 23716 17332
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 15292 17144 15344 17196
rect 10048 17076 10100 17128
rect 12440 17076 12492 17128
rect 12624 17076 12676 17128
rect 14096 17076 14148 17128
rect 8300 17008 8352 17060
rect 8668 17008 8720 17060
rect 11152 17008 11204 17060
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 7380 16940 7432 16992
rect 11612 16940 11664 16992
rect 15476 17076 15528 17128
rect 16948 17144 17000 17196
rect 17868 17144 17920 17196
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 22284 17144 22336 17196
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 24124 17280 24176 17332
rect 24216 17144 24268 17196
rect 13728 16983 13780 16992
rect 13728 16949 13737 16983
rect 13737 16949 13771 16983
rect 13771 16949 13780 16983
rect 13728 16940 13780 16949
rect 14280 16940 14332 16992
rect 14740 16940 14792 16992
rect 15108 16940 15160 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 19156 17076 19208 17128
rect 19616 17076 19668 17128
rect 21364 17076 21416 17128
rect 21640 17076 21692 17128
rect 22928 17076 22980 17128
rect 23572 17076 23624 17128
rect 20628 17008 20680 17060
rect 24124 17008 24176 17060
rect 24492 17008 24544 17060
rect 20168 16940 20220 16992
rect 20812 16940 20864 16992
rect 25688 17076 25740 17128
rect 26516 17008 26568 17060
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 6644 16736 6696 16788
rect 7288 16779 7340 16788
rect 7288 16745 7297 16779
rect 7297 16745 7331 16779
rect 7331 16745 7340 16779
rect 7288 16736 7340 16745
rect 3884 16643 3936 16652
rect 3884 16609 3893 16643
rect 3893 16609 3927 16643
rect 3927 16609 3936 16643
rect 3884 16600 3936 16609
rect 5908 16668 5960 16720
rect 7472 16668 7524 16720
rect 4712 16600 4764 16652
rect 7656 16668 7708 16720
rect 9036 16779 9088 16788
rect 9036 16745 9045 16779
rect 9045 16745 9079 16779
rect 9079 16745 9088 16779
rect 9036 16736 9088 16745
rect 9956 16736 10008 16788
rect 8300 16668 8352 16720
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 9496 16711 9548 16720
rect 9496 16677 9505 16711
rect 9505 16677 9539 16711
rect 9539 16677 9548 16711
rect 9496 16668 9548 16677
rect 1952 16439 2004 16448
rect 1952 16405 1961 16439
rect 1961 16405 1995 16439
rect 1995 16405 2004 16439
rect 1952 16396 2004 16405
rect 4160 16464 4212 16516
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 7564 16532 7616 16584
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 8392 16532 8444 16584
rect 8668 16532 8720 16584
rect 8852 16532 8904 16584
rect 10324 16668 10376 16720
rect 10600 16668 10652 16720
rect 15108 16736 15160 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 15660 16668 15712 16720
rect 19524 16736 19576 16788
rect 20168 16736 20220 16788
rect 20352 16736 20404 16788
rect 21456 16736 21508 16788
rect 10968 16532 11020 16584
rect 11612 16600 11664 16652
rect 12716 16600 12768 16652
rect 13728 16600 13780 16652
rect 14924 16600 14976 16652
rect 15752 16600 15804 16652
rect 11704 16532 11756 16584
rect 10600 16464 10652 16516
rect 12532 16464 12584 16516
rect 12716 16464 12768 16516
rect 14280 16464 14332 16516
rect 15016 16464 15068 16516
rect 19340 16600 19392 16652
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 22652 16600 22704 16652
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 23664 16532 23716 16584
rect 24860 16532 24912 16584
rect 25504 16532 25556 16584
rect 17316 16464 17368 16516
rect 17684 16464 17736 16516
rect 19340 16464 19392 16516
rect 5172 16396 5224 16448
rect 5632 16396 5684 16448
rect 11980 16396 12032 16448
rect 12348 16396 12400 16448
rect 13820 16396 13872 16448
rect 17224 16396 17276 16448
rect 19156 16396 19208 16448
rect 21364 16396 21416 16448
rect 21732 16396 21784 16448
rect 23940 16396 23992 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 3516 16192 3568 16244
rect 3884 16235 3936 16244
rect 3884 16201 3893 16235
rect 3893 16201 3927 16235
rect 3927 16201 3936 16235
rect 3884 16192 3936 16201
rect 5632 16192 5684 16244
rect 6276 16192 6328 16244
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 2136 16056 2188 16065
rect 3424 16056 3476 16108
rect 6460 16124 6512 16176
rect 6736 16192 6788 16244
rect 5264 16056 5316 16108
rect 8024 16099 8076 16108
rect 8024 16065 8033 16099
rect 8033 16065 8067 16099
rect 8067 16065 8076 16099
rect 8024 16056 8076 16065
rect 2228 15988 2280 16040
rect 2872 15920 2924 15972
rect 5356 15988 5408 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 7012 15988 7064 16040
rect 8484 16124 8536 16176
rect 10324 16192 10376 16244
rect 9036 16056 9088 16108
rect 11888 16124 11940 16176
rect 12716 16124 12768 16176
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 11520 16056 11572 16108
rect 7840 15963 7892 15972
rect 7840 15929 7849 15963
rect 7849 15929 7883 15963
rect 7883 15929 7892 15963
rect 7840 15920 7892 15929
rect 5540 15852 5592 15904
rect 6092 15852 6144 15904
rect 8300 15852 8352 15904
rect 8760 15852 8812 15904
rect 8944 15852 8996 15904
rect 10784 15920 10836 15972
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12348 15988 12400 16040
rect 20996 16192 21048 16244
rect 21916 16192 21968 16244
rect 22652 16192 22704 16244
rect 23848 16235 23900 16244
rect 23848 16201 23857 16235
rect 23857 16201 23891 16235
rect 23891 16201 23900 16235
rect 23848 16192 23900 16201
rect 13728 16124 13780 16176
rect 13544 16056 13596 16108
rect 15200 16056 15252 16108
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 11980 15852 12032 15904
rect 12348 15852 12400 15904
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 18788 16124 18840 16176
rect 19984 16124 20036 16176
rect 19616 16056 19668 16108
rect 18880 16031 18932 16040
rect 18880 15997 18889 16031
rect 18889 15997 18923 16031
rect 18923 15997 18932 16031
rect 18880 15988 18932 15997
rect 16488 15920 16540 15972
rect 21824 16056 21876 16108
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 20996 16031 21048 16040
rect 20996 15997 21005 16031
rect 21005 15997 21039 16031
rect 21039 15997 21048 16031
rect 20996 15988 21048 15997
rect 21272 15988 21324 16040
rect 24952 16124 25004 16176
rect 22744 16056 22796 16108
rect 22192 15988 22244 16040
rect 13360 15852 13412 15904
rect 14096 15852 14148 15904
rect 14188 15852 14240 15904
rect 14648 15852 14700 15904
rect 15292 15852 15344 15904
rect 16212 15852 16264 15904
rect 16396 15852 16448 15904
rect 19156 15852 19208 15904
rect 22560 15852 22612 15904
rect 23204 16056 23256 16108
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 23940 16031 23992 16040
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 23296 15895 23348 15904
rect 23296 15861 23305 15895
rect 23305 15861 23339 15895
rect 23339 15861 23348 15895
rect 23296 15852 23348 15861
rect 25228 15895 25280 15904
rect 25228 15861 25237 15895
rect 25237 15861 25271 15895
rect 25271 15861 25280 15895
rect 25228 15852 25280 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 2136 15648 2188 15700
rect 2596 15648 2648 15700
rect 4068 15648 4120 15700
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 8024 15691 8076 15700
rect 8024 15657 8033 15691
rect 8033 15657 8067 15691
rect 8067 15657 8076 15691
rect 8024 15648 8076 15657
rect 2872 15580 2924 15632
rect 5264 15580 5316 15632
rect 7380 15580 7432 15632
rect 8576 15648 8628 15700
rect 9312 15648 9364 15700
rect 4252 15444 4304 15496
rect 6920 15444 6972 15496
rect 7748 15444 7800 15496
rect 9864 15580 9916 15632
rect 11888 15580 11940 15632
rect 16856 15648 16908 15700
rect 17316 15648 17368 15700
rect 15568 15580 15620 15632
rect 16396 15623 16448 15632
rect 16396 15589 16405 15623
rect 16405 15589 16439 15623
rect 16439 15589 16448 15623
rect 16396 15580 16448 15589
rect 16580 15623 16632 15632
rect 16580 15589 16589 15623
rect 16589 15589 16623 15623
rect 16623 15589 16632 15623
rect 16580 15580 16632 15589
rect 18696 15691 18748 15700
rect 18696 15657 18705 15691
rect 18705 15657 18739 15691
rect 18739 15657 18748 15691
rect 18696 15648 18748 15657
rect 19892 15648 19944 15700
rect 22836 15580 22888 15632
rect 23388 15648 23440 15700
rect 24584 15580 24636 15632
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 4712 15351 4764 15360
rect 4712 15317 4721 15351
rect 4721 15317 4755 15351
rect 4755 15317 4764 15351
rect 4712 15308 4764 15317
rect 5908 15351 5960 15360
rect 5908 15317 5917 15351
rect 5917 15317 5951 15351
rect 5951 15317 5960 15351
rect 5908 15308 5960 15317
rect 9588 15376 9640 15428
rect 10692 15376 10744 15428
rect 10784 15419 10836 15428
rect 10784 15385 10793 15419
rect 10793 15385 10827 15419
rect 10827 15385 10836 15419
rect 10784 15376 10836 15385
rect 12348 15376 12400 15428
rect 12716 15376 12768 15428
rect 14188 15512 14240 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 16856 15512 16908 15564
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 21364 15555 21416 15564
rect 21364 15521 21373 15555
rect 21373 15521 21407 15555
rect 21407 15521 21416 15555
rect 21364 15512 21416 15521
rect 13820 15444 13872 15496
rect 13912 15444 13964 15496
rect 20536 15444 20588 15496
rect 10600 15308 10652 15360
rect 11612 15308 11664 15360
rect 14096 15308 14148 15360
rect 15016 15376 15068 15428
rect 16672 15376 16724 15428
rect 17316 15376 17368 15428
rect 17684 15376 17736 15428
rect 18604 15376 18656 15428
rect 21180 15376 21232 15428
rect 23296 15512 23348 15564
rect 22560 15444 22612 15496
rect 23388 15444 23440 15496
rect 25412 15444 25464 15496
rect 16028 15308 16080 15360
rect 19432 15308 19484 15360
rect 19524 15351 19576 15360
rect 19524 15317 19533 15351
rect 19533 15317 19567 15351
rect 19567 15317 19576 15351
rect 19524 15308 19576 15317
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 20904 15308 20956 15360
rect 22192 15308 22244 15360
rect 22376 15308 22428 15360
rect 22560 15351 22612 15360
rect 22560 15317 22569 15351
rect 22569 15317 22603 15351
rect 22603 15317 22612 15351
rect 22560 15308 22612 15317
rect 23572 15308 23624 15360
rect 25964 15308 26016 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 4252 15147 4304 15156
rect 4252 15113 4261 15147
rect 4261 15113 4295 15147
rect 4295 15113 4304 15147
rect 4252 15104 4304 15113
rect 4344 15104 4396 15156
rect 7012 15104 7064 15156
rect 10048 15104 10100 15156
rect 10416 15104 10468 15156
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 12624 15104 12676 15156
rect 13728 15104 13780 15156
rect 13820 15104 13872 15156
rect 16028 15104 16080 15156
rect 6920 15079 6972 15088
rect 6920 15045 6929 15079
rect 6929 15045 6963 15079
rect 6963 15045 6972 15079
rect 6920 15036 6972 15045
rect 9680 15079 9732 15088
rect 9680 15045 9689 15079
rect 9689 15045 9723 15079
rect 9723 15045 9732 15079
rect 9680 15036 9732 15045
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 9680 14832 9732 14884
rect 11888 15036 11940 15088
rect 12716 15036 12768 15088
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 13360 14968 13412 15020
rect 16764 15036 16816 15088
rect 18696 15104 18748 15156
rect 18880 15104 18932 15156
rect 21548 15147 21600 15156
rect 21548 15113 21557 15147
rect 21557 15113 21591 15147
rect 21591 15113 21600 15147
rect 21548 15104 21600 15113
rect 17224 15036 17276 15088
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 16580 14968 16632 15020
rect 10692 14900 10744 14952
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 11980 14900 12032 14952
rect 14740 14900 14792 14952
rect 16764 14900 16816 14952
rect 14464 14832 14516 14884
rect 16488 14832 16540 14884
rect 17132 14900 17184 14952
rect 17684 14900 17736 14952
rect 18604 14900 18656 14952
rect 19340 15036 19392 15088
rect 22376 15036 22428 15088
rect 23940 15104 23992 15156
rect 24768 15104 24820 15156
rect 23756 15036 23808 15088
rect 25136 15079 25188 15088
rect 25136 15045 25145 15079
rect 25145 15045 25179 15079
rect 25179 15045 25188 15079
rect 25136 15036 25188 15045
rect 19340 14943 19392 14952
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 20628 14900 20680 14952
rect 20812 14900 20864 14952
rect 22284 14900 22336 14952
rect 13820 14764 13872 14816
rect 15108 14764 15160 14816
rect 25596 14832 25648 14884
rect 18328 14764 18380 14816
rect 18696 14764 18748 14816
rect 20720 14764 20772 14816
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 25504 14764 25556 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 12440 14560 12492 14612
rect 18696 14560 18748 14612
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 19616 14560 19668 14612
rect 20260 14560 20312 14612
rect 13820 14492 13872 14544
rect 18512 14492 18564 14544
rect 18604 14492 18656 14544
rect 22100 14560 22152 14612
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 20720 14492 20772 14544
rect 22560 14492 22612 14544
rect 2688 14424 2740 14476
rect 5540 14424 5592 14476
rect 11612 14424 11664 14476
rect 12624 14424 12676 14476
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 15108 14424 15160 14476
rect 10416 14356 10468 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 12348 14356 12400 14408
rect 12716 14356 12768 14408
rect 13452 14356 13504 14408
rect 12256 14288 12308 14340
rect 14464 14288 14516 14340
rect 15016 14288 15068 14340
rect 18328 14424 18380 14476
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 22008 14424 22060 14476
rect 22744 14424 22796 14476
rect 23480 14424 23532 14476
rect 24308 14424 24360 14476
rect 13728 14220 13780 14272
rect 13820 14220 13872 14272
rect 14924 14220 14976 14272
rect 16672 14220 16724 14272
rect 17224 14288 17276 14340
rect 18052 14288 18104 14340
rect 20720 14356 20772 14408
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 21548 14356 21600 14408
rect 19432 14288 19484 14340
rect 24492 14356 24544 14408
rect 24860 14356 24912 14408
rect 23756 14288 23808 14340
rect 17776 14220 17828 14272
rect 18604 14220 18656 14272
rect 19248 14220 19300 14272
rect 20168 14220 20220 14272
rect 21088 14220 21140 14272
rect 21548 14220 21600 14272
rect 22744 14220 22796 14272
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 23664 14263 23716 14272
rect 23664 14229 23673 14263
rect 23673 14229 23707 14263
rect 23707 14229 23716 14263
rect 23664 14220 23716 14229
rect 23848 14220 23900 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 10508 14016 10560 14068
rect 10232 13948 10284 14000
rect 11612 14059 11664 14068
rect 11612 14025 11621 14059
rect 11621 14025 11655 14059
rect 11655 14025 11664 14059
rect 11612 14016 11664 14025
rect 12716 14016 12768 14068
rect 13360 14016 13412 14068
rect 9404 13880 9456 13932
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 12348 13880 12400 13932
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 14280 13948 14332 14000
rect 14464 13948 14516 14000
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 19340 14016 19392 14068
rect 20812 14016 20864 14068
rect 20996 14016 21048 14068
rect 17684 13948 17736 14000
rect 17776 13948 17828 14000
rect 9588 13744 9640 13796
rect 15016 13880 15068 13932
rect 17224 13880 17276 13932
rect 17868 13880 17920 13932
rect 18880 13948 18932 14000
rect 20444 13948 20496 14000
rect 22468 14016 22520 14068
rect 24768 14016 24820 14068
rect 23756 13948 23808 14000
rect 20720 13880 20772 13932
rect 21824 13880 21876 13932
rect 22192 13880 22244 13932
rect 22284 13880 22336 13932
rect 25136 13923 25188 13932
rect 25136 13889 25145 13923
rect 25145 13889 25179 13923
rect 25179 13889 25188 13923
rect 25136 13880 25188 13889
rect 25412 13880 25464 13932
rect 12716 13744 12768 13796
rect 13728 13744 13780 13796
rect 14556 13812 14608 13864
rect 16396 13812 16448 13864
rect 17592 13744 17644 13796
rect 19248 13812 19300 13864
rect 21180 13812 21232 13864
rect 20628 13744 20680 13796
rect 24308 13812 24360 13864
rect 25044 13812 25096 13864
rect 24216 13744 24268 13796
rect 24676 13744 24728 13796
rect 13360 13676 13412 13728
rect 13820 13676 13872 13728
rect 16028 13676 16080 13728
rect 16764 13676 16816 13728
rect 17408 13676 17460 13728
rect 19616 13676 19668 13728
rect 19984 13676 20036 13728
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 22192 13676 22244 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 13912 13515 13964 13524
rect 13912 13481 13921 13515
rect 13921 13481 13955 13515
rect 13955 13481 13964 13515
rect 13912 13472 13964 13481
rect 13360 13404 13412 13456
rect 15936 13472 15988 13524
rect 16028 13515 16080 13524
rect 16028 13481 16037 13515
rect 16037 13481 16071 13515
rect 16071 13481 16080 13515
rect 16028 13472 16080 13481
rect 19616 13472 19668 13524
rect 20168 13472 20220 13524
rect 20628 13472 20680 13524
rect 17776 13404 17828 13456
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 14556 13336 14608 13388
rect 15016 13336 15068 13388
rect 15108 13336 15160 13388
rect 16304 13336 16356 13388
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 18512 13336 18564 13388
rect 11244 13200 11296 13252
rect 10048 13132 10100 13184
rect 10692 13132 10744 13184
rect 18052 13268 18104 13320
rect 11980 13200 12032 13252
rect 12716 13200 12768 13252
rect 14188 13200 14240 13252
rect 14556 13243 14608 13252
rect 14556 13209 14565 13243
rect 14565 13209 14599 13243
rect 14599 13209 14608 13243
rect 14556 13200 14608 13209
rect 15016 13200 15068 13252
rect 13360 13132 13412 13184
rect 16764 13200 16816 13252
rect 17224 13200 17276 13252
rect 21088 13404 21140 13456
rect 19984 13336 20036 13388
rect 26056 13404 26108 13456
rect 25136 13379 25188 13388
rect 25136 13345 25145 13379
rect 25145 13345 25179 13379
rect 25179 13345 25188 13379
rect 25136 13336 25188 13345
rect 22100 13200 22152 13252
rect 22192 13243 22244 13252
rect 22192 13209 22201 13243
rect 22201 13209 22235 13243
rect 22235 13209 22244 13243
rect 22192 13200 22244 13209
rect 26056 13200 26108 13252
rect 16304 13132 16356 13184
rect 17592 13132 17644 13184
rect 18880 13132 18932 13184
rect 19064 13132 19116 13184
rect 23480 13132 23532 13184
rect 23756 13132 23808 13184
rect 24400 13132 24452 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 11244 12928 11296 12980
rect 11796 12928 11848 12980
rect 12716 12971 12768 12980
rect 12716 12937 12725 12971
rect 12725 12937 12759 12971
rect 12759 12937 12768 12971
rect 12716 12928 12768 12937
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 14280 12928 14332 12937
rect 17224 12860 17276 12912
rect 17776 12928 17828 12980
rect 18880 12928 18932 12980
rect 19800 12928 19852 12980
rect 22100 12928 22152 12980
rect 22192 12928 22244 12980
rect 25136 12928 25188 12980
rect 25228 12928 25280 12980
rect 12348 12835 12400 12844
rect 12348 12801 12357 12835
rect 12357 12801 12391 12835
rect 12391 12801 12400 12835
rect 12348 12792 12400 12801
rect 14372 12792 14424 12844
rect 16764 12792 16816 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 17500 12724 17552 12776
rect 18328 12724 18380 12776
rect 19156 12860 19208 12912
rect 19616 12860 19668 12912
rect 20536 12792 20588 12844
rect 18972 12724 19024 12776
rect 22376 12860 22428 12912
rect 22560 12860 22612 12912
rect 23388 12792 23440 12844
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 7288 12656 7340 12708
rect 18512 12656 18564 12708
rect 18604 12699 18656 12708
rect 18604 12665 18613 12699
rect 18613 12665 18647 12699
rect 18647 12665 18656 12699
rect 18604 12656 18656 12665
rect 20628 12656 20680 12708
rect 11336 12588 11388 12640
rect 19064 12631 19116 12640
rect 19064 12597 19073 12631
rect 19073 12597 19107 12631
rect 19107 12597 19116 12631
rect 19064 12588 19116 12597
rect 19432 12588 19484 12640
rect 19984 12588 20036 12640
rect 20352 12588 20404 12640
rect 20812 12588 20864 12640
rect 21364 12588 21416 12640
rect 24952 12588 25004 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 14464 12384 14516 12436
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 22100 12384 22152 12436
rect 22376 12384 22428 12436
rect 16764 12248 16816 12300
rect 17040 12248 17092 12300
rect 17224 12248 17276 12300
rect 20996 12248 21048 12300
rect 21364 12248 21416 12300
rect 22192 12248 22244 12300
rect 24308 12248 24360 12300
rect 5448 12180 5500 12232
rect 14372 12180 14424 12232
rect 15660 12180 15712 12232
rect 16304 12112 16356 12164
rect 16488 12112 16540 12164
rect 17040 12044 17092 12096
rect 19340 12180 19392 12232
rect 20812 12180 20864 12232
rect 18696 12155 18748 12164
rect 18696 12121 18705 12155
rect 18705 12121 18739 12155
rect 18739 12121 18748 12155
rect 18696 12112 18748 12121
rect 18880 12155 18932 12164
rect 18880 12121 18889 12155
rect 18889 12121 18923 12155
rect 18923 12121 18932 12155
rect 18880 12112 18932 12121
rect 19708 12155 19760 12164
rect 19708 12121 19717 12155
rect 19717 12121 19751 12155
rect 19751 12121 19760 12155
rect 19708 12112 19760 12121
rect 19984 12112 20036 12164
rect 21456 12180 21508 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 19800 12044 19852 12096
rect 20628 12044 20680 12096
rect 23388 12044 23440 12096
rect 24952 12044 25004 12096
rect 25228 12087 25280 12096
rect 25228 12053 25237 12087
rect 25237 12053 25271 12087
rect 25271 12053 25280 12087
rect 25228 12044 25280 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 5816 11772 5868 11824
rect 12716 11772 12768 11824
rect 14096 11840 14148 11892
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 13360 11772 13412 11824
rect 13820 11636 13872 11688
rect 14464 11772 14516 11824
rect 16488 11840 16540 11892
rect 15844 11815 15896 11824
rect 15844 11781 15853 11815
rect 15853 11781 15887 11815
rect 15887 11781 15896 11815
rect 15844 11772 15896 11781
rect 19340 11840 19392 11892
rect 21548 11840 21600 11892
rect 22192 11840 22244 11892
rect 22284 11840 22336 11892
rect 17316 11772 17368 11824
rect 19800 11772 19852 11824
rect 20996 11772 21048 11824
rect 24860 11772 24912 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 20812 11704 20864 11756
rect 21548 11704 21600 11756
rect 22284 11747 22336 11756
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22284 11704 22336 11713
rect 23940 11747 23992 11756
rect 23940 11713 23949 11747
rect 23949 11713 23983 11747
rect 23983 11713 23992 11747
rect 23940 11704 23992 11713
rect 12808 11500 12860 11552
rect 18604 11636 18656 11688
rect 18512 11568 18564 11620
rect 19156 11568 19208 11620
rect 22744 11568 22796 11620
rect 19708 11500 19760 11552
rect 19892 11500 19944 11552
rect 20352 11500 20404 11552
rect 21180 11543 21232 11552
rect 21180 11509 21189 11543
rect 21189 11509 21223 11543
rect 21223 11509 21232 11543
rect 21180 11500 21232 11509
rect 21548 11543 21600 11552
rect 21548 11509 21557 11543
rect 21557 11509 21591 11543
rect 21591 11509 21600 11543
rect 21548 11500 21600 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 14832 11296 14884 11348
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 16948 11296 17000 11348
rect 17408 11339 17460 11348
rect 17408 11305 17417 11339
rect 17417 11305 17451 11339
rect 17451 11305 17460 11339
rect 17408 11296 17460 11305
rect 18788 11296 18840 11348
rect 9128 11228 9180 11280
rect 18512 11228 18564 11280
rect 17868 11160 17920 11212
rect 15200 11092 15252 11144
rect 15752 11092 15804 11144
rect 16672 11092 16724 11144
rect 17132 11092 17184 11144
rect 19432 11296 19484 11348
rect 19156 11228 19208 11280
rect 17040 11024 17092 11076
rect 17960 11024 18012 11076
rect 18144 11024 18196 11076
rect 19340 11160 19392 11212
rect 19800 11160 19852 11212
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 20812 11160 20864 11212
rect 24860 11160 24912 11212
rect 25136 11160 25188 11212
rect 25412 11160 25464 11212
rect 14740 10956 14792 11008
rect 20168 11135 20220 11144
rect 20168 11101 20177 11135
rect 20177 11101 20211 11135
rect 20211 11101 20220 11135
rect 20168 11092 20220 11101
rect 20628 11092 20680 11144
rect 20996 11092 21048 11144
rect 22008 11092 22060 11144
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 24676 11092 24728 11144
rect 25320 11092 25372 11144
rect 20076 11024 20128 11076
rect 25412 11024 25464 11076
rect 19800 10956 19852 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 8760 10752 8812 10804
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 16672 10795 16724 10804
rect 16672 10761 16681 10795
rect 16681 10761 16715 10795
rect 16715 10761 16724 10795
rect 16672 10752 16724 10761
rect 17132 10752 17184 10804
rect 17592 10752 17644 10804
rect 17868 10752 17920 10804
rect 19432 10752 19484 10804
rect 20076 10795 20128 10804
rect 20076 10761 20085 10795
rect 20085 10761 20119 10795
rect 20119 10761 20128 10795
rect 20076 10752 20128 10761
rect 20168 10795 20220 10804
rect 20168 10761 20177 10795
rect 20177 10761 20211 10795
rect 20211 10761 20220 10795
rect 20168 10752 20220 10761
rect 20352 10752 20404 10804
rect 18236 10684 18288 10736
rect 16304 10659 16356 10668
rect 16304 10625 16313 10659
rect 16313 10625 16347 10659
rect 16347 10625 16356 10659
rect 16304 10616 16356 10625
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 14372 10548 14424 10600
rect 19156 10616 19208 10668
rect 19708 10548 19760 10600
rect 21272 10659 21324 10668
rect 21272 10625 21281 10659
rect 21281 10625 21315 10659
rect 21315 10625 21324 10659
rect 21272 10616 21324 10625
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 24860 10684 24912 10736
rect 24400 10548 24452 10600
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 13636 10480 13688 10532
rect 20812 10480 20864 10532
rect 21916 10480 21968 10532
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 15660 10208 15712 10260
rect 15016 10140 15068 10192
rect 19984 10208 20036 10260
rect 22652 10208 22704 10260
rect 18420 10072 18472 10124
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 19892 10072 19944 10124
rect 18328 9936 18380 9988
rect 18604 9936 18656 9988
rect 20076 10004 20128 10056
rect 20904 10072 20956 10124
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 22744 10140 22796 10192
rect 23296 10072 23348 10124
rect 23388 10072 23440 10124
rect 23480 10004 23532 10056
rect 24952 10004 25004 10056
rect 19156 9936 19208 9988
rect 20904 9936 20956 9988
rect 21180 9936 21232 9988
rect 19340 9868 19392 9920
rect 19432 9911 19484 9920
rect 19432 9877 19441 9911
rect 19441 9877 19475 9911
rect 19475 9877 19484 9911
rect 19432 9868 19484 9877
rect 19892 9868 19944 9920
rect 20168 9868 20220 9920
rect 24032 9979 24084 9988
rect 24032 9945 24041 9979
rect 24041 9945 24075 9979
rect 24075 9945 24084 9979
rect 24032 9936 24084 9945
rect 23388 9868 23440 9920
rect 24952 9911 25004 9920
rect 24952 9877 24961 9911
rect 24961 9877 24995 9911
rect 24995 9877 25004 9911
rect 24952 9868 25004 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 19432 9664 19484 9716
rect 16580 9528 16632 9580
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 17776 9528 17828 9580
rect 19156 9528 19208 9580
rect 20168 9596 20220 9648
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 20904 9528 20956 9580
rect 21088 9528 21140 9580
rect 21456 9571 21508 9580
rect 21456 9537 21465 9571
rect 21465 9537 21499 9571
rect 21499 9537 21508 9571
rect 21456 9528 21508 9537
rect 23296 9639 23348 9648
rect 23296 9605 23305 9639
rect 23305 9605 23339 9639
rect 23339 9605 23348 9639
rect 23296 9596 23348 9605
rect 26148 9596 26200 9648
rect 16028 9324 16080 9376
rect 19616 9392 19668 9444
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 19708 9324 19760 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 21456 9324 21508 9376
rect 26424 9324 26476 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 14464 9120 14516 9172
rect 17592 9120 17644 9172
rect 19432 9163 19484 9172
rect 19432 9129 19441 9163
rect 19441 9129 19475 9163
rect 19475 9129 19484 9163
rect 19432 9120 19484 9129
rect 20996 9120 21048 9172
rect 21548 9120 21600 9172
rect 23480 9120 23532 9172
rect 24584 9163 24636 9172
rect 24584 9129 24593 9163
rect 24593 9129 24627 9163
rect 24627 9129 24636 9163
rect 24584 9120 24636 9129
rect 25136 9120 25188 9172
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 19708 8984 19760 9036
rect 24952 9052 25004 9104
rect 18328 8959 18380 8968
rect 18328 8925 18337 8959
rect 18337 8925 18371 8959
rect 18371 8925 18380 8959
rect 18328 8916 18380 8925
rect 19984 8916 20036 8968
rect 21456 8984 21508 9036
rect 22008 8984 22060 9036
rect 24860 8984 24912 9036
rect 21088 8916 21140 8968
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 21548 8916 21600 8968
rect 9312 8848 9364 8900
rect 13820 8848 13872 8900
rect 24124 8848 24176 8900
rect 21548 8780 21600 8832
rect 22192 8780 22244 8832
rect 23480 8780 23532 8832
rect 26148 8780 26200 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 14004 8508 14056 8560
rect 19524 8440 19576 8492
rect 19984 8551 20036 8560
rect 19984 8517 19993 8551
rect 19993 8517 20027 8551
rect 20027 8517 20036 8551
rect 19984 8508 20036 8517
rect 20168 8551 20220 8560
rect 20168 8517 20177 8551
rect 20177 8517 20211 8551
rect 20211 8517 20220 8551
rect 20168 8508 20220 8517
rect 20536 8508 20588 8560
rect 20720 8440 20772 8492
rect 19156 8372 19208 8424
rect 21640 8372 21692 8424
rect 26516 8576 26568 8628
rect 24860 8508 24912 8560
rect 22192 8440 22244 8492
rect 22284 8372 22336 8424
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 20628 8347 20680 8356
rect 20628 8313 20637 8347
rect 20637 8313 20671 8347
rect 20671 8313 20680 8347
rect 20628 8304 20680 8313
rect 20904 8304 20956 8356
rect 25228 8304 25280 8356
rect 21640 8236 21692 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 15384 8032 15436 8084
rect 22192 8032 22244 8084
rect 24216 8032 24268 8084
rect 21364 7964 21416 8016
rect 16396 7896 16448 7948
rect 18972 7828 19024 7880
rect 19340 7828 19392 7880
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 21640 7828 21692 7880
rect 24492 8007 24544 8016
rect 24492 7973 24501 8007
rect 24501 7973 24535 8007
rect 24535 7973 24544 8007
rect 24492 7964 24544 7973
rect 24860 7896 24912 7948
rect 24676 7828 24728 7880
rect 19064 7760 19116 7812
rect 20352 7692 20404 7744
rect 20904 7692 20956 7744
rect 24952 7760 25004 7812
rect 25964 7760 26016 7812
rect 22008 7735 22060 7744
rect 22008 7701 22017 7735
rect 22017 7701 22051 7735
rect 22051 7701 22060 7735
rect 22008 7692 22060 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 6828 7488 6880 7540
rect 19248 7488 19300 7540
rect 25412 7488 25464 7540
rect 24860 7420 24912 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 20904 7352 20956 7404
rect 21732 7352 21784 7404
rect 21916 7352 21968 7404
rect 21180 7216 21232 7268
rect 21548 7284 21600 7336
rect 25412 7352 25464 7404
rect 26148 7352 26200 7404
rect 24676 7216 24728 7268
rect 25136 7216 25188 7268
rect 20076 7148 20128 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 21548 6944 21600 6996
rect 24584 6876 24636 6928
rect 25044 6876 25096 6928
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 22836 6740 22888 6792
rect 24952 6808 25004 6860
rect 25412 6808 25464 6860
rect 23940 6740 23992 6792
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 24860 6740 24912 6749
rect 20352 6672 20404 6724
rect 23296 6672 23348 6724
rect 24584 6672 24636 6724
rect 25688 6672 25740 6724
rect 17224 6604 17276 6656
rect 22836 6604 22888 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 23664 6400 23716 6452
rect 24860 6332 24912 6384
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 20444 6264 20496 6316
rect 22008 6264 22060 6316
rect 25872 6264 25924 6316
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 23480 6060 23532 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 22652 5856 22704 5908
rect 25320 5899 25372 5908
rect 25320 5865 25329 5899
rect 25329 5865 25363 5899
rect 25363 5865 25372 5899
rect 25320 5856 25372 5865
rect 19708 5788 19760 5840
rect 25780 5788 25832 5840
rect 21824 5720 21876 5772
rect 20628 5652 20680 5704
rect 22560 5652 22612 5704
rect 22836 5695 22888 5704
rect 22836 5661 22845 5695
rect 22845 5661 22879 5695
rect 22879 5661 22888 5695
rect 22836 5652 22888 5661
rect 24952 5652 25004 5704
rect 19616 5584 19668 5636
rect 25044 5584 25096 5636
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 21456 5312 21508 5364
rect 18328 5244 18380 5296
rect 19892 5176 19944 5228
rect 22468 5176 22520 5228
rect 24860 5244 24912 5296
rect 24676 5151 24728 5160
rect 24676 5117 24685 5151
rect 24685 5117 24719 5151
rect 24719 5117 24728 5151
rect 24676 5108 24728 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 8668 4768 8720 4820
rect 25136 4811 25188 4820
rect 25136 4777 25145 4811
rect 25145 4777 25179 4811
rect 25179 4777 25188 4811
rect 25136 4768 25188 4777
rect 24584 4700 24636 4752
rect 24676 4743 24728 4752
rect 24676 4709 24685 4743
rect 24685 4709 24719 4743
rect 24719 4709 24728 4743
rect 24676 4700 24728 4709
rect 7012 4564 7064 4616
rect 22744 4632 22796 4684
rect 25596 4632 25648 4684
rect 21180 4496 21232 4548
rect 24952 4496 25004 4548
rect 26056 4428 26108 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 22100 4020 22152 4072
rect 23204 4020 23256 4072
rect 25044 4088 25096 4140
rect 25504 4088 25556 4140
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 24952 3952 25004 4004
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 23480 3544 23532 3596
rect 7472 3476 7524 3528
rect 19800 3476 19852 3528
rect 24676 3476 24728 3528
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 24952 3408 25004 3460
rect 7196 3340 7248 3392
rect 22284 3340 22336 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 25964 3136 26016 3188
rect 6736 3000 6788 3052
rect 24860 3068 24912 3120
rect 25136 3111 25188 3120
rect 25136 3077 25145 3111
rect 25145 3077 25179 3111
rect 25179 3077 25188 3111
rect 25136 3068 25188 3077
rect 18880 3000 18932 3052
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 24032 3043 24084 3052
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 25044 2932 25096 2984
rect 6736 2796 6788 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 7012 2592 7064 2644
rect 19340 2592 19392 2644
rect 22836 2592 22888 2644
rect 23388 2592 23440 2644
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 23388 2456 23440 2508
rect 24584 2388 24636 2440
rect 24952 2320 25004 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1674 26200 1730 27000
rect 1952 26376 2004 26382
rect 1952 26318 2004 26324
rect 1582 25936 1638 25945
rect 1582 25871 1638 25880
rect 1490 23760 1546 23769
rect 1490 23695 1546 23704
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 20058 1440 22578
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1504 18766 1532 23695
rect 1596 21622 1624 25871
rect 1688 22794 1716 26200
rect 1766 23760 1822 23769
rect 1766 23695 1822 23704
rect 1860 23724 1912 23730
rect 1780 23322 1808 23695
rect 1860 23666 1912 23672
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1872 23089 1900 23666
rect 1858 23080 1914 23089
rect 1858 23015 1914 23024
rect 1688 22766 1900 22794
rect 1674 22672 1730 22681
rect 1674 22607 1730 22616
rect 1584 21616 1636 21622
rect 1584 21558 1636 21564
rect 1596 19310 1624 21558
rect 1688 20534 1716 22607
rect 1766 21992 1822 22001
rect 1766 21927 1768 21936
rect 1820 21927 1822 21936
rect 1768 21898 1820 21904
rect 1766 21448 1822 21457
rect 1766 21383 1822 21392
rect 1676 20528 1728 20534
rect 1676 20470 1728 20476
rect 1688 20058 1716 20470
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1780 17338 1808 21383
rect 1872 19310 1900 22766
rect 1964 22642 1992 26318
rect 2042 26200 2098 27000
rect 2410 26200 2466 27000
rect 2778 26466 2834 27000
rect 2778 26450 3096 26466
rect 2778 26444 3108 26450
rect 2778 26438 3056 26444
rect 2778 26200 2834 26438
rect 3056 26386 3108 26392
rect 3146 26330 3202 27000
rect 3424 26444 3476 26450
rect 3424 26386 3476 26392
rect 2884 26302 3202 26330
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1952 21888 2004 21894
rect 1952 21830 2004 21836
rect 1964 20806 1992 21830
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 2056 19786 2084 26200
rect 2228 23520 2280 23526
rect 2228 23462 2280 23468
rect 2134 23080 2190 23089
rect 2134 23015 2190 23024
rect 2044 19780 2096 19786
rect 2044 19722 2096 19728
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2148 18986 2176 23015
rect 2056 18958 2176 18986
rect 2056 18290 2084 18958
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2148 18290 2176 18566
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 1950 17776 2006 17785
rect 1950 17711 1952 17720
rect 2004 17711 2006 17720
rect 1952 17682 2004 17688
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 2134 17232 2190 17241
rect 2134 17167 2136 17176
rect 2188 17167 2190 17176
rect 2136 17138 2188 17144
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 13433 1992 16390
rect 2134 16144 2190 16153
rect 2134 16079 2136 16088
rect 2188 16079 2190 16088
rect 2136 16050 2188 16056
rect 2148 15706 2176 16050
rect 2240 16046 2268 23462
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2332 22166 2360 23054
rect 2424 22234 2452 26200
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2688 22432 2740 22438
rect 2688 22374 2740 22380
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2320 22160 2372 22166
rect 2320 22102 2372 22108
rect 2412 20800 2464 20806
rect 2412 20742 2464 20748
rect 2424 20262 2452 20742
rect 2596 20392 2648 20398
rect 2594 20360 2596 20369
rect 2648 20360 2650 20369
rect 2594 20295 2650 20304
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 18902 2452 20198
rect 2412 18896 2464 18902
rect 2412 18838 2464 18844
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2608 15706 2636 18702
rect 2700 18698 2728 22374
rect 2792 19394 2820 22578
rect 2884 22098 2912 26302
rect 3146 26200 3202 26302
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2976 21434 3004 22170
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 2884 21406 3004 21434
rect 2884 21010 2912 21406
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 3344 21146 3372 21490
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 3068 20466 3096 20742
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 3436 20398 3464 26386
rect 3514 26200 3570 27000
rect 3882 26330 3938 27000
rect 3882 26302 4108 26330
rect 3882 26200 3938 26302
rect 3528 21486 3556 26200
rect 3700 24880 3752 24886
rect 3606 24848 3662 24857
rect 3700 24822 3752 24828
rect 3606 24783 3662 24792
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3620 20534 3648 24783
rect 3608 20528 3660 20534
rect 3608 20470 3660 20476
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3606 20224 3662 20233
rect 2950 20156 3258 20165
rect 3606 20159 3662 20168
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2792 19366 2912 19394
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2792 18290 2820 19178
rect 2884 18426 2912 19366
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3238 17640 3294 17649
rect 3238 17575 3294 17584
rect 3252 17542 3280 17575
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2700 14482 2728 17478
rect 3344 17202 3372 18022
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 2792 16590 2820 17031
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 3436 16114 3464 19110
rect 3514 19000 3570 19009
rect 3514 18935 3570 18944
rect 3528 16250 3556 18935
rect 3620 17270 3648 20159
rect 3712 19310 3740 24822
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3804 18834 3832 23802
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3884 22092 3936 22098
rect 3884 22034 3936 22040
rect 3896 18970 3924 22034
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 3608 17264 3660 17270
rect 3608 17206 3660 17212
rect 3882 16688 3938 16697
rect 3882 16623 3884 16632
rect 3936 16623 3938 16632
rect 3884 16594 3936 16600
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2884 15638 2912 15914
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 3896 14929 3924 16186
rect 3988 15688 4016 23054
rect 4080 22094 4108 26302
rect 4250 26200 4306 27000
rect 4618 26200 4674 27000
rect 4986 26330 5042 27000
rect 5354 26330 5410 27000
rect 4986 26302 5120 26330
rect 4986 26200 5042 26302
rect 4160 24676 4212 24682
rect 4160 24618 4212 24624
rect 4172 24206 4200 24618
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 4172 22574 4200 23666
rect 4264 22710 4292 26200
rect 4632 23050 4660 26200
rect 4802 25664 4858 25673
rect 4802 25599 4858 25608
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4620 22500 4672 22506
rect 4620 22442 4672 22448
rect 4080 22066 4384 22094
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4264 21418 4292 21966
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 4252 21412 4304 21418
rect 4252 21354 4304 21360
rect 4080 20262 4108 21354
rect 4264 21010 4292 21354
rect 4356 21010 4384 22066
rect 4528 21956 4580 21962
rect 4528 21898 4580 21904
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4344 21004 4396 21010
rect 4344 20946 4396 20952
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4172 20058 4200 20878
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4448 19922 4476 21830
rect 4436 19916 4488 19922
rect 4436 19858 4488 19864
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4172 18358 4200 19314
rect 4160 18352 4212 18358
rect 4066 18320 4122 18329
rect 4160 18294 4212 18300
rect 4066 18255 4068 18264
rect 4120 18255 4122 18264
rect 4068 18226 4120 18232
rect 4080 17882 4108 18226
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4172 16522 4200 17070
rect 4264 16946 4292 19790
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4356 18290 4384 18634
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4448 18222 4476 19654
rect 4540 19514 4568 21898
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 4448 17882 4476 18158
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4632 17202 4660 22442
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4264 16918 4384 16946
rect 4250 16824 4306 16833
rect 4250 16759 4306 16768
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4068 15700 4120 15706
rect 3988 15660 4068 15688
rect 4068 15642 4120 15648
rect 4264 15502 4292 16759
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4264 15162 4292 15438
rect 4356 15162 4384 16918
rect 4724 16658 4752 24278
rect 4816 24206 4844 25599
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4988 24064 5040 24070
rect 4988 24006 5040 24012
rect 4896 23044 4948 23050
rect 4896 22986 4948 22992
rect 4802 21584 4858 21593
rect 4802 21519 4804 21528
rect 4856 21519 4858 21528
rect 4804 21490 4856 21496
rect 4908 18834 4936 22986
rect 5000 19242 5028 24006
rect 5092 21486 5120 26302
rect 5184 26302 5410 26330
rect 5184 23798 5212 26302
rect 5354 26200 5410 26302
rect 5722 26200 5778 27000
rect 6090 26200 6146 27000
rect 6458 26200 6514 27000
rect 6826 26200 6882 27000
rect 7194 26330 7250 27000
rect 7562 26330 7618 27000
rect 7930 26330 7986 27000
rect 7194 26302 7328 26330
rect 7194 26200 7250 26302
rect 5356 24336 5408 24342
rect 5356 24278 5408 24284
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5172 23792 5224 23798
rect 5172 23734 5224 23740
rect 5172 23588 5224 23594
rect 5172 23530 5224 23536
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5184 19938 5212 23530
rect 5092 19910 5212 19938
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4988 18896 5040 18902
rect 4986 18864 4988 18873
rect 5040 18864 5042 18873
rect 4896 18828 4948 18834
rect 4986 18799 5042 18808
rect 4896 18770 4948 18776
rect 4986 18048 5042 18057
rect 4986 17983 5042 17992
rect 4802 17776 4858 17785
rect 4802 17711 4858 17720
rect 4816 17678 4844 17711
rect 5000 17678 5028 17983
rect 5092 17746 5120 19910
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 5184 16454 5212 19246
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5276 16114 5304 24142
rect 5368 22094 5396 24278
rect 5632 24132 5684 24138
rect 5632 24074 5684 24080
rect 5644 23730 5672 24074
rect 5632 23724 5684 23730
rect 5632 23666 5684 23672
rect 5446 23216 5502 23225
rect 5446 23151 5502 23160
rect 5460 23118 5488 23151
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5736 22710 5764 26200
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 5538 22536 5594 22545
rect 5538 22471 5594 22480
rect 5368 22066 5488 22094
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 19961 5396 20198
rect 5354 19952 5410 19961
rect 5354 19887 5410 19896
rect 5356 18896 5408 18902
rect 5356 18838 5408 18844
rect 5368 18630 5396 18838
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5368 16046 5396 17750
rect 5460 17746 5488 22066
rect 5552 21978 5580 22471
rect 5828 22094 5856 24550
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 5736 22066 5856 22094
rect 5552 21950 5672 21978
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5552 17882 5580 21830
rect 5644 20806 5672 21950
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5630 19272 5686 19281
rect 5630 19207 5686 19216
rect 5644 18426 5672 19207
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 15632 5316 15638
rect 5262 15600 5264 15609
rect 5316 15600 5318 15609
rect 5262 15535 5318 15544
rect 4710 15464 4766 15473
rect 4710 15399 4766 15408
rect 4724 15366 4752 15399
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 3882 14920 3938 14929
rect 3882 14855 3938 14864
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 1950 13424 2006 13433
rect 1950 13359 2006 13368
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 5460 12238 5488 17478
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 15910 5580 17070
rect 5736 16833 5764 22066
rect 6012 19334 6040 22374
rect 6104 22098 6132 26200
rect 6182 26072 6238 26081
rect 6182 26007 6238 26016
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 5920 19306 6040 19334
rect 5920 18834 5948 19306
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5814 18728 5870 18737
rect 5814 18663 5870 18672
rect 5828 18630 5856 18663
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5722 16824 5778 16833
rect 5722 16759 5778 16768
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5644 16250 5672 16390
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5448 12232 5500 12238
rect 5552 12209 5580 14418
rect 5448 12174 5500 12180
rect 5538 12200 5594 12209
rect 5538 12135 5594 12144
rect 5828 11830 5856 18022
rect 5920 16726 5948 18566
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 6104 15910 6132 19858
rect 6196 18426 6224 26007
rect 6274 24304 6330 24313
rect 6472 24274 6500 26200
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6274 24239 6330 24248
rect 6460 24268 6512 24274
rect 6288 19718 6316 24239
rect 6460 24210 6512 24216
rect 6748 24206 6776 24346
rect 6736 24200 6788 24206
rect 6734 24168 6736 24177
rect 6788 24168 6790 24177
rect 6734 24103 6790 24112
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6564 23497 6592 24006
rect 6550 23488 6606 23497
rect 6550 23423 6606 23432
rect 6840 22094 6868 26200
rect 7010 24168 7066 24177
rect 7010 24103 7066 24112
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6932 22710 6960 23462
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 6840 22066 6960 22094
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6366 21312 6422 21321
rect 6366 21247 6422 21256
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 6276 19236 6328 19242
rect 6276 19178 6328 19184
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6196 17202 6224 18362
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6288 16250 6316 19178
rect 6380 18222 6408 21247
rect 6644 20868 6696 20874
rect 6644 20810 6696 20816
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6472 16182 6500 20742
rect 6656 20058 6684 20810
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6564 19514 6592 19790
rect 6748 19666 6776 21830
rect 6932 21010 6960 22066
rect 7024 21350 7052 24103
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7024 20942 7052 21286
rect 7116 21026 7144 22646
rect 7300 21486 7328 26302
rect 7392 26302 7618 26330
rect 7392 23798 7420 26302
rect 7562 26200 7618 26302
rect 7668 26302 7986 26330
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 7116 20998 7236 21026
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 6826 20360 6882 20369
rect 6826 20295 6882 20304
rect 6840 19990 6868 20295
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6828 19984 6880 19990
rect 6828 19926 6880 19932
rect 6656 19638 6776 19666
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6564 18834 6592 19246
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6656 17762 6684 19638
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6564 17734 6684 17762
rect 6564 17338 6592 17734
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5920 14521 5948 15302
rect 5906 14512 5962 14521
rect 5906 14447 5962 14456
rect 6564 13977 6592 16934
rect 6656 16794 6684 17614
rect 6748 17610 6776 19450
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6840 17082 6868 19246
rect 6932 17202 6960 20198
rect 7010 19408 7066 19417
rect 7010 19343 7066 19352
rect 7024 18426 7052 19343
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7024 17678 7052 18362
rect 7116 17882 7144 20878
rect 7208 19938 7236 20998
rect 7286 20088 7342 20097
rect 7286 20023 7288 20032
rect 7340 20023 7342 20032
rect 7288 19994 7340 20000
rect 7208 19910 7328 19938
rect 7194 19816 7250 19825
rect 7194 19751 7250 19760
rect 7208 18154 7236 19751
rect 7300 19553 7328 19910
rect 7286 19544 7342 19553
rect 7286 19479 7342 19488
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 7300 18970 7328 19178
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 7392 18034 7420 21490
rect 7484 20602 7512 24686
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7484 19854 7512 20538
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7300 18006 7420 18034
rect 7104 17876 7156 17882
rect 7300 17864 7328 18006
rect 7300 17836 7420 17864
rect 7104 17818 7156 17824
rect 7286 17776 7342 17785
rect 7286 17711 7342 17720
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6840 17054 7052 17082
rect 6918 16824 6974 16833
rect 6644 16788 6696 16794
rect 6918 16759 6974 16768
rect 6644 16730 6696 16736
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6748 16250 6776 16526
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6550 13968 6606 13977
rect 6550 13903 6606 13912
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 6840 7546 6868 15982
rect 6932 15502 6960 16759
rect 7024 16046 7052 17054
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6932 15094 6960 15438
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 7024 11801 7052 15098
rect 7116 13705 7144 17478
rect 7300 17338 7328 17711
rect 7392 17338 7420 17836
rect 7484 17785 7512 19246
rect 7470 17776 7526 17785
rect 7470 17711 7526 17720
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7392 16998 7420 17138
rect 7380 16992 7432 16998
rect 7286 16960 7342 16969
rect 7380 16934 7432 16940
rect 7286 16895 7342 16904
rect 7300 16794 7328 16895
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7286 16008 7342 16017
rect 7286 15943 7342 15952
rect 7102 13696 7158 13705
rect 7102 13631 7158 13640
rect 7300 12714 7328 15943
rect 7392 15638 7420 16934
rect 7484 16726 7512 17614
rect 7576 17270 7604 23666
rect 7668 23050 7696 26302
rect 7930 26200 7986 26302
rect 8298 26200 8354 27000
rect 8666 26330 8722 27000
rect 9034 26330 9090 27000
rect 8404 26302 8722 26330
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 7656 23044 7708 23050
rect 7656 22986 7708 22992
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7668 18272 7696 22578
rect 7760 19446 7788 24142
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8312 22098 8340 26200
rect 8404 24138 8432 26302
rect 8666 26200 8722 26302
rect 8772 26302 9090 26330
rect 8666 25936 8722 25945
rect 8666 25871 8722 25880
rect 8392 24132 8444 24138
rect 8392 24074 8444 24080
rect 8576 24132 8628 24138
rect 8576 24074 8628 24080
rect 8484 23248 8536 23254
rect 8484 23190 8536 23196
rect 8392 23044 8444 23050
rect 8392 22986 8444 22992
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7852 20913 7880 21966
rect 8404 21894 8432 22986
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8496 21162 8524 23190
rect 8404 21134 8524 21162
rect 8298 21040 8354 21049
rect 8298 20975 8354 20984
rect 7838 20904 7894 20913
rect 7838 20839 7894 20848
rect 8312 20806 8340 20975
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8404 20534 8432 21134
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8390 19544 8446 19553
rect 8390 19479 8446 19488
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 8404 19310 8432 19479
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7852 18290 7880 18838
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8312 18426 8340 18634
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18426 8432 18566
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8496 18290 8524 21014
rect 7840 18284 7892 18290
rect 7668 18244 7788 18272
rect 7654 18184 7710 18193
rect 7654 18119 7656 18128
rect 7708 18119 7710 18128
rect 7656 18090 7708 18096
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7668 16946 7696 17206
rect 7760 17202 7788 18244
rect 7840 18226 7892 18232
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8588 18170 8616 24074
rect 8404 18142 8616 18170
rect 7838 17912 7894 17921
rect 8404 17882 8432 18142
rect 8680 18068 8708 25871
rect 8772 22710 8800 26302
rect 9034 26200 9090 26302
rect 9402 26200 9458 27000
rect 9770 26330 9826 27000
rect 9692 26302 9826 26330
rect 9218 24712 9274 24721
rect 9218 24647 9274 24656
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 9126 22672 9182 22681
rect 9126 22607 9182 22616
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 9048 22098 9076 22510
rect 9036 22092 9088 22098
rect 9036 22034 9088 22040
rect 9048 21554 9076 22034
rect 9140 22030 9168 22607
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8758 21448 8814 21457
rect 8758 21383 8814 21392
rect 8772 21010 8800 21383
rect 8760 21004 8812 21010
rect 8760 20946 8812 20952
rect 8772 19854 8800 20946
rect 9048 20466 9076 21490
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8496 18040 8708 18068
rect 7838 17847 7894 17856
rect 8392 17876 8444 17882
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7576 16918 7696 16946
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7576 16590 7604 16918
rect 7656 16720 7708 16726
rect 7760 16708 7788 17138
rect 7708 16680 7788 16708
rect 7656 16662 7708 16668
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7852 16266 7880 17847
rect 8392 17818 8444 17824
rect 8298 17776 8354 17785
rect 8298 17711 8354 17720
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7944 16590 7972 17138
rect 8312 17066 8340 17711
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8404 17338 8432 17478
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8496 17270 8524 18040
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 7932 16584 7984 16590
rect 8312 16561 8340 16662
rect 8392 16584 8444 16590
rect 7932 16526 7984 16532
rect 8298 16552 8354 16561
rect 8392 16526 8444 16532
rect 8298 16487 8354 16496
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7760 16238 7880 16266
rect 7760 15706 7788 16238
rect 8022 16144 8078 16153
rect 8022 16079 8024 16088
rect 8076 16079 8078 16088
rect 8024 16050 8076 16056
rect 7838 16008 7894 16017
rect 7838 15943 7840 15952
rect 7892 15943 7894 15952
rect 7840 15914 7892 15920
rect 8036 15706 8064 16050
rect 8300 15904 8352 15910
rect 8298 15872 8300 15881
rect 8352 15872 8354 15881
rect 8298 15807 8354 15816
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7760 15502 7788 15642
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8404 12753 8432 16526
rect 8496 16182 8524 17206
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8588 15706 8616 17818
rect 8680 17066 8708 17818
rect 8772 17490 8800 19382
rect 8864 19378 8892 19926
rect 8956 19922 8984 20334
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 9048 19378 9076 20402
rect 9232 20058 9260 24647
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9324 23322 9352 23598
rect 9312 23316 9364 23322
rect 9312 23258 9364 23264
rect 9416 23118 9444 26200
rect 9692 24274 9720 26302
rect 9770 26200 9826 26302
rect 10138 26200 10194 27000
rect 10506 26200 10562 27000
rect 10874 26200 10930 27000
rect 11242 26200 11298 27000
rect 11610 26330 11666 27000
rect 11610 26302 11928 26330
rect 11610 26200 11666 26302
rect 9772 24336 9824 24342
rect 9772 24278 9824 24284
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9784 23497 9812 24278
rect 10152 23662 10180 26200
rect 10230 25800 10286 25809
rect 10230 25735 10286 25744
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 9770 23488 9826 23497
rect 9770 23423 9826 23432
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 9324 20534 9352 22986
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 22778 9444 22918
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9404 22432 9456 22438
rect 9402 22400 9404 22409
rect 9456 22400 9458 22409
rect 9402 22335 9458 22344
rect 9402 21992 9458 22001
rect 9402 21927 9404 21936
rect 9456 21927 9458 21936
rect 9404 21898 9456 21904
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9416 20641 9444 21558
rect 9402 20632 9458 20641
rect 9402 20567 9458 20576
rect 9312 20528 9364 20534
rect 9312 20470 9364 20476
rect 9508 20448 9536 23054
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 9416 20420 9536 20448
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9232 19854 9260 19994
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 8852 19372 8904 19378
rect 9036 19372 9088 19378
rect 8852 19314 8904 19320
rect 8956 19320 9036 19334
rect 8956 19314 9088 19320
rect 8956 19306 9076 19314
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 18630 8892 19110
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8956 18290 8984 19306
rect 9034 18864 9090 18873
rect 9034 18799 9090 18808
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 17746 8984 18226
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8772 17462 8892 17490
rect 8758 17368 8814 17377
rect 8758 17303 8814 17312
rect 8772 17202 8800 17303
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8772 16969 8800 17138
rect 8758 16960 8814 16969
rect 8758 16895 8814 16904
rect 8864 16590 8892 17462
rect 8956 17202 8984 17682
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9048 16946 9076 18799
rect 8956 16918 9076 16946
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8680 13161 8708 16526
rect 8956 15910 8984 16918
rect 9034 16824 9090 16833
rect 9034 16759 9036 16768
rect 9088 16759 9090 16768
rect 9036 16730 9088 16736
rect 9048 16114 9076 16730
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8666 13152 8722 13161
rect 8666 13087 8722 13096
rect 8390 12744 8446 12753
rect 7288 12708 7340 12714
rect 8390 12679 8446 12688
rect 7288 12650 7340 12656
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7010 11792 7066 11801
rect 7010 11727 7066 11736
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8772 10810 8800 15846
rect 9140 11286 9168 19654
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 9232 18358 9260 19450
rect 9324 19446 9352 19994
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9416 18834 9444 20420
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9508 18698 9536 19722
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9310 18320 9366 18329
rect 9310 18255 9366 18264
rect 9324 15706 9352 18255
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9416 13938 9444 18022
rect 9600 17610 9628 18770
rect 9692 17678 9720 22374
rect 9770 22264 9826 22273
rect 9770 22199 9826 22208
rect 9784 22166 9812 22199
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 10244 22094 10272 25735
rect 10322 24984 10378 24993
rect 10322 24919 10378 24928
rect 10152 22066 10272 22094
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9784 21729 9812 21898
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 10046 21856 10102 21865
rect 9770 21720 9826 21729
rect 9770 21655 9826 21664
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9784 18222 9812 20742
rect 9876 19174 9904 21830
rect 9968 20806 9996 21830
rect 10046 21791 10102 21800
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9876 18306 9904 18566
rect 9968 18465 9996 19654
rect 9954 18456 10010 18465
rect 9954 18391 10010 18400
rect 9876 18278 9996 18306
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9784 17270 9812 18022
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9508 16561 9536 16662
rect 9494 16552 9550 16561
rect 9494 16487 9550 16496
rect 9876 15638 9904 18158
rect 9968 16794 9996 18278
rect 10060 18204 10088 21791
rect 10152 18630 10180 22066
rect 10336 21978 10364 24919
rect 10520 23186 10548 26200
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10244 21950 10364 21978
rect 10244 18873 10272 21950
rect 10324 21616 10376 21622
rect 10324 21558 10376 21564
rect 10336 20466 10364 21558
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10520 21010 10548 21286
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10428 19938 10456 20742
rect 10520 20398 10548 20946
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10612 19990 10640 20470
rect 10600 19984 10652 19990
rect 10428 19910 10548 19938
rect 10600 19926 10652 19932
rect 10414 19816 10470 19825
rect 10414 19751 10470 19760
rect 10428 19718 10456 19751
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10230 18864 10286 18873
rect 10230 18799 10286 18808
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10060 18176 10180 18204
rect 10152 17728 10180 18176
rect 10244 18154 10272 18702
rect 10336 18290 10364 19110
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10152 17700 10272 17728
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10060 17134 10088 17546
rect 10152 17270 10180 17546
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10046 16824 10102 16833
rect 9956 16788 10008 16794
rect 10046 16759 10102 16768
rect 9956 16730 10008 16736
rect 9968 16114 9996 16730
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 10060 15502 10088 16759
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9600 13802 9628 15370
rect 10060 15162 10088 15438
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9692 14890 9720 15030
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 10244 14006 10272 17700
rect 10336 17610 10364 18226
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10336 16250 10364 16662
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10428 15162 10456 19178
rect 10520 18222 10548 19910
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 10612 16522 10640 16662
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10704 15722 10732 23802
rect 10888 23798 10916 26200
rect 11256 24274 11284 26200
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10980 21690 11008 24006
rect 11428 23656 11480 23662
rect 11428 23598 11480 23604
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11060 23248 11112 23254
rect 11060 23190 11112 23196
rect 11072 23089 11100 23190
rect 11058 23080 11114 23089
rect 11058 23015 11114 23024
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 11072 21010 11100 22034
rect 11150 21720 11206 21729
rect 11150 21655 11206 21664
rect 11164 21622 11192 21655
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11256 21486 11284 22374
rect 11348 21486 11376 23258
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11058 20904 11114 20913
rect 11058 20839 11114 20848
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10874 20224 10930 20233
rect 10796 20058 10824 20198
rect 10874 20159 10930 20168
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10782 19952 10838 19961
rect 10782 19887 10838 19896
rect 10796 15978 10824 19887
rect 10888 19825 10916 20159
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10874 19816 10930 19825
rect 10874 19751 10930 19760
rect 10980 19514 11008 19858
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10980 18902 11008 19246
rect 10968 18896 11020 18902
rect 11072 18873 11100 20839
rect 11256 20806 11284 21422
rect 11334 20904 11390 20913
rect 11334 20839 11390 20848
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11348 20505 11376 20839
rect 11334 20496 11390 20505
rect 11334 20431 11390 20440
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11164 19786 11192 19994
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11348 19258 11376 20431
rect 11256 19230 11376 19258
rect 10968 18838 11020 18844
rect 11058 18864 11114 18873
rect 11058 18799 11114 18808
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10888 18086 10916 18294
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10980 16590 11008 18158
rect 11072 17202 11100 18226
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10612 15694 10732 15722
rect 10612 15366 10640 15694
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10506 15056 10562 15065
rect 10506 14991 10508 15000
rect 10560 14991 10562 15000
rect 10508 14962 10560 14968
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10428 13870 10456 14350
rect 10520 14074 10548 14962
rect 10704 14958 10732 15370
rect 10796 15337 10824 15370
rect 10782 15328 10838 15337
rect 10782 15263 10838 15272
rect 10966 15192 11022 15201
rect 10966 15127 10968 15136
rect 11020 15127 11022 15136
rect 10968 15098 11020 15104
rect 11164 15026 11192 17002
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10704 14414 10732 14894
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 10060 9042 10088 13126
rect 10428 13025 10456 13806
rect 10704 13190 10732 14350
rect 11256 13410 11284 19230
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 17542 11376 19110
rect 11440 19009 11468 23598
rect 11520 22432 11572 22438
rect 11518 22400 11520 22409
rect 11572 22400 11574 22409
rect 11518 22335 11574 22344
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11532 20505 11560 20538
rect 11624 20534 11652 24890
rect 11900 24818 11928 26302
rect 11978 26200 12034 27000
rect 12346 26200 12402 27000
rect 12714 26200 12770 27000
rect 13082 26200 13138 27000
rect 13450 26330 13506 27000
rect 13372 26302 13506 26330
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11808 24290 11836 24346
rect 11808 24262 11928 24290
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23526 11836 24006
rect 11900 23730 11928 24262
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11992 23662 12020 26200
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11704 22704 11756 22710
rect 11704 22646 11756 22652
rect 11716 21486 11744 22646
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11716 20602 11744 21422
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11612 20528 11664 20534
rect 11518 20496 11574 20505
rect 11612 20470 11664 20476
rect 11518 20431 11574 20440
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 19514 11652 19790
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11716 19378 11744 20538
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11808 19258 11836 23462
rect 11886 21992 11942 22001
rect 11886 21927 11942 21936
rect 11900 21894 11928 21927
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11900 20534 11928 21490
rect 11992 21321 12020 23462
rect 12084 23186 12112 24754
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12268 24138 12296 24550
rect 12360 24274 12388 26200
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12176 23730 12204 24074
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 12452 23526 12480 24142
rect 12440 23520 12492 23526
rect 12728 23497 12756 26200
rect 12808 25016 12860 25022
rect 12808 24958 12860 24964
rect 12440 23462 12492 23468
rect 12714 23488 12770 23497
rect 12714 23423 12770 23432
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 12346 22944 12402 22953
rect 12346 22879 12402 22888
rect 12360 22778 12388 22879
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12164 22704 12216 22710
rect 12164 22646 12216 22652
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 12084 22166 12112 22510
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 11978 21312 12034 21321
rect 11978 21247 12034 21256
rect 12084 21010 12112 21422
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11532 19230 11836 19258
rect 11426 19000 11482 19009
rect 11426 18935 11482 18944
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 17105 11376 17478
rect 11334 17096 11390 17105
rect 11334 17031 11390 17040
rect 11532 16266 11560 19230
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18766 11744 19110
rect 11704 18760 11756 18766
rect 11756 18720 11836 18748
rect 11704 18702 11756 18708
rect 11704 18624 11756 18630
rect 11610 18592 11666 18601
rect 11704 18566 11756 18572
rect 11610 18527 11666 18536
rect 11624 16998 11652 18527
rect 11716 17746 11744 18566
rect 11808 18290 11836 18720
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17202 11744 17682
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11440 16238 11560 16266
rect 11440 15609 11468 16238
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11532 15745 11560 16050
rect 11518 15736 11574 15745
rect 11518 15671 11574 15680
rect 11426 15600 11482 15609
rect 11426 15535 11482 15544
rect 11624 15366 11652 16594
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16046 11744 16526
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11624 14482 11652 15302
rect 11716 14958 11744 15982
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11610 14104 11666 14113
rect 11610 14039 11612 14048
rect 11664 14039 11666 14048
rect 11612 14010 11664 14016
rect 11256 13382 11376 13410
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10414 13016 10470 13025
rect 11256 12986 11284 13194
rect 10414 12951 10470 12960
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11348 12646 11376 13382
rect 11808 12986 11836 18226
rect 11900 16182 11928 20198
rect 12176 19530 12204 22646
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12268 22098 12296 22510
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12728 22273 12756 22374
rect 12714 22264 12770 22273
rect 12714 22199 12770 22208
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12728 21690 12756 22102
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12440 21412 12492 21418
rect 12820 21400 12848 24958
rect 13096 24954 13124 26200
rect 13084 24948 13136 24954
rect 13084 24890 13136 24896
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 23322 13400 26302
rect 13450 26200 13506 26302
rect 13818 26330 13874 27000
rect 13818 26302 13952 26330
rect 13818 26200 13874 26302
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13556 22710 13584 24754
rect 13728 24676 13780 24682
rect 13728 24618 13780 24624
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13648 23594 13676 24278
rect 13636 23588 13688 23594
rect 13636 23530 13688 23536
rect 13634 23080 13690 23089
rect 13634 23015 13690 23024
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 12912 21894 12940 21966
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12440 21354 12492 21360
rect 12728 21372 12848 21400
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 20777 12296 21286
rect 12254 20768 12310 20777
rect 12452 20754 12480 21354
rect 12532 21344 12584 21350
rect 12728 21332 12756 21372
rect 12912 21350 12940 21830
rect 13096 21622 13124 21966
rect 13176 21956 13228 21962
rect 13176 21898 13228 21904
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 13188 21554 13216 21898
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 12532 21286 12584 21292
rect 12636 21304 12756 21332
rect 12900 21344 12952 21350
rect 12544 20942 12572 21286
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12452 20726 12572 20754
rect 12254 20703 12310 20712
rect 12438 20632 12494 20641
rect 12438 20567 12440 20576
rect 12492 20567 12494 20576
rect 12440 20538 12492 20544
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 11992 19502 12204 19530
rect 11992 16454 12020 19502
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11886 15736 11942 15745
rect 11886 15671 11942 15680
rect 11900 15638 11928 15671
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11900 14793 11928 15030
rect 11992 14958 12020 15846
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11886 14784 11942 14793
rect 11886 14719 11942 14728
rect 11992 13258 12020 14894
rect 12084 14385 12112 19110
rect 12070 14376 12126 14385
rect 12176 14362 12204 19314
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12268 17610 12296 18566
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12268 17270 12296 17546
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12360 16454 12388 18158
rect 12452 17762 12480 20266
rect 12544 19310 12572 20726
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12544 18057 12572 18362
rect 12530 18048 12586 18057
rect 12530 17983 12586 17992
rect 12636 17921 12664 21304
rect 12900 21286 12952 21292
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12622 17912 12678 17921
rect 12622 17847 12678 17856
rect 12728 17762 12756 20878
rect 12820 19972 12848 20946
rect 12912 20806 12940 20946
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20602 13216 20742
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12900 19984 12952 19990
rect 12820 19944 12900 19972
rect 12900 19926 12952 19932
rect 13372 19122 13400 22578
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13556 22234 13584 22374
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13464 20398 13492 21422
rect 13556 21146 13584 22170
rect 13648 22030 13676 23015
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13740 21690 13768 24618
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13832 23662 13860 24074
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13924 23186 13952 26302
rect 14186 26200 14242 27000
rect 14554 26200 14610 27000
rect 14922 26200 14978 27000
rect 15290 26200 15346 27000
rect 15658 26200 15714 27000
rect 16026 26330 16082 27000
rect 15856 26302 16082 26330
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14108 24410 14136 24550
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13912 22160 13964 22166
rect 13912 22102 13964 22108
rect 13818 21992 13874 22001
rect 13818 21927 13874 21936
rect 13832 21894 13860 21927
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13924 21690 13952 22102
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13912 21412 13964 21418
rect 13912 21354 13964 21360
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13648 21049 13676 21082
rect 13634 21040 13690 21049
rect 13634 20975 13690 20984
rect 13924 20602 13952 21354
rect 14016 20942 14044 24210
rect 14094 23352 14150 23361
rect 14200 23322 14228 26200
rect 14568 24274 14596 26200
rect 14936 25022 14964 26200
rect 14924 25016 14976 25022
rect 14924 24958 14976 24964
rect 15016 24676 15068 24682
rect 15016 24618 15068 24624
rect 14556 24268 14608 24274
rect 14556 24210 14608 24216
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14832 24064 14884 24070
rect 14832 24006 14884 24012
rect 14752 23798 14780 24006
rect 14740 23792 14792 23798
rect 14740 23734 14792 23740
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14094 23287 14150 23296
rect 14188 23316 14240 23322
rect 14108 22817 14136 23287
rect 14188 23258 14240 23264
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14094 22808 14150 22817
rect 14094 22743 14150 22752
rect 14200 22710 14228 23054
rect 14554 22808 14610 22817
rect 14554 22743 14610 22752
rect 14188 22704 14240 22710
rect 14188 22646 14240 22652
rect 14200 22030 14228 22646
rect 14568 22574 14596 22743
rect 14660 22574 14688 23190
rect 14752 22778 14780 23598
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14554 22400 14610 22409
rect 14554 22335 14610 22344
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14004 20936 14056 20942
rect 14004 20878 14056 20884
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 19310 13492 20334
rect 13556 20233 13584 20402
rect 13542 20224 13598 20233
rect 13542 20159 13598 20168
rect 13818 20224 13874 20233
rect 13818 20159 13874 20168
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13544 19848 13596 19854
rect 13740 19836 13768 19926
rect 13596 19808 13768 19836
rect 13544 19790 13596 19796
rect 13542 19680 13598 19689
rect 13542 19615 13598 19624
rect 13726 19680 13782 19689
rect 13726 19615 13782 19624
rect 13556 19417 13584 19615
rect 13542 19408 13598 19417
rect 13542 19343 13598 19352
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13740 19174 13768 19615
rect 13832 19514 13860 20159
rect 13924 19854 13952 20538
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13728 19168 13780 19174
rect 13372 19094 13676 19122
rect 13728 19110 13780 19116
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13358 19000 13414 19009
rect 13358 18935 13414 18944
rect 13372 18426 13400 18935
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13084 18216 13136 18222
rect 12820 18164 13084 18170
rect 12820 18158 13136 18164
rect 12820 18142 13124 18158
rect 12820 18086 12848 18142
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13464 17814 13492 18566
rect 13452 17808 13504 17814
rect 12452 17746 12664 17762
rect 12452 17740 12676 17746
rect 12452 17734 12624 17740
rect 12728 17734 12848 17762
rect 13452 17750 13504 17756
rect 12624 17682 12676 17688
rect 12440 17536 12492 17542
rect 12438 17504 12440 17513
rect 12532 17536 12584 17542
rect 12492 17504 12494 17513
rect 12532 17478 12584 17484
rect 12438 17439 12494 17448
rect 12452 17134 12480 17439
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12544 16522 12572 17478
rect 12636 17134 12664 17682
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12728 16658 12756 17546
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 16522 12756 16594
rect 12532 16516 12584 16522
rect 12532 16458 12584 16464
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 16046 12388 16390
rect 12728 16182 12756 16458
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12348 15904 12400 15910
rect 12346 15872 12348 15881
rect 12400 15872 12402 15881
rect 12346 15807 12402 15816
rect 12728 15434 12756 16118
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 12360 14414 12388 15370
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12636 14793 12664 15098
rect 12728 15094 12756 15370
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12622 14784 12678 14793
rect 12622 14719 12678 14728
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12348 14408 12400 14414
rect 12176 14346 12296 14362
rect 12348 14350 12400 14356
rect 12176 14340 12308 14346
rect 12176 14334 12256 14340
rect 12070 14311 12126 14320
rect 12256 14282 12308 14288
rect 12360 13938 12388 14350
rect 12452 13938 12480 14554
rect 12636 14482 12664 14719
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12728 14074 12756 14350
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12346 13288 12402 13297
rect 11980 13252 12032 13258
rect 12728 13258 12756 13738
rect 12346 13223 12402 13232
rect 12716 13252 12768 13258
rect 11980 13194 12032 13200
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 12360 12850 12388 13223
rect 12716 13194 12768 13200
rect 12728 12986 12756 13194
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12728 10577 12756 11766
rect 12820 11558 12848 17734
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15337 13400 15846
rect 13358 15328 13414 15337
rect 13358 15263 13414 15272
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14074 13400 14962
rect 13464 14414 13492 17206
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13556 14482 13584 16050
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13372 13462 13400 13670
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 11830 13400 13126
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12714 10568 12770 10577
rect 13648 10538 13676 19094
rect 13832 18766 13860 19450
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13832 18426 13860 18702
rect 13924 18698 13952 19654
rect 13912 18692 13964 18698
rect 13912 18634 13964 18640
rect 13820 18420 13872 18426
rect 14016 18408 14044 20742
rect 14108 20534 14136 21830
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14200 20233 14228 21966
rect 14370 21176 14426 21185
rect 14370 21111 14426 21120
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14186 20224 14242 20233
rect 14186 20159 14242 20168
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14108 19378 14136 19926
rect 14292 19530 14320 20878
rect 14200 19502 14320 19530
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14108 18970 14136 19178
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 13820 18362 13872 18368
rect 13924 18380 14044 18408
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16658 13768 16934
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13740 15162 13768 16118
rect 13832 15502 13860 16390
rect 13924 15502 13952 18380
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14016 17882 14044 18226
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13832 14822 13860 15098
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13910 14784 13966 14793
rect 13910 14719 13966 14728
rect 13818 14648 13874 14657
rect 13740 14606 13818 14634
rect 13740 14278 13768 14606
rect 13818 14583 13874 14592
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13832 14278 13860 14486
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13726 13832 13782 13841
rect 13726 13767 13728 13776
rect 13780 13767 13782 13776
rect 13728 13738 13780 13744
rect 13820 13728 13872 13734
rect 13924 13682 13952 14719
rect 13872 13676 13952 13682
rect 13820 13670 13952 13676
rect 13832 13654 13952 13670
rect 13924 13530 13952 13654
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 12714 10503 12770 10512
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 13832 8906 13860 11630
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 9324 6458 9352 8842
rect 14016 8566 14044 17478
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14108 15910 14136 17070
rect 14200 16289 14228 19502
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14292 18970 14320 19382
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16522 14320 16934
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 14186 16280 14242 16289
rect 14186 16215 14242 16224
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 15688 14228 15846
rect 14292 15745 14320 16458
rect 14108 15660 14228 15688
rect 14278 15736 14334 15745
rect 14278 15671 14334 15680
rect 14108 15366 14136 15660
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 15026 14136 15302
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14200 13258 14228 15506
rect 14292 14482 14320 15506
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 14006 14320 14418
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14292 13394 14320 13942
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14292 12986 14320 13330
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14292 12434 14320 12922
rect 14384 12850 14412 21111
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 14476 19786 14504 19926
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14476 19514 14504 19722
rect 14568 19514 14596 22335
rect 14752 22234 14780 22714
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 20602 14780 21286
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14660 19334 14688 19790
rect 14752 19378 14780 20538
rect 14568 19306 14688 19334
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14476 18426 14504 18770
rect 14568 18698 14596 19306
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14646 19136 14702 19145
rect 14646 19071 14702 19080
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14554 18320 14610 18329
rect 14554 18255 14610 18264
rect 14462 17912 14518 17921
rect 14462 17847 14518 17856
rect 14476 17678 14504 17847
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14568 17490 14596 18255
rect 14476 17462 14596 17490
rect 14476 15473 14504 17462
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14462 15464 14518 15473
rect 14462 15399 14518 15408
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14476 14346 14504 14826
rect 14568 14482 14596 15982
rect 14660 15910 14688 19071
rect 14752 18902 14780 19178
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14752 16998 14780 18838
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14646 15736 14702 15745
rect 14646 15671 14702 15680
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14476 13841 14504 13942
rect 14568 13870 14596 14418
rect 14556 13864 14608 13870
rect 14462 13832 14518 13841
rect 14556 13806 14608 13812
rect 14462 13767 14518 13776
rect 14476 13376 14504 13767
rect 14556 13388 14608 13394
rect 14476 13348 14556 13376
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14476 12442 14504 13348
rect 14556 13330 14608 13336
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14108 12406 14320 12434
rect 14464 12436 14516 12442
rect 14108 11898 14136 12406
rect 14464 12378 14516 12384
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14384 10606 14412 12174
rect 14476 11830 14504 12378
rect 14568 11898 14596 13194
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14660 9674 14688 15671
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 11014 14780 14894
rect 14844 11354 14872 24006
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 14936 23322 14964 23462
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 14936 22710 14964 23258
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14922 22536 14978 22545
rect 14922 22471 14924 22480
rect 14976 22471 14978 22480
rect 14924 22442 14976 22448
rect 15028 22409 15056 24618
rect 15198 24440 15254 24449
rect 15198 24375 15254 24384
rect 15212 24177 15240 24375
rect 15198 24168 15254 24177
rect 15198 24103 15254 24112
rect 15014 22400 15070 22409
rect 15014 22335 15070 22344
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 14936 21350 14964 22170
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 15014 21040 15070 21049
rect 15014 20975 15070 20984
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14936 19242 14964 19722
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14936 17746 14964 18702
rect 15028 18601 15056 20975
rect 15120 19378 15148 21490
rect 15212 21146 15240 21490
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15212 20874 15240 21082
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 15212 20534 15240 20810
rect 15200 20528 15252 20534
rect 15304 20505 15332 26200
rect 15476 25016 15528 25022
rect 15476 24958 15528 24964
rect 15488 24342 15516 24958
rect 15566 24576 15622 24585
rect 15566 24511 15622 24520
rect 15580 24342 15608 24511
rect 15476 24336 15528 24342
rect 15476 24278 15528 24284
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15580 23798 15608 24006
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15396 22982 15424 23462
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15476 22976 15528 22982
rect 15672 22953 15700 26200
rect 15476 22918 15528 22924
rect 15658 22944 15714 22953
rect 15200 20470 15252 20476
rect 15290 20496 15346 20505
rect 15212 19854 15240 20470
rect 15290 20431 15346 20440
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15212 18816 15240 19790
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 19553 15332 19654
rect 15290 19544 15346 19553
rect 15290 19479 15346 19488
rect 15120 18788 15240 18816
rect 15120 18630 15148 18788
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15108 18624 15160 18630
rect 15014 18592 15070 18601
rect 15108 18566 15160 18572
rect 15014 18527 15070 18536
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14936 16658 14964 17682
rect 15120 17610 15148 18566
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15014 17232 15070 17241
rect 15014 17167 15070 17176
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 15028 16522 15056 17167
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16794 15148 16934
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 15434 15056 16458
rect 15212 16114 15240 18634
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15304 15910 15332 17138
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 14346 15056 15370
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15120 14482 15148 14758
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 12434 14964 14214
rect 15028 13938 15056 14282
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15028 13394 15056 13874
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15028 13258 15056 13330
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14936 12406 15056 12434
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 15028 10198 15056 12406
rect 15120 11898 15148 13330
rect 15198 12336 15254 12345
rect 15198 12271 15254 12280
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15212 11150 15240 12271
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 14476 9646 14688 9674
rect 14476 9178 14504 9646
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 15396 8090 15424 22918
rect 15488 21457 15516 22918
rect 15658 22879 15714 22888
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15474 21448 15530 21457
rect 15474 21383 15530 21392
rect 15476 20596 15528 20602
rect 15580 20584 15608 21490
rect 15672 21486 15700 22646
rect 15856 22094 15884 26302
rect 16026 26200 16082 26302
rect 16394 26200 16450 27000
rect 16762 26330 16818 27000
rect 16592 26302 16818 26330
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 16224 24274 16252 24890
rect 16408 24449 16436 26200
rect 16394 24440 16450 24449
rect 16394 24375 16450 24384
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 15934 23216 15990 23225
rect 15934 23151 15990 23160
rect 15764 22066 15884 22094
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15528 20556 15608 20584
rect 15476 20538 15528 20544
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15488 19514 15516 19722
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15488 18222 15516 18362
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15580 17746 15608 18906
rect 15672 18698 15700 19110
rect 15660 18692 15712 18698
rect 15660 18634 15712 18640
rect 15672 18290 15700 18634
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15488 17134 15516 17546
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15580 15638 15608 17682
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15672 17241 15700 17546
rect 15658 17232 15714 17241
rect 15658 17167 15714 17176
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15672 13161 15700 16662
rect 15764 16658 15792 22066
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15856 21554 15884 21898
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15844 20800 15896 20806
rect 15842 20768 15844 20777
rect 15896 20768 15898 20777
rect 15842 20703 15898 20712
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15856 16425 15884 18294
rect 15948 17746 15976 23151
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 16040 20806 16068 21354
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 20058 16068 20198
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18698 16068 19246
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15842 16416 15898 16425
rect 15842 16351 15898 16360
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15750 15872 15806 15881
rect 15750 15807 15806 15816
rect 15658 13152 15714 13161
rect 15658 13087 15714 13096
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15672 10266 15700 12174
rect 15764 11150 15792 15807
rect 15856 12900 15884 16050
rect 15948 13530 15976 17274
rect 16040 16794 16068 18634
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16040 15162 16068 15302
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13530 16068 13670
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15856 12872 16068 12900
rect 15842 11928 15898 11937
rect 15842 11863 15898 11872
rect 15856 11830 15884 11863
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15764 10810 15792 11086
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 16040 9382 16068 12872
rect 16132 11354 16160 23734
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16210 22944 16266 22953
rect 16210 22879 16266 22888
rect 16224 22234 16252 22879
rect 16316 22778 16344 23258
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16316 21554 16344 22714
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16302 21448 16358 21457
rect 16302 21383 16304 21392
rect 16356 21383 16358 21392
rect 16304 21354 16356 21360
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16224 21146 16252 21286
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16224 20788 16252 20946
rect 16316 20942 16344 21354
rect 16408 21332 16436 23462
rect 16500 22710 16528 24142
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16500 21486 16528 22442
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16408 21304 16528 21332
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16224 20760 16344 20788
rect 16210 20360 16266 20369
rect 16210 20295 16266 20304
rect 16224 20262 16252 20295
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16224 18698 16252 19450
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16224 18290 16252 18634
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16224 17241 16252 18226
rect 16210 17232 16266 17241
rect 16210 17167 16266 17176
rect 16224 15910 16252 17167
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16210 15600 16266 15609
rect 16210 15535 16266 15544
rect 16224 13025 16252 15535
rect 16316 13394 16344 20760
rect 16408 19990 16436 20946
rect 16500 20777 16528 21304
rect 16486 20768 16542 20777
rect 16486 20703 16542 20712
rect 16396 19984 16448 19990
rect 16396 19926 16448 19932
rect 16486 18456 16542 18465
rect 16486 18391 16542 18400
rect 16500 15978 16528 18391
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15638 16436 15846
rect 16592 15638 16620 26302
rect 16762 26200 16818 26302
rect 17130 26200 17186 27000
rect 17498 26200 17554 27000
rect 17866 26200 17922 27000
rect 18234 26330 18290 27000
rect 18234 26302 18552 26330
rect 18234 26200 18290 26302
rect 16946 24440 17002 24449
rect 16856 24404 16908 24410
rect 16946 24375 16948 24384
rect 16856 24346 16908 24352
rect 17000 24375 17002 24384
rect 16948 24346 17000 24352
rect 16764 23248 16816 23254
rect 16764 23190 16816 23196
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16684 22778 16712 23054
rect 16776 22982 16804 23190
rect 16868 23118 16896 24346
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16776 22817 16804 22918
rect 16762 22808 16818 22817
rect 16672 22772 16724 22778
rect 16762 22743 16818 22752
rect 16672 22714 16724 22720
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16856 22636 16908 22642
rect 16960 22624 16988 23258
rect 16908 22596 16988 22624
rect 16856 22578 16908 22584
rect 16776 22545 16804 22578
rect 16762 22536 16818 22545
rect 16762 22471 16818 22480
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16868 22094 16896 22442
rect 16868 22066 16988 22094
rect 16762 21992 16818 22001
rect 16762 21927 16764 21936
rect 16816 21927 16818 21936
rect 16764 21898 16816 21904
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16684 21146 16712 21626
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16776 20874 16804 21354
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16670 20224 16726 20233
rect 16776 20210 16804 20470
rect 16868 20233 16896 21830
rect 16726 20182 16804 20210
rect 16670 20159 16726 20168
rect 16776 20074 16804 20182
rect 16854 20224 16910 20233
rect 16854 20159 16910 20168
rect 16776 20046 16896 20074
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16684 19718 16712 19926
rect 16764 19848 16816 19854
rect 16762 19816 16764 19825
rect 16816 19816 16818 19825
rect 16762 19751 16818 19760
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16776 19514 16804 19654
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16868 19378 16896 20046
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16776 18873 16804 18906
rect 16762 18864 16818 18873
rect 16960 18834 16988 22066
rect 17052 21554 17080 23666
rect 17144 23050 17172 26200
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 17236 22930 17264 24550
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17328 23089 17356 24006
rect 17512 23497 17540 26200
rect 17880 24721 17908 26200
rect 18236 24948 18288 24954
rect 18236 24890 18288 24896
rect 17866 24712 17922 24721
rect 17866 24647 17922 24656
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17604 23662 17632 24550
rect 18248 24342 18276 24890
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18236 24336 18288 24342
rect 18236 24278 18288 24284
rect 17960 24268 18012 24274
rect 17960 24210 18012 24216
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 17972 24177 18000 24210
rect 17958 24168 18014 24177
rect 17958 24103 18014 24112
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23662 18368 24210
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17868 23520 17920 23526
rect 17498 23488 17554 23497
rect 17920 23480 18000 23508
rect 17868 23462 17920 23468
rect 17498 23423 17554 23432
rect 17972 23186 18000 23480
rect 18064 23322 18092 23598
rect 18142 23488 18198 23497
rect 18142 23423 18198 23432
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17314 23080 17370 23089
rect 17314 23015 17370 23024
rect 17408 22976 17460 22982
rect 17236 22902 17356 22930
rect 17684 22976 17736 22982
rect 17408 22918 17460 22924
rect 17682 22944 17684 22953
rect 17736 22944 17738 22953
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 17144 22098 17172 22374
rect 17236 22234 17264 22646
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17132 22092 17184 22098
rect 17328 22094 17356 22902
rect 17132 22034 17184 22040
rect 17236 22066 17356 22094
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 17144 21418 17172 21898
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 19514 17080 21286
rect 17236 21146 17264 22066
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16762 18799 16818 18808
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16592 15026 16620 15574
rect 16684 15434 16712 17682
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16500 14414 16528 14826
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16210 13016 16266 13025
rect 16210 12951 16266 12960
rect 16316 12170 16344 13126
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16302 10704 16358 10713
rect 16302 10639 16304 10648
rect 16356 10639 16358 10648
rect 16304 10610 16356 10616
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 16408 7954 16436 13806
rect 16500 13394 16528 14350
rect 16684 14278 16712 15370
rect 16776 15094 16804 18226
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16868 15706 16896 16934
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16776 14521 16804 14894
rect 16762 14512 16818 14521
rect 16762 14447 16818 14456
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16670 13560 16726 13569
rect 16670 13495 16726 13504
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16684 13297 16712 13495
rect 16670 13288 16726 13297
rect 16776 13258 16804 13670
rect 16670 13223 16726 13232
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16762 12880 16818 12889
rect 16868 12850 16896 15506
rect 16762 12815 16764 12824
rect 16816 12815 16818 12824
rect 16856 12844 16908 12850
rect 16764 12786 16816 12792
rect 16856 12786 16908 12792
rect 16670 12472 16726 12481
rect 16868 12434 16896 12786
rect 16670 12407 16726 12416
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11898 16528 12106
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 9674 16528 11834
rect 16684 11150 16712 12407
rect 16776 12406 16896 12434
rect 16776 12306 16804 12406
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16960 11354 16988 17138
rect 17052 12306 17080 17546
rect 17144 16833 17172 20878
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17236 18902 17264 20334
rect 17328 19310 17356 21422
rect 17420 20942 17448 22918
rect 17682 22879 17738 22888
rect 17788 22574 17816 23122
rect 18064 23118 18092 23258
rect 18156 23225 18184 23423
rect 18340 23322 18368 23598
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18142 23216 18198 23225
rect 18142 23151 18198 23160
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18328 23044 18380 23050
rect 18328 22986 18380 22992
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 21593 17540 21966
rect 17604 21729 17632 22374
rect 18340 22273 18368 22986
rect 18432 22982 18460 24822
rect 18524 24698 18552 26302
rect 18602 26200 18658 27000
rect 18696 26376 18748 26382
rect 18970 26330 19026 27000
rect 18748 26324 19026 26330
rect 18696 26318 19026 26324
rect 18708 26302 19026 26318
rect 18970 26200 19026 26302
rect 19338 26200 19394 27000
rect 19706 26200 19762 27000
rect 20074 26200 20130 27000
rect 20442 26200 20498 27000
rect 20810 26200 20866 27000
rect 21178 26200 21234 27000
rect 21546 26330 21602 27000
rect 21284 26302 21602 26330
rect 21284 26217 21312 26302
rect 21270 26208 21326 26217
rect 18616 24818 18644 26200
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18524 24670 19104 24698
rect 18878 24576 18934 24585
rect 18878 24511 18934 24520
rect 18512 24200 18564 24206
rect 18564 24160 18644 24188
rect 18512 24142 18564 24148
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18420 22976 18472 22982
rect 18420 22918 18472 22924
rect 18326 22264 18382 22273
rect 18326 22199 18382 22208
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17776 21888 17828 21894
rect 18156 21876 18184 22034
rect 18236 21888 18288 21894
rect 18156 21848 18236 21876
rect 17776 21830 17828 21836
rect 18236 21830 18288 21836
rect 17590 21720 17646 21729
rect 17590 21655 17646 21664
rect 17696 21622 17724 21830
rect 17684 21616 17736 21622
rect 17498 21584 17554 21593
rect 17684 21558 17736 21564
rect 17498 21519 17500 21528
rect 17552 21519 17554 21528
rect 17500 21490 17552 21496
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17406 20632 17462 20641
rect 17406 20567 17462 20576
rect 17420 19961 17448 20567
rect 17406 19952 17462 19961
rect 17512 19922 17540 21286
rect 17684 20868 17736 20874
rect 17684 20810 17736 20816
rect 17406 19887 17462 19896
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17406 19408 17462 19417
rect 17512 19394 17540 19858
rect 17462 19366 17540 19394
rect 17406 19343 17462 19352
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17236 17377 17264 18634
rect 17328 17542 17356 19246
rect 17512 18290 17540 19366
rect 17604 18902 17632 19858
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17420 17678 17448 18158
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17222 17368 17278 17377
rect 17222 17303 17278 17312
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17130 16824 17186 16833
rect 17130 16759 17186 16768
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17144 14958 17172 16526
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 15570 17264 16390
rect 17328 15706 17356 16458
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17224 15088 17276 15094
rect 17328 15076 17356 15370
rect 17276 15048 17356 15076
rect 17224 15030 17276 15036
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17222 14920 17278 14929
rect 17222 14855 17278 14864
rect 17236 14464 17264 14855
rect 17144 14436 17264 14464
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16684 10810 16712 11086
rect 17052 11082 17080 12038
rect 17144 11150 17172 14436
rect 17224 14340 17276 14346
rect 17328 14328 17356 15048
rect 17276 14300 17356 14328
rect 17224 14282 17276 14288
rect 17236 13938 17264 14282
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17236 13258 17264 13874
rect 17420 13734 17448 17070
rect 17512 14074 17540 18022
rect 17604 17882 17632 18838
rect 17696 18057 17724 20810
rect 17788 19417 17816 21830
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18524 21690 18552 23462
rect 18616 22794 18644 24160
rect 18696 24064 18748 24070
rect 18696 24006 18748 24012
rect 18708 23662 18736 24006
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18696 23248 18748 23254
rect 18696 23190 18748 23196
rect 18708 22982 18736 23190
rect 18800 23050 18828 23462
rect 18788 23044 18840 23050
rect 18788 22986 18840 22992
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18616 22766 18736 22794
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18616 22234 18644 22646
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 17868 21412 17920 21418
rect 17868 21354 17920 21360
rect 17774 19408 17830 19417
rect 17774 19343 17830 19352
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17682 18048 17738 18057
rect 17682 17983 17738 17992
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 17338 17632 17614
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17696 17270 17724 17546
rect 17788 17542 17816 18566
rect 17880 18272 17908 21354
rect 18340 21078 18368 21422
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18328 21072 18380 21078
rect 18328 21014 18380 21020
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17960 20596 18012 20602
rect 18432 20584 18460 21082
rect 17960 20538 18012 20544
rect 18156 20556 18460 20584
rect 17972 19718 18000 20538
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 18064 19718 18092 19926
rect 18156 19922 18184 20556
rect 18616 20534 18644 22170
rect 18708 21185 18736 22766
rect 18694 21176 18750 21185
rect 18694 21111 18750 21120
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18708 20602 18736 20946
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18604 20528 18656 20534
rect 18340 20476 18604 20482
rect 18340 20470 18656 20476
rect 18340 20466 18644 20470
rect 18328 20460 18644 20466
rect 18380 20454 18644 20460
rect 18328 20402 18380 20408
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18248 19718 18276 20198
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18340 19446 18368 20402
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17960 18284 18012 18290
rect 17880 18244 17960 18272
rect 17960 18226 18012 18232
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 17338 17816 17478
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17880 17202 17908 17818
rect 18248 17542 18276 18090
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 17202 18368 19110
rect 18604 18828 18656 18834
rect 18432 18788 18604 18816
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17590 15464 17646 15473
rect 17696 15434 17724 16458
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17590 15399 17646 15408
rect 17684 15428 17736 15434
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17604 13954 17632 15399
rect 17684 15370 17736 15376
rect 17696 14958 17724 15370
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14482 18368 14758
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18052 14340 18104 14346
rect 17880 14300 18052 14328
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 14006 17816 14214
rect 17880 14056 17908 14300
rect 18052 14282 18104 14288
rect 18432 14260 18460 18788
rect 18604 18770 18656 18776
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18524 14550 18552 18090
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17270 18644 17546
rect 18604 17264 18656 17270
rect 18708 17241 18736 19858
rect 18604 17206 18656 17212
rect 18694 17232 18750 17241
rect 18616 15434 18644 17206
rect 18694 17167 18750 17176
rect 18800 16561 18828 19926
rect 18892 18358 18920 24511
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 18984 22234 19012 23122
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18984 21554 19012 21830
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18984 21146 19012 21490
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18786 16552 18842 16561
rect 18786 16487 18842 16496
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18616 14958 18644 15370
rect 18708 15162 18736 15642
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18708 14618 18736 14758
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 18340 14232 18460 14260
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17880 14028 18092 14056
rect 17512 13926 17632 13954
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 12918 17264 13194
rect 17224 12912 17276 12918
rect 17276 12872 17356 12900
rect 17224 12854 17276 12860
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 17052 10674 17080 11018
rect 17144 10810 17172 11086
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16500 9646 16620 9674
rect 16592 9586 16620 9646
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 17236 6662 17264 12242
rect 17328 11830 17356 12872
rect 17512 12866 17540 13926
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17604 13190 17632 13738
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17512 12838 17632 12866
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12442 17540 12718
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17406 11384 17462 11393
rect 17406 11319 17408 11328
rect 17460 11319 17462 11328
rect 17408 11290 17460 11296
rect 17604 10810 17632 12838
rect 17696 12730 17724 13942
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17788 12986 17816 13398
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17696 12702 17816 12730
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17788 9586 17816 12702
rect 17880 11218 17908 13874
rect 18064 13326 18092 14028
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12782 18368 14232
rect 18524 13394 18552 14486
rect 18616 14278 18644 14486
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18602 13696 18658 13705
rect 18602 13631 18658 13640
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18616 12832 18644 13631
rect 18432 12804 18644 12832
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18432 12434 18460 12804
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18340 12406 18460 12434
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17866 11112 17922 11121
rect 17866 11047 17922 11056
rect 17960 11076 18012 11082
rect 17880 10810 17908 11047
rect 18144 11076 18196 11082
rect 18012 11036 18144 11064
rect 17960 11018 18012 11024
rect 18144 11018 18196 11024
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18248 10062 18276 10678
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18340 9994 18368 12406
rect 18524 11880 18552 12650
rect 18432 11852 18552 11880
rect 18432 10130 18460 11852
rect 18616 11694 18644 12650
rect 18694 12200 18750 12209
rect 18694 12135 18696 12144
rect 18748 12135 18750 12144
rect 18696 12106 18748 12112
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18524 11286 18552 11562
rect 18512 11280 18564 11286
rect 18708 11257 18736 12106
rect 18800 11354 18828 16118
rect 18892 16046 18920 17478
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18892 15162 18920 15982
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18892 14006 18920 15098
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12986 18920 13126
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18984 12900 19012 19654
rect 19076 19145 19104 24670
rect 19246 23488 19302 23497
rect 19352 23474 19380 26200
rect 19430 25392 19486 25401
rect 19430 25327 19486 25336
rect 19302 23446 19380 23474
rect 19246 23423 19302 23432
rect 19248 23180 19300 23186
rect 19300 23140 19380 23168
rect 19248 23122 19300 23128
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 19168 21962 19196 22918
rect 19352 22030 19380 23140
rect 19444 22642 19472 25327
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19430 22536 19486 22545
rect 19430 22471 19486 22480
rect 19444 22438 19472 22471
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 19352 21350 19380 21966
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20942 19380 21286
rect 19536 21146 19564 24006
rect 19614 23488 19670 23497
rect 19614 23423 19670 23432
rect 19628 22778 19656 23423
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19616 22568 19668 22574
rect 19616 22510 19668 22516
rect 19628 21962 19656 22510
rect 19720 22506 19748 26200
rect 20088 25022 20116 26200
rect 20456 26081 20484 26200
rect 20442 26072 20498 26081
rect 20442 26007 20498 26016
rect 20626 25664 20682 25673
rect 20626 25599 20682 25608
rect 20076 25016 20128 25022
rect 20076 24958 20128 24964
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 19800 23520 19852 23526
rect 19904 23497 19932 24346
rect 20548 24206 20576 24686
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 20180 23497 20208 24142
rect 20260 23792 20312 23798
rect 20640 23769 20668 25599
rect 20260 23734 20312 23740
rect 20626 23760 20682 23769
rect 19800 23462 19852 23468
rect 19890 23488 19946 23497
rect 19708 22500 19760 22506
rect 19708 22442 19760 22448
rect 19812 22166 19840 23462
rect 19890 23423 19946 23432
rect 20166 23488 20222 23497
rect 20166 23423 20222 23432
rect 20272 23050 20300 23734
rect 20626 23695 20628 23704
rect 20680 23695 20682 23704
rect 20628 23666 20680 23672
rect 20824 23361 20852 26200
rect 21192 25809 21220 26200
rect 21546 26200 21602 26302
rect 21914 26200 21970 27000
rect 22190 26344 22246 26353
rect 22190 26279 22246 26288
rect 21270 26143 21326 26152
rect 21928 25945 21956 26200
rect 22204 26058 22232 26279
rect 22282 26200 22338 27000
rect 22650 26330 22706 27000
rect 23018 26330 23074 27000
rect 23386 26330 23442 27000
rect 22388 26302 22706 26330
rect 22296 26058 22324 26200
rect 22204 26030 22324 26058
rect 21914 25936 21970 25945
rect 21914 25871 21970 25880
rect 21178 25800 21234 25809
rect 21178 25735 21234 25744
rect 22098 24712 22154 24721
rect 21456 24676 21508 24682
rect 22098 24647 22154 24656
rect 21456 24618 21508 24624
rect 21270 24304 21326 24313
rect 21270 24239 21326 24248
rect 21284 24070 21312 24239
rect 21468 24206 21496 24618
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 20810 23352 20866 23361
rect 20810 23287 20866 23296
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20272 22778 20300 22986
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 19800 22160 19852 22166
rect 19800 22102 19852 22108
rect 19616 21956 19668 21962
rect 19616 21898 19668 21904
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20618 19380 20878
rect 19260 20590 19380 20618
rect 19260 20398 19288 20590
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19522 20360 19578 20369
rect 19260 19174 19288 20334
rect 19522 20295 19578 20304
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19825 19380 19858
rect 19536 19825 19564 20295
rect 19338 19816 19394 19825
rect 19338 19751 19394 19760
rect 19522 19816 19578 19825
rect 19522 19751 19578 19760
rect 19352 19718 19380 19751
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19536 19417 19564 19450
rect 19522 19408 19578 19417
rect 19522 19343 19578 19352
rect 19248 19168 19300 19174
rect 19062 19136 19118 19145
rect 19248 19110 19300 19116
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19062 19071 19118 19080
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19076 13190 19104 18838
rect 19168 18698 19196 18838
rect 19260 18766 19288 19110
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19156 18692 19208 18698
rect 19156 18634 19208 18640
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16454 19196 17070
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19168 12918 19196 15846
rect 19260 14278 19288 18022
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19352 16658 19380 17274
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 15094 19380 16458
rect 19444 15366 19472 19110
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19536 16969 19564 18634
rect 19628 17252 19656 21898
rect 19720 21729 19748 21898
rect 19706 21720 19762 21729
rect 19706 21655 19762 21664
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19996 20641 20024 20810
rect 19982 20632 20038 20641
rect 19982 20567 20038 20576
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19996 20398 20024 20470
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19904 19446 19932 20334
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20088 19446 20116 19790
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19904 19310 19932 19382
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19996 19174 20024 19314
rect 20168 19236 20220 19242
rect 20168 19178 20220 19184
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19800 18828 19852 18834
rect 19720 18788 19800 18816
rect 19720 18329 19748 18788
rect 19800 18770 19852 18776
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19706 18320 19762 18329
rect 19996 18290 20024 18566
rect 19706 18255 19762 18264
rect 19984 18284 20036 18290
rect 19720 18222 19748 18255
rect 19984 18226 20036 18232
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17320 19748 17478
rect 19720 17292 19840 17320
rect 19628 17224 19748 17252
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19522 16960 19578 16969
rect 19522 16895 19578 16904
rect 19524 16788 19576 16794
rect 19628 16776 19656 17070
rect 19576 16748 19656 16776
rect 19524 16730 19576 16736
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19352 14074 19380 14894
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19444 14346 19472 14554
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19156 12912 19208 12918
rect 18984 12872 19104 12900
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 19076 12730 19104 12872
rect 19156 12854 19208 12860
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18512 11222 18564 11228
rect 18694 11248 18750 11257
rect 18694 11183 18750 11192
rect 18602 11112 18658 11121
rect 18602 11047 18658 11056
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18616 9994 18644 11047
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17604 9489 17632 9522
rect 17590 9480 17646 9489
rect 17590 9415 17646 9424
rect 17604 9178 17632 9415
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 8680 4826 8708 6258
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18340 5302 18368 8910
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6748 2854 6776 2994
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 6748 800 6776 2790
rect 7024 2650 7052 4558
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7208 2446 7236 3334
rect 7484 3194 7512 3470
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 18892 3058 18920 12106
rect 18984 7886 19012 12718
rect 19076 12702 19196 12730
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19076 7818 19104 12582
rect 19168 11744 19196 12702
rect 19260 12345 19288 13806
rect 19246 12336 19302 12345
rect 19246 12271 19302 12280
rect 19352 12238 19380 14010
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19352 11898 19380 12174
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11762 19472 12582
rect 19432 11756 19484 11762
rect 19168 11716 19288 11744
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19168 11286 19196 11562
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19168 9994 19196 10610
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19168 8430 19196 9522
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 19260 7546 19288 11716
rect 19432 11698 19484 11704
rect 19430 11656 19486 11665
rect 19430 11591 19486 11600
rect 19444 11354 19472 11591
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19430 11248 19486 11257
rect 19340 11212 19392 11218
rect 19430 11183 19486 11192
rect 19340 11154 19392 11160
rect 19352 10849 19380 11154
rect 19338 10840 19394 10849
rect 19444 10810 19472 11183
rect 19338 10775 19394 10784
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19352 7886 19380 9862
rect 19444 9722 19472 9862
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19430 9208 19486 9217
rect 19430 9143 19432 9152
rect 19484 9143 19486 9152
rect 19432 9114 19484 9120
rect 19536 8498 19564 15302
rect 19628 14618 19656 16050
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19628 13530 19656 13670
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19628 11064 19656 12854
rect 19720 12753 19748 17224
rect 19812 12986 19840 17292
rect 19904 15706 19932 18158
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 16182 20024 18022
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19706 12744 19762 12753
rect 19706 12679 19762 12688
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19720 11558 19748 12106
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11830 19840 12038
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19904 11558 19932 15302
rect 19996 13734 20024 15982
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19996 12646 20024 13330
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 20088 12434 20116 17682
rect 20180 17082 20208 19178
rect 20272 17338 20300 21286
rect 20456 20602 20484 22170
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20732 21894 20760 22034
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20180 17054 20300 17082
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16794 20208 16934
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20272 14770 20300 17054
rect 20364 16794 20392 19654
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20180 14742 20300 14770
rect 20180 14657 20208 14742
rect 20166 14648 20222 14657
rect 20166 14583 20222 14592
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20180 13530 20208 14214
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 19996 12406 20116 12434
rect 19996 12170 20024 12406
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 20074 11792 20130 11801
rect 20074 11727 20130 11736
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19628 11036 19735 11064
rect 19614 10976 19670 10985
rect 19707 10962 19735 11036
rect 19812 11014 19840 11154
rect 19800 11008 19852 11014
rect 19707 10934 19748 10962
rect 19800 10950 19852 10956
rect 19614 10911 19670 10920
rect 19628 9450 19656 10911
rect 19720 10606 19748 10934
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19904 10418 19932 11154
rect 20088 11082 20116 11727
rect 20166 11384 20222 11393
rect 20166 11319 20222 11328
rect 20180 11150 20208 11319
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20088 10962 20116 11018
rect 20088 10934 20208 10962
rect 20074 10840 20130 10849
rect 20180 10810 20208 10934
rect 20074 10775 20076 10784
rect 20128 10775 20130 10784
rect 20168 10804 20220 10810
rect 20076 10746 20128 10752
rect 20168 10746 20220 10752
rect 19812 10390 19932 10418
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 9160 19748 9318
rect 19628 9132 19748 9160
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19628 5642 19656 9132
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19720 5846 19748 8978
rect 19708 5840 19760 5846
rect 19708 5782 19760 5788
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19812 3534 19840 10390
rect 19890 10296 19946 10305
rect 19890 10231 19946 10240
rect 19984 10260 20036 10266
rect 19904 10130 19932 10231
rect 19984 10202 20036 10208
rect 19996 10146 20024 10202
rect 19892 10124 19944 10130
rect 19996 10118 20208 10146
rect 19892 10066 19944 10072
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 5234 19932 9862
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19996 8566 20024 8910
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20088 7206 20116 9998
rect 20180 9926 20208 10118
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20180 8566 20208 9590
rect 20168 8560 20220 8566
rect 20168 8502 20220 8508
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 19352 2650 19380 2926
rect 20272 2774 20300 14554
rect 20456 14006 20484 18022
rect 20548 15502 20576 21626
rect 20628 21616 20680 21622
rect 20904 21616 20956 21622
rect 20680 21576 20904 21604
rect 20628 21558 20680 21564
rect 20904 21558 20956 21564
rect 21008 21486 21036 22918
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21100 21962 21128 22714
rect 21192 22234 21220 23122
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21100 20874 21128 21898
rect 21192 21146 21220 22170
rect 21284 22137 21312 23258
rect 21730 23080 21786 23089
rect 21640 23044 21692 23050
rect 21730 23015 21786 23024
rect 21640 22986 21692 22992
rect 21652 22778 21680 22986
rect 21640 22772 21692 22778
rect 21640 22714 21692 22720
rect 21362 22672 21418 22681
rect 21362 22607 21418 22616
rect 21376 22574 21404 22607
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21456 22432 21508 22438
rect 21456 22374 21508 22380
rect 21270 22128 21326 22137
rect 21270 22063 21326 22072
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21284 21026 21312 21830
rect 21468 21622 21496 22374
rect 21744 21622 21772 23015
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21192 20998 21312 21026
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 21100 20602 21128 20810
rect 21192 20806 21220 20998
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20732 20058 20760 20334
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20732 19786 20760 19994
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20626 19680 20682 19689
rect 20626 19615 20682 19624
rect 20640 17066 20668 19615
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 20718 19408 20774 19417
rect 20718 19343 20774 19352
rect 21008 19360 21036 19450
rect 21088 19372 21140 19378
rect 20732 18698 20760 19343
rect 21008 19332 21088 19360
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20732 17921 20760 18090
rect 20718 17912 20774 17921
rect 20718 17847 20774 17856
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20824 16998 20852 19178
rect 20902 18728 20958 18737
rect 20902 18663 20958 18672
rect 20916 18222 20944 18663
rect 21008 18630 21036 19332
rect 21088 19314 21140 19320
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20824 14958 20852 16934
rect 21008 16250 21036 18566
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20996 16040 21048 16046
rect 20994 16008 20996 16017
rect 21048 16008 21050 16017
rect 20994 15943 21050 15952
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20640 13802 20668 14894
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14550 20760 14758
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20732 13938 20760 14350
rect 20824 14074 20852 14350
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 20640 13530 20668 13738
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 12434 20392 12582
rect 20364 12406 20484 12434
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20364 10810 20392 11494
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20350 8392 20406 8401
rect 20350 8327 20406 8336
rect 20364 7750 20392 8327
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20352 6724 20404 6730
rect 20352 6666 20404 6672
rect 20364 6458 20392 6666
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20456 6322 20484 12406
rect 20548 8566 20576 12786
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20640 12102 20668 12650
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20640 9586 20668 11086
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20732 8498 20760 13670
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 12238 20852 12582
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20824 11762 20852 12174
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20824 11218 20852 11698
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20640 5710 20668 8298
rect 20824 6798 20852 10474
rect 20916 10130 20944 15302
rect 20994 14376 21050 14385
rect 20994 14311 21050 14320
rect 21008 14074 21036 14311
rect 21100 14278 21128 18158
rect 21192 15570 21220 19450
rect 21284 19281 21312 20810
rect 21376 20330 21404 21082
rect 21468 21078 21496 21558
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 21548 21412 21600 21418
rect 21548 21354 21600 21360
rect 21456 21072 21508 21078
rect 21456 21014 21508 21020
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 21376 19310 21404 19722
rect 21364 19304 21416 19310
rect 21270 19272 21326 19281
rect 21364 19246 21416 19252
rect 21270 19207 21326 19216
rect 21376 18698 21404 19246
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21376 17134 21404 18634
rect 21468 18086 21496 20742
rect 21560 18426 21588 21354
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21652 19718 21680 20946
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21652 18834 21680 19654
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21652 18426 21680 18566
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21100 13462 21128 14214
rect 21192 13870 21220 15370
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21088 13456 21140 13462
rect 21088 13398 21140 13404
rect 21284 12434 21312 15982
rect 21376 15570 21404 16390
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 12646 21404 14758
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21192 12406 21312 12434
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 21008 11830 21036 12242
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 21192 11558 21220 12406
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20916 9761 20944 9930
rect 20902 9752 20958 9761
rect 20902 9687 20958 9696
rect 20916 9586 20944 9687
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 21008 9178 21036 11086
rect 21086 10296 21142 10305
rect 21086 10231 21142 10240
rect 21100 9586 21128 10231
rect 21192 9994 21220 11494
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21284 10577 21312 10610
rect 21270 10568 21326 10577
rect 21270 10503 21326 10512
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21284 9602 21312 10503
rect 21376 10130 21404 12242
rect 21468 12238 21496 16730
rect 21560 15162 21588 18362
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21652 17134 21680 17546
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21744 16454 21772 21422
rect 21836 20602 21864 23598
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 21928 21894 21956 23530
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 21928 20890 21956 21830
rect 22112 21457 22140 24647
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22296 23662 22324 24142
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 22204 23050 22232 23530
rect 22296 23186 22324 23598
rect 22388 23322 22416 26302
rect 22650 26200 22706 26302
rect 22848 26302 23074 26330
rect 22742 24440 22798 24449
rect 22742 24375 22798 24384
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22480 23644 22508 24074
rect 22560 23656 22612 23662
rect 22480 23616 22560 23644
rect 22560 23598 22612 23604
rect 22572 23322 22600 23598
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22664 23202 22692 24210
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22572 23174 22692 23202
rect 22466 23080 22522 23089
rect 22192 23044 22244 23050
rect 22466 23015 22522 23024
rect 22192 22986 22244 22992
rect 22204 21962 22232 22986
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22098 21448 22154 21457
rect 22098 21383 22154 21392
rect 22296 20890 22324 22510
rect 22388 21894 22416 22714
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 21928 20862 22048 20890
rect 22020 20806 22048 20862
rect 22112 20862 22324 20890
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21836 18970 21864 19110
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21836 16114 21864 16526
rect 21928 16250 21956 20742
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22020 19417 22048 20538
rect 22006 19408 22062 19417
rect 22112 19378 22140 20862
rect 22282 20360 22338 20369
rect 22282 20295 22338 20304
rect 22190 19408 22246 19417
rect 22006 19343 22062 19352
rect 22100 19372 22152 19378
rect 22190 19343 22192 19352
rect 22100 19314 22152 19320
rect 22244 19343 22246 19352
rect 22192 19314 22244 19320
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 22020 19174 22048 19246
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21638 15464 21694 15473
rect 21638 15399 21694 15408
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21560 14414 21588 15098
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21560 11898 21588 14214
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21560 11558 21588 11698
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21192 9574 21312 9602
rect 21454 9616 21510 9625
rect 21192 9466 21220 9574
rect 21454 9551 21456 9560
rect 21508 9551 21510 9560
rect 21456 9522 21508 9528
rect 21100 9438 21220 9466
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 21100 8974 21128 9438
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20916 7886 20944 8298
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 7410 20944 7686
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 21192 4554 21220 7210
rect 21284 6866 21312 9318
rect 21468 9042 21496 9318
rect 21560 9178 21588 11494
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21364 8968 21416 8974
rect 21548 8968 21600 8974
rect 21364 8910 21416 8916
rect 21468 8916 21548 8922
rect 21468 8910 21600 8916
rect 21376 8022 21404 8910
rect 21468 8894 21588 8910
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21468 5370 21496 8894
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21560 7886 21588 8774
rect 21652 8430 21680 15399
rect 21730 14512 21786 14521
rect 22020 14482 22048 19110
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22204 17882 22232 18566
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22112 14618 22140 17206
rect 22204 16046 22232 17818
rect 22296 17338 22324 20295
rect 22388 19990 22416 21830
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 22480 19009 22508 23015
rect 22572 21894 22600 23174
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22664 22030 22692 22578
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22572 20097 22600 20334
rect 22558 20088 22614 20097
rect 22558 20023 22614 20032
rect 22466 19000 22522 19009
rect 22466 18935 22522 18944
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22296 17202 22324 17274
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 21730 14447 21786 14456
rect 22008 14476 22060 14482
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21652 7886 21680 8230
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21744 7410 21772 14447
rect 22008 14418 22060 14424
rect 22204 13938 22232 15302
rect 22296 14958 22324 16594
rect 22388 15366 22416 17274
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22296 14618 22324 14894
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22296 13938 22324 14554
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21560 7002 21588 7278
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21836 5778 21864 13874
rect 22296 13818 22324 13874
rect 22112 13790 22324 13818
rect 22006 13424 22062 13433
rect 22006 13359 22062 13368
rect 22020 11150 22048 13359
rect 22112 13258 22140 13790
rect 22192 13728 22244 13734
rect 22190 13696 22192 13705
rect 22244 13696 22246 13705
rect 22388 13682 22416 15030
rect 22480 14226 22508 18770
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22572 17746 22600 18294
rect 22664 17882 22692 20334
rect 22756 18816 22784 24375
rect 22848 22438 22876 26302
rect 23018 26200 23074 26302
rect 23308 26302 23442 26330
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23020 24132 23072 24138
rect 23020 24074 23072 24080
rect 23032 23798 23060 24074
rect 23020 23792 23072 23798
rect 23020 23734 23072 23740
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23308 23338 23336 26302
rect 23386 26200 23442 26302
rect 24490 26200 24546 27000
rect 24858 26200 24914 27000
rect 24950 26480 25006 26489
rect 24950 26415 25006 26424
rect 24398 26072 24454 26081
rect 24398 26007 24454 26016
rect 24214 25528 24270 25537
rect 24214 25463 24270 25472
rect 23386 25120 23442 25129
rect 23386 25055 23442 25064
rect 23400 24449 23428 25055
rect 24124 24608 24176 24614
rect 24124 24550 24176 24556
rect 23386 24440 23442 24449
rect 23386 24375 23442 24384
rect 23756 24404 23808 24410
rect 23756 24346 23808 24352
rect 23308 23310 23428 23338
rect 23400 23225 23428 23310
rect 23386 23216 23442 23225
rect 23296 23180 23348 23186
rect 23386 23151 23442 23160
rect 23296 23122 23348 23128
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22940 22710 22968 22918
rect 22928 22704 22980 22710
rect 22928 22646 22980 22652
rect 23308 22574 23336 23122
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 21554 23336 22510
rect 23386 22400 23442 22409
rect 23386 22335 23442 22344
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22848 18970 22876 21286
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23204 20868 23256 20874
rect 23204 20810 23256 20816
rect 23216 20602 23244 20810
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 23308 20466 23336 21490
rect 23400 21457 23428 22335
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23386 21448 23442 21457
rect 23386 21383 23442 21392
rect 23492 21010 23520 21898
rect 23676 21690 23704 22986
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23768 21350 23796 24346
rect 24136 24070 24164 24550
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 23860 23730 23888 24006
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 23940 23248 23992 23254
rect 23940 23190 23992 23196
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23860 21962 23888 22646
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23492 20602 23520 20946
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23308 19922 23336 20402
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23308 19378 23336 19858
rect 23400 19854 23428 20538
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23388 19848 23440 19854
rect 23386 19816 23388 19825
rect 23440 19816 23442 19825
rect 23386 19751 23442 19760
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22756 18788 22968 18816
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18426 22784 18566
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22572 17202 22600 17682
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22664 16658 22692 17818
rect 22756 17610 22784 18362
rect 22848 17762 22876 18634
rect 22940 18358 22968 18788
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 23216 18193 23244 18634
rect 23308 18426 23336 19314
rect 23400 19145 23428 19450
rect 23386 19136 23442 19145
rect 23386 19071 23442 19080
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23400 18737 23428 18838
rect 23386 18728 23442 18737
rect 23386 18663 23442 18672
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23386 18320 23442 18329
rect 23386 18255 23388 18264
rect 23440 18255 23442 18264
rect 23388 18226 23440 18232
rect 23202 18184 23258 18193
rect 23202 18119 23258 18128
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 22926 17776 22982 17785
rect 22848 17734 22926 17762
rect 22926 17711 22928 17720
rect 22980 17711 22982 17720
rect 22928 17682 22980 17688
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22848 17270 22876 17614
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22940 17270 22968 17478
rect 23032 17338 23060 17818
rect 23202 17776 23258 17785
rect 23202 17711 23258 17720
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 22836 17264 22888 17270
rect 22836 17206 22888 17212
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 22940 17134 22968 17206
rect 22928 17128 22980 17134
rect 23216 17105 23244 17711
rect 22928 17070 22980 17076
rect 23202 17096 23258 17105
rect 23202 17031 23258 17040
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23400 16810 23428 18022
rect 23308 16782 23428 16810
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22572 15502 22600 15846
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22572 14550 22600 15302
rect 22560 14544 22612 14550
rect 22664 14521 22692 16186
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 23204 16108 23256 16114
rect 23308 16096 23336 16782
rect 23386 16688 23442 16697
rect 23386 16623 23442 16632
rect 23256 16068 23336 16096
rect 23204 16050 23256 16056
rect 22560 14486 22612 14492
rect 22650 14512 22706 14521
rect 22756 14482 22784 16050
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22650 14447 22706 14456
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22848 14362 22876 15574
rect 23308 15570 23336 15846
rect 23400 15706 23428 16623
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23400 15502 23428 15642
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23492 14482 23520 19654
rect 23584 17746 23612 19994
rect 23676 18873 23704 20742
rect 23768 20534 23796 21286
rect 23860 20806 23888 21626
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23754 19544 23810 19553
rect 23754 19479 23810 19488
rect 23662 18864 23718 18873
rect 23662 18799 23718 18808
rect 23676 18426 23704 18799
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23768 18086 23796 19479
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23584 17134 23612 17682
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23676 16590 23704 17274
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 22664 14334 22876 14362
rect 22480 14198 22600 14226
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22190 13631 22246 13640
rect 22296 13654 22416 13682
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22112 12986 22140 13194
rect 22204 12986 22232 13194
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22112 12594 22140 12922
rect 22112 12566 22232 12594
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22112 10674 22140 12378
rect 22204 12306 22232 12566
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22296 11898 22324 13654
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22388 12442 22416 12854
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 21928 7410 21956 10474
rect 22006 9072 22062 9081
rect 22006 9007 22008 9016
rect 22060 9007 22062 9016
rect 22008 8978 22060 8984
rect 22204 8838 22232 11834
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22204 8090 22232 8434
rect 22296 8430 22324 11698
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 22020 6322 22048 7686
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 22480 5234 22508 14010
rect 22572 12918 22600 14198
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22664 12730 22692 14334
rect 22744 14272 22796 14278
rect 23296 14272 23348 14278
rect 22744 14214 22796 14220
rect 22834 14240 22890 14249
rect 22572 12702 22692 12730
rect 22572 5710 22600 12702
rect 22756 11626 22784 14214
rect 23296 14214 23348 14220
rect 22834 14175 22890 14184
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22664 10266 22692 11086
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 5914 22692 6734
rect 22652 5908 22704 5914
rect 22652 5850 22704 5856
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22756 4690 22784 10134
rect 22848 6798 22876 14175
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23308 10130 23336 14214
rect 23480 13184 23532 13190
rect 23400 13144 23480 13172
rect 23400 12850 23428 13144
rect 23480 13126 23532 13132
rect 23584 12889 23612 15302
rect 23676 15076 23704 16526
rect 23768 15337 23796 17478
rect 23860 16250 23888 20198
rect 23952 17678 23980 23190
rect 24044 20942 24072 23734
rect 24136 22982 24164 24006
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24124 21956 24176 21962
rect 24124 21898 24176 21904
rect 24136 21622 24164 21898
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24122 21176 24178 21185
rect 24122 21111 24178 21120
rect 24032 20936 24084 20942
rect 24136 20913 24164 21111
rect 24032 20878 24084 20884
rect 24122 20904 24178 20913
rect 24122 20839 24178 20848
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 24044 19446 24072 20470
rect 24136 19718 24164 20742
rect 24228 20058 24256 25463
rect 24306 24984 24362 24993
rect 24306 24919 24362 24928
rect 24320 23322 24348 24919
rect 24412 23798 24440 26007
rect 24400 23792 24452 23798
rect 24400 23734 24452 23740
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24308 23316 24360 23322
rect 24308 23258 24360 23264
rect 24308 22976 24360 22982
rect 24308 22918 24360 22924
rect 24320 22778 24348 22918
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24412 19718 24440 23462
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23940 17672 23992 17678
rect 24044 17649 24072 18022
rect 24136 17814 24164 19654
rect 24412 19292 24440 19654
rect 24320 19264 24440 19292
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24320 18034 24348 19264
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24412 18222 24440 18566
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24124 17808 24176 17814
rect 24124 17750 24176 17756
rect 23940 17614 23992 17620
rect 24030 17640 24086 17649
rect 24030 17575 24086 17584
rect 24044 17320 24072 17575
rect 24124 17332 24176 17338
rect 24044 17292 24124 17320
rect 24124 17274 24176 17280
rect 24228 17202 24256 18022
rect 24320 18006 24440 18034
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23952 16046 23980 16390
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23754 15328 23810 15337
rect 23754 15263 23810 15272
rect 23952 15162 23980 15982
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 23756 15088 23808 15094
rect 23676 15048 23756 15076
rect 23756 15030 23808 15036
rect 23768 14346 23796 15030
rect 23756 14340 23808 14346
rect 23756 14282 23808 14288
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23570 12880 23626 12889
rect 23388 12844 23440 12850
rect 23570 12815 23626 12824
rect 23388 12786 23440 12792
rect 23400 12102 23428 12786
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23400 9926 23428 10066
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23294 9752 23350 9761
rect 23294 9687 23350 9696
rect 23308 9654 23336 9687
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22848 5710 22876 6598
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 21180 4548 21232 4554
rect 21180 4490 21232 4496
rect 23308 4162 23336 6666
rect 23216 4134 23336 4162
rect 23216 4078 23244 4134
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 20180 2746 20300 2774
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 800 20208 2746
rect 22020 1170 22048 3402
rect 22112 1601 22140 4014
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22296 3058 22324 3334
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23400 2650 23428 9862
rect 23492 9178 23520 9998
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23492 8838 23520 9114
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23676 6458 23704 14214
rect 23768 14006 23796 14282
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23756 14000 23808 14006
rect 23756 13942 23808 13948
rect 23768 13190 23796 13942
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23860 11665 23888 14214
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23846 11656 23902 11665
rect 23846 11591 23902 11600
rect 23952 6798 23980 11698
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23492 3602 23520 6054
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 24044 3058 24072 9930
rect 24136 8906 24164 17002
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24320 13870 24348 14418
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24216 13796 24268 13802
rect 24216 13738 24268 13744
rect 24228 12850 24256 13738
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24124 8900 24176 8906
rect 24124 8842 24176 8848
rect 24228 8090 24256 12786
rect 24320 12306 24348 13806
rect 24412 13297 24440 18006
rect 24504 17066 24532 26200
rect 24766 24848 24822 24857
rect 24766 24783 24822 24792
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24596 23633 24624 24006
rect 24688 23866 24716 24006
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24780 23633 24808 24783
rect 24582 23624 24638 23633
rect 24582 23559 24638 23568
rect 24766 23624 24822 23633
rect 24766 23559 24822 23568
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24872 21486 24900 22714
rect 24964 22574 24992 26415
rect 25226 26200 25282 27000
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 24952 22568 25004 22574
rect 24952 22510 25004 22516
rect 24952 22024 25004 22030
rect 24950 21992 24952 22001
rect 25004 21992 25006 22001
rect 24950 21927 25006 21936
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24582 21176 24638 21185
rect 24582 21111 24638 21120
rect 24596 20874 24624 21111
rect 24676 21072 24728 21078
rect 24676 21014 24728 21020
rect 24584 20868 24636 20874
rect 24584 20810 24636 20816
rect 24688 20641 24716 21014
rect 24674 20632 24730 20641
rect 24674 20567 24730 20576
rect 25056 20074 25084 24142
rect 25148 23798 25176 25191
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 24964 20046 25084 20074
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24688 18630 24716 18906
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24596 18057 24624 18566
rect 24582 18048 24638 18057
rect 24582 17983 24638 17992
rect 24674 17096 24730 17105
rect 24492 17060 24544 17066
rect 24674 17031 24730 17040
rect 24492 17002 24544 17008
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24596 15638 24624 16050
rect 24584 15632 24636 15638
rect 24584 15574 24636 15580
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24398 13288 24454 13297
rect 24398 13223 24454 13232
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 24412 10606 24440 13126
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 24504 8022 24532 14350
rect 24582 13832 24638 13841
rect 24688 13802 24716 17031
rect 24780 15162 24808 19858
rect 24964 17882 24992 20046
rect 25042 19952 25098 19961
rect 25042 19887 25044 19896
rect 25096 19887 25098 19896
rect 25044 19858 25096 19864
rect 25148 19514 25176 23122
rect 25240 22778 25268 24210
rect 25780 23792 25832 23798
rect 25780 23734 25832 23740
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25228 22500 25280 22506
rect 25228 22442 25280 22448
rect 25240 21962 25268 22442
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25240 19310 25268 20198
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 25056 18086 25084 18770
rect 25148 18766 25176 19110
rect 25240 18834 25268 19246
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25332 18222 25360 23666
rect 25504 23112 25556 23118
rect 25504 23054 25556 23060
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 25424 21894 25452 22374
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25412 21344 25464 21350
rect 25412 21286 25464 21292
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24872 16289 24900 16526
rect 24858 16280 24914 16289
rect 24858 16215 24914 16224
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24780 14074 24808 15098
rect 24858 14648 24914 14657
rect 24858 14583 24914 14592
rect 24872 14414 24900 14583
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24964 14226 24992 16118
rect 25228 15904 25280 15910
rect 25424 15881 25452 21286
rect 25516 16590 25544 23054
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25608 17746 25636 22918
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25700 17134 25728 19450
rect 25688 17128 25740 17134
rect 25688 17070 25740 17076
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25686 16280 25742 16289
rect 25686 16215 25742 16224
rect 25228 15846 25280 15852
rect 25410 15872 25466 15881
rect 25240 15609 25268 15846
rect 25410 15807 25466 15816
rect 25226 15600 25282 15609
rect 25226 15535 25282 15544
rect 25424 15502 25452 15807
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25134 15192 25190 15201
rect 25134 15127 25190 15136
rect 25148 15094 25176 15127
rect 25136 15088 25188 15094
rect 25188 15048 25268 15076
rect 25136 15030 25188 15036
rect 24872 14198 24992 14226
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24582 13767 24638 13776
rect 24676 13796 24728 13802
rect 24596 12238 24624 13767
rect 24676 13738 24728 13744
rect 24674 13016 24730 13025
rect 24674 12951 24730 12960
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 9178 24624 12174
rect 24688 11150 24716 12951
rect 24766 12200 24822 12209
rect 24766 12135 24822 12144
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24674 10976 24730 10985
rect 24674 10911 24730 10920
rect 24688 9518 24716 10911
rect 24780 10606 24808 12135
rect 24872 11914 24900 14198
rect 25134 13968 25190 13977
rect 25134 13903 25136 13912
rect 25188 13903 25190 13912
rect 25136 13874 25188 13880
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24964 12102 24992 12582
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24872 11886 24992 11914
rect 24860 11824 24912 11830
rect 24858 11792 24860 11801
rect 24912 11792 24914 11801
rect 24858 11727 24914 11736
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24872 11218 24900 11319
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24768 10600 24820 10606
rect 24872 10577 24900 10678
rect 24768 10542 24820 10548
rect 24858 10568 24914 10577
rect 24858 10503 24914 10512
rect 24766 10160 24822 10169
rect 24766 10095 24822 10104
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24780 8430 24808 10095
rect 24964 10062 24992 11886
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24872 9042 24900 9279
rect 24964 9110 24992 9862
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24860 8560 24912 8566
rect 24858 8528 24860 8537
rect 24912 8528 24914 8537
rect 24858 8463 24914 8472
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24858 8120 24914 8129
rect 24858 8055 24914 8064
rect 24492 8016 24544 8022
rect 24492 7958 24544 7964
rect 24872 7954 24900 8055
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7274 24716 7822
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24676 7268 24728 7274
rect 24676 7210 24728 7216
rect 24584 6928 24636 6934
rect 24584 6870 24636 6876
rect 24596 6730 24624 6870
rect 24584 6724 24636 6730
rect 24584 6666 24636 6672
rect 24674 6488 24730 6497
rect 24674 6423 24730 6432
rect 24688 5166 24716 6423
rect 24780 6254 24808 7647
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24872 7313 24900 7414
rect 24858 7304 24914 7313
rect 24858 7239 24914 7248
rect 24964 7154 24992 7754
rect 24872 7126 24992 7154
rect 24872 6798 24900 7126
rect 25056 6934 25084 13806
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25148 12986 25176 13330
rect 25240 12986 25268 15048
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25504 14816 25556 14822
rect 25504 14758 25556 14764
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25134 12608 25190 12617
rect 25134 12543 25190 12552
rect 25148 11830 25176 12543
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25148 9178 25176 11154
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 25148 7478 25176 8871
rect 25240 8362 25268 12038
rect 25424 11218 25452 13874
rect 25412 11212 25464 11218
rect 25412 11154 25464 11160
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 25044 6928 25096 6934
rect 24950 6896 25006 6905
rect 25044 6870 25096 6876
rect 24950 6831 24952 6840
rect 25004 6831 25006 6840
rect 24952 6802 25004 6808
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24872 6089 24900 6326
rect 24858 6080 24914 6089
rect 24858 6015 24914 6024
rect 24952 5704 25004 5710
rect 24950 5672 24952 5681
rect 25004 5672 25006 5681
rect 24950 5607 25006 5616
rect 25044 5636 25096 5642
rect 25044 5578 25096 5584
rect 24860 5296 24912 5302
rect 24766 5264 24822 5273
rect 24860 5238 24912 5244
rect 24766 5199 24822 5208
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 22848 2009 22876 2586
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 22834 2000 22890 2009
rect 22834 1935 22890 1944
rect 22098 1592 22154 1601
rect 22098 1527 22154 1536
rect 22098 1184 22154 1193
rect 22020 1142 22098 1170
rect 22098 1119 22154 1128
rect 6734 0 6790 800
rect 20166 0 20222 800
rect 23400 377 23428 2450
rect 24596 2446 24624 4694
rect 24688 3534 24716 4694
rect 24780 4078 24808 5199
rect 24872 4865 24900 5238
rect 24858 4856 24914 4865
rect 24858 4791 24914 4800
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24964 4457 24992 4490
rect 24950 4448 25006 4457
rect 24950 4383 25006 4392
rect 25056 4146 25084 5578
rect 25148 4826 25176 7210
rect 25332 5914 25360 11086
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25424 7546 25452 11018
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25424 6866 25452 7346
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25516 4146 25544 14758
rect 25608 4690 25636 14826
rect 25700 6730 25728 16215
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25792 5846 25820 23734
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26054 21176 26110 21185
rect 26054 21111 26110 21120
rect 26068 20738 26096 21111
rect 26056 20732 26108 20738
rect 26056 20674 26108 20680
rect 26056 18896 26108 18902
rect 26056 18838 26108 18844
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25884 6322 25912 18022
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25976 10713 26004 15302
rect 26068 13462 26096 18838
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 25962 10704 26018 10713
rect 25962 10639 26018 10648
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 25872 6316 25924 6322
rect 25872 6258 25924 6264
rect 25780 5840 25832 5846
rect 25780 5782 25832 5788
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25134 4040 25190 4049
rect 24952 4004 25004 4010
rect 25134 3975 25190 3984
rect 24952 3946 25004 3952
rect 24964 3641 24992 3946
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24952 3460 25004 3466
rect 24952 3402 25004 3408
rect 24964 3233 24992 3402
rect 24950 3224 25006 3233
rect 24950 3159 25006 3168
rect 25148 3126 25176 3975
rect 25976 3194 26004 7754
rect 26068 4486 26096 13194
rect 26160 9654 26188 21830
rect 26424 20732 26476 20738
rect 26424 20674 26476 20680
rect 26148 9648 26200 9654
rect 26148 9590 26200 9596
rect 26436 9382 26464 20674
rect 26516 17060 26568 17066
rect 26516 17002 26568 17008
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 26160 7410 26188 8774
rect 26528 8634 26556 17002
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25136 3120 25188 3126
rect 25136 3062 25188 3068
rect 24872 2825 24900 3062
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24950 2408 25006 2417
rect 24950 2343 24952 2352
rect 25004 2343 25006 2352
rect 24952 2314 25004 2320
rect 25056 785 25084 2926
rect 25042 776 25098 785
rect 25042 711 25098 720
rect 23386 368 23442 377
rect 23386 303 23442 312
<< via2 >>
rect 1582 25880 1638 25936
rect 1490 23704 1546 23760
rect 1766 23704 1822 23760
rect 1858 23024 1914 23080
rect 1674 22616 1730 22672
rect 1766 21956 1822 21992
rect 1766 21936 1768 21956
rect 1768 21936 1820 21956
rect 1820 21936 1822 21956
rect 1766 21392 1822 21448
rect 2134 23024 2190 23080
rect 1950 17740 2006 17776
rect 1950 17720 1952 17740
rect 1952 17720 2004 17740
rect 2004 17720 2006 17740
rect 2134 17196 2190 17232
rect 2134 17176 2136 17196
rect 2136 17176 2188 17196
rect 2188 17176 2190 17196
rect 2134 16108 2190 16144
rect 2134 16088 2136 16108
rect 2136 16088 2188 16108
rect 2188 16088 2190 16108
rect 2594 20340 2596 20360
rect 2596 20340 2648 20360
rect 2648 20340 2650 20360
rect 2594 20304 2650 20340
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 3606 24792 3662 24848
rect 3606 20168 3662 20224
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3238 17584 3294 17640
rect 2778 17040 2834 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 3514 18944 3570 19000
rect 3882 16652 3938 16688
rect 3882 16632 3884 16652
rect 3884 16632 3936 16652
rect 3936 16632 3938 16652
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 4802 25608 4858 25664
rect 4066 18284 4122 18320
rect 4066 18264 4068 18284
rect 4068 18264 4120 18284
rect 4120 18264 4122 18284
rect 4250 16768 4306 16824
rect 4802 21548 4858 21584
rect 4802 21528 4804 21548
rect 4804 21528 4856 21548
rect 4856 21528 4858 21548
rect 4986 18844 4988 18864
rect 4988 18844 5040 18864
rect 5040 18844 5042 18864
rect 4986 18808 5042 18844
rect 4986 17992 5042 18048
rect 4802 17720 4858 17776
rect 5446 23160 5502 23216
rect 5538 22480 5594 22536
rect 5354 19896 5410 19952
rect 5630 19216 5686 19272
rect 5262 15580 5264 15600
rect 5264 15580 5316 15600
rect 5316 15580 5318 15600
rect 5262 15544 5318 15580
rect 4710 15408 4766 15464
rect 3882 14864 3938 14920
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 1950 13368 2006 13424
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 6182 26016 6238 26072
rect 5814 18672 5870 18728
rect 5722 16768 5778 16824
rect 5538 12144 5594 12200
rect 6274 24248 6330 24304
rect 6734 24148 6736 24168
rect 6736 24148 6788 24168
rect 6788 24148 6790 24168
rect 6734 24112 6790 24148
rect 6550 23432 6606 23488
rect 7010 24112 7066 24168
rect 6366 21256 6422 21312
rect 6826 20304 6882 20360
rect 5906 14456 5962 14512
rect 7010 19352 7066 19408
rect 7286 20052 7342 20088
rect 7286 20032 7288 20052
rect 7288 20032 7340 20052
rect 7340 20032 7342 20052
rect 7194 19760 7250 19816
rect 7286 19488 7342 19544
rect 7286 17720 7342 17776
rect 6918 16768 6974 16824
rect 6550 13912 6606 13968
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 7470 17720 7526 17776
rect 7286 16904 7342 16960
rect 7286 15952 7342 16008
rect 7102 13640 7158 13696
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 8666 25880 8722 25936
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8298 20984 8354 21040
rect 7838 20848 7894 20904
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 8390 19488 8446 19544
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7654 18148 7710 18184
rect 7654 18128 7656 18148
rect 7656 18128 7708 18148
rect 7708 18128 7710 18148
rect 7838 17856 7894 17912
rect 9218 24656 9274 24712
rect 9126 22616 9182 22672
rect 8758 21392 8814 21448
rect 8298 17720 8354 17776
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8298 16496 8354 16552
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8022 16108 8078 16144
rect 8022 16088 8024 16108
rect 8024 16088 8076 16108
rect 8076 16088 8078 16108
rect 7838 15972 7894 16008
rect 7838 15952 7840 15972
rect 7840 15952 7892 15972
rect 7892 15952 7894 15972
rect 8298 15852 8300 15872
rect 8300 15852 8352 15872
rect 8352 15852 8354 15872
rect 8298 15816 8354 15852
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 10230 25744 10286 25800
rect 9770 23432 9826 23488
rect 9402 22380 9404 22400
rect 9404 22380 9456 22400
rect 9456 22380 9458 22400
rect 9402 22344 9458 22380
rect 9402 21956 9458 21992
rect 9402 21936 9404 21956
rect 9404 21936 9456 21956
rect 9456 21936 9458 21956
rect 9402 20576 9458 20632
rect 9034 18808 9090 18864
rect 8758 17312 8814 17368
rect 8758 16904 8814 16960
rect 9034 16788 9090 16824
rect 9034 16768 9036 16788
rect 9036 16768 9088 16788
rect 9088 16768 9090 16788
rect 8666 13096 8722 13152
rect 8390 12688 8446 12744
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7010 11736 7066 11792
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 9310 18264 9366 18320
rect 9770 22208 9826 22264
rect 10322 24928 10378 24984
rect 9770 21664 9826 21720
rect 10046 21800 10102 21856
rect 9954 18400 10010 18456
rect 9494 16496 9550 16552
rect 10414 19760 10470 19816
rect 10230 18808 10286 18864
rect 10046 16768 10102 16824
rect 11058 23024 11114 23080
rect 11150 21664 11206 21720
rect 11058 20848 11114 20904
rect 10874 20168 10930 20224
rect 10782 19896 10838 19952
rect 10874 19760 10930 19816
rect 11334 20848 11390 20904
rect 11334 20440 11390 20496
rect 11058 18808 11114 18864
rect 10506 15020 10562 15056
rect 10506 15000 10508 15020
rect 10508 15000 10560 15020
rect 10560 15000 10562 15020
rect 10782 15272 10838 15328
rect 10966 15156 11022 15192
rect 10966 15136 10968 15156
rect 10968 15136 11020 15156
rect 11020 15136 11022 15156
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 11518 22380 11520 22400
rect 11520 22380 11572 22400
rect 11572 22380 11574 22400
rect 11518 22344 11574 22380
rect 11518 20440 11574 20496
rect 11886 21936 11942 21992
rect 12714 23432 12770 23488
rect 12346 22888 12402 22944
rect 11978 21256 12034 21312
rect 11426 18944 11482 19000
rect 11334 17040 11390 17096
rect 11610 18536 11666 18592
rect 11518 15680 11574 15736
rect 11426 15544 11482 15600
rect 11610 14068 11666 14104
rect 11610 14048 11612 14068
rect 11612 14048 11664 14068
rect 11664 14048 11666 14068
rect 10414 12960 10470 13016
rect 12714 22208 12770 22264
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13634 23024 13690 23080
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12254 20712 12310 20768
rect 12438 20596 12494 20632
rect 12438 20576 12440 20596
rect 12440 20576 12492 20596
rect 12492 20576 12494 20596
rect 11886 15680 11942 15736
rect 11886 14728 11942 14784
rect 12070 14320 12126 14376
rect 12530 17992 12586 18048
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12622 17856 12678 17912
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 13818 21936 13874 21992
rect 13634 20984 13690 21040
rect 14094 23296 14150 23352
rect 14094 22752 14150 22808
rect 14554 22752 14610 22808
rect 14554 22344 14610 22400
rect 13542 20168 13598 20224
rect 13818 20168 13874 20224
rect 13542 19624 13598 19680
rect 13726 19624 13782 19680
rect 13542 19352 13598 19408
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13358 18944 13414 19000
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12438 17484 12440 17504
rect 12440 17484 12492 17504
rect 12492 17484 12494 17504
rect 12438 17448 12494 17484
rect 12346 15852 12348 15872
rect 12348 15852 12400 15872
rect 12400 15852 12402 15872
rect 12346 15816 12402 15852
rect 12622 14728 12678 14784
rect 12346 13232 12402 13288
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13358 15272 13414 15328
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12714 10512 12770 10568
rect 14370 21120 14426 21176
rect 14186 20168 14242 20224
rect 13910 14728 13966 14784
rect 13818 14592 13874 14648
rect 13726 13796 13782 13832
rect 13726 13776 13728 13796
rect 13728 13776 13780 13796
rect 13780 13776 13782 13796
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 14186 16224 14242 16280
rect 14278 15680 14334 15736
rect 14646 19080 14702 19136
rect 14554 18264 14610 18320
rect 14462 17856 14518 17912
rect 14462 15408 14518 15464
rect 14646 15680 14702 15736
rect 14462 13776 14518 13832
rect 14922 22500 14978 22536
rect 14922 22480 14924 22500
rect 14924 22480 14976 22500
rect 14976 22480 14978 22500
rect 15198 24384 15254 24440
rect 15198 24112 15254 24168
rect 15014 22344 15070 22400
rect 15014 20984 15070 21040
rect 15566 24520 15622 24576
rect 15290 20440 15346 20496
rect 15290 19488 15346 19544
rect 15014 18536 15070 18592
rect 15014 17176 15070 17232
rect 15198 12280 15254 12336
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 15658 22888 15714 22944
rect 15474 21392 15530 21448
rect 16394 24384 16450 24440
rect 15934 23160 15990 23216
rect 15658 17176 15714 17232
rect 15842 20748 15844 20768
rect 15844 20748 15896 20768
rect 15896 20748 15898 20768
rect 15842 20712 15898 20748
rect 15842 16360 15898 16416
rect 15750 15816 15806 15872
rect 15658 13096 15714 13152
rect 15842 11872 15898 11928
rect 16210 22888 16266 22944
rect 16302 21412 16358 21448
rect 16302 21392 16304 21412
rect 16304 21392 16356 21412
rect 16356 21392 16358 21412
rect 16210 20304 16266 20360
rect 16210 17176 16266 17232
rect 16210 15544 16266 15600
rect 16486 20712 16542 20768
rect 16486 18400 16542 18456
rect 16946 24404 17002 24440
rect 16946 24384 16948 24404
rect 16948 24384 17000 24404
rect 17000 24384 17002 24404
rect 16762 22752 16818 22808
rect 16762 22480 16818 22536
rect 16762 21956 16818 21992
rect 16762 21936 16764 21956
rect 16764 21936 16816 21956
rect 16816 21936 16818 21956
rect 16670 20168 16726 20224
rect 16854 20168 16910 20224
rect 16762 19796 16764 19816
rect 16764 19796 16816 19816
rect 16816 19796 16818 19816
rect 16762 19760 16818 19796
rect 16762 18808 16818 18864
rect 17866 24656 17922 24712
rect 17958 24112 18014 24168
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17498 23432 17554 23488
rect 18142 23432 18198 23488
rect 17314 23024 17370 23080
rect 17682 22924 17684 22944
rect 17684 22924 17736 22944
rect 17736 22924 17738 22944
rect 16210 12960 16266 13016
rect 16302 10668 16358 10704
rect 16302 10648 16304 10668
rect 16304 10648 16356 10668
rect 16356 10648 16358 10668
rect 16762 14456 16818 14512
rect 16670 13504 16726 13560
rect 16670 13232 16726 13288
rect 16762 12844 16818 12880
rect 16762 12824 16764 12844
rect 16764 12824 16816 12844
rect 16816 12824 16818 12844
rect 16670 12416 16726 12472
rect 17682 22888 17738 22924
rect 18142 23160 18198 23216
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 18878 24520 18934 24576
rect 18326 22208 18382 22264
rect 17590 21664 17646 21720
rect 17498 21548 17554 21584
rect 17498 21528 17500 21548
rect 17500 21528 17552 21548
rect 17552 21528 17554 21548
rect 17406 20576 17462 20632
rect 17406 19896 17462 19952
rect 17406 19352 17462 19408
rect 17222 17312 17278 17368
rect 17130 16768 17186 16824
rect 17222 14864 17278 14920
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17774 19352 17830 19408
rect 17682 17992 17738 18048
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18694 21120 18750 21176
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17590 15408 17646 15464
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18694 17176 18750 17232
rect 18786 16496 18842 16552
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 17406 11348 17462 11384
rect 17406 11328 17408 11348
rect 17408 11328 17460 11348
rect 17460 11328 17462 11348
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18602 13640 18658 13696
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17866 11056 17922 11112
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18694 12164 18750 12200
rect 18694 12144 18696 12164
rect 18696 12144 18748 12164
rect 18748 12144 18750 12164
rect 19246 23432 19302 23488
rect 19430 25336 19486 25392
rect 19430 22480 19486 22536
rect 19614 23432 19670 23488
rect 20442 26016 20498 26072
rect 20626 25608 20682 25664
rect 19890 23432 19946 23488
rect 20166 23432 20222 23488
rect 20626 23724 20682 23760
rect 20626 23704 20628 23724
rect 20628 23704 20680 23724
rect 20680 23704 20682 23724
rect 21270 26152 21326 26208
rect 22190 26288 22246 26344
rect 21914 25880 21970 25936
rect 21178 25744 21234 25800
rect 22098 24656 22154 24712
rect 21270 24248 21326 24304
rect 20810 23296 20866 23352
rect 19522 20304 19578 20360
rect 19338 19760 19394 19816
rect 19522 19760 19578 19816
rect 19522 19352 19578 19408
rect 19062 19080 19118 19136
rect 19706 21664 19762 21720
rect 19982 20576 20038 20632
rect 19706 18264 19762 18320
rect 19522 16904 19578 16960
rect 18694 11192 18750 11248
rect 18602 11056 18658 11112
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17590 9424 17646 9480
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19246 12280 19302 12336
rect 19430 11600 19486 11656
rect 19430 11192 19486 11248
rect 19338 10784 19394 10840
rect 19430 9172 19486 9208
rect 19430 9152 19432 9172
rect 19432 9152 19484 9172
rect 19484 9152 19486 9172
rect 19706 12688 19762 12744
rect 20166 14592 20222 14648
rect 20074 11736 20130 11792
rect 19614 10920 19670 10976
rect 20166 11328 20222 11384
rect 20074 10804 20130 10840
rect 20074 10784 20076 10804
rect 20076 10784 20128 10804
rect 20128 10784 20130 10804
rect 19890 10240 19946 10296
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 21730 23024 21786 23080
rect 21362 22616 21418 22672
rect 21270 22072 21326 22128
rect 20626 19624 20682 19680
rect 20718 19352 20774 19408
rect 20718 17856 20774 17912
rect 20902 18672 20958 18728
rect 20994 15988 20996 16008
rect 20996 15988 21048 16008
rect 21048 15988 21050 16008
rect 20994 15952 21050 15988
rect 20350 8336 20406 8392
rect 20994 14320 21050 14376
rect 21270 19216 21326 19272
rect 20902 9696 20958 9752
rect 21086 10240 21142 10296
rect 21270 10512 21326 10568
rect 22742 24384 22798 24440
rect 22466 23024 22522 23080
rect 22098 21392 22154 21448
rect 22006 19352 22062 19408
rect 22282 20304 22338 20360
rect 22190 19372 22246 19408
rect 22190 19352 22192 19372
rect 22192 19352 22244 19372
rect 22244 19352 22246 19372
rect 21638 15408 21694 15464
rect 21454 9580 21510 9616
rect 21454 9560 21456 9580
rect 21456 9560 21508 9580
rect 21508 9560 21510 9580
rect 21730 14456 21786 14512
rect 22558 20032 22614 20088
rect 22466 18944 22522 19000
rect 22006 13368 22062 13424
rect 22190 13676 22192 13696
rect 22192 13676 22244 13696
rect 22244 13676 22246 13696
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 24950 26424 25006 26480
rect 24398 26016 24454 26072
rect 24214 25472 24270 25528
rect 23386 25064 23442 25120
rect 23386 24384 23442 24440
rect 23386 23160 23442 23216
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23386 22344 23442 22400
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23386 21392 23442 21448
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23386 19796 23388 19816
rect 23388 19796 23440 19816
rect 23440 19796 23442 19816
rect 23386 19760 23442 19796
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23386 19080 23442 19136
rect 23386 18672 23442 18728
rect 23386 18284 23442 18320
rect 23386 18264 23388 18284
rect 23388 18264 23440 18284
rect 23440 18264 23442 18284
rect 23202 18128 23258 18184
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22926 17740 22982 17776
rect 22926 17720 22928 17740
rect 22928 17720 22980 17740
rect 22980 17720 22982 17740
rect 23202 17720 23258 17776
rect 23202 17040 23258 17096
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23386 16632 23442 16688
rect 22650 14456 22706 14512
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 23754 19488 23810 19544
rect 23662 18808 23718 18864
rect 22190 13640 22246 13676
rect 22006 9036 22062 9072
rect 22006 9016 22008 9036
rect 22008 9016 22060 9036
rect 22060 9016 22062 9036
rect 22834 14184 22890 14240
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 24122 21120 24178 21176
rect 24122 20848 24178 20904
rect 24306 24928 24362 24984
rect 24030 17584 24086 17640
rect 23754 15272 23810 15328
rect 23570 12824 23626 12880
rect 23294 9696 23350 9752
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23846 11600 23902 11656
rect 24766 24792 24822 24848
rect 24582 23568 24638 23624
rect 24766 23568 24822 23624
rect 25134 25200 25190 25256
rect 24950 21972 24952 21992
rect 24952 21972 25004 21992
rect 25004 21972 25006 21992
rect 24950 21936 25006 21972
rect 24582 21120 24638 21176
rect 24674 20576 24730 20632
rect 24582 17992 24638 18048
rect 24674 17040 24730 17096
rect 24398 13232 24454 13288
rect 24582 13776 24638 13832
rect 25042 19916 25098 19952
rect 25042 19896 25044 19916
rect 25044 19896 25096 19916
rect 25096 19896 25098 19916
rect 24858 16224 24914 16280
rect 24858 14592 24914 14648
rect 25686 16224 25742 16280
rect 25410 15816 25466 15872
rect 25226 15544 25282 15600
rect 25134 15136 25190 15192
rect 24674 12960 24730 13016
rect 24766 12144 24822 12200
rect 24674 10920 24730 10976
rect 25134 13932 25190 13968
rect 25134 13912 25136 13932
rect 25136 13912 25188 13932
rect 25188 13912 25190 13932
rect 24858 11772 24860 11792
rect 24860 11772 24912 11792
rect 24912 11772 24914 11792
rect 24858 11736 24914 11772
rect 24858 11328 24914 11384
rect 24858 10512 24914 10568
rect 24766 10104 24822 10160
rect 24858 9288 24914 9344
rect 24858 8508 24860 8528
rect 24860 8508 24912 8528
rect 24912 8508 24914 8528
rect 24858 8472 24914 8508
rect 24858 8064 24914 8120
rect 24766 7656 24822 7712
rect 24674 6432 24730 6488
rect 24858 7248 24914 7304
rect 25134 12552 25190 12608
rect 25134 8880 25190 8936
rect 24950 6860 25006 6896
rect 24950 6840 24952 6860
rect 24952 6840 25004 6860
rect 25004 6840 25006 6860
rect 24858 6024 24914 6080
rect 24950 5652 24952 5672
rect 24952 5652 25004 5672
rect 25004 5652 25006 5672
rect 24950 5616 25006 5652
rect 24766 5208 24822 5264
rect 22834 1944 22890 2000
rect 22098 1536 22154 1592
rect 22098 1128 22154 1184
rect 24858 4800 24914 4856
rect 24950 4392 25006 4448
rect 26054 21120 26110 21176
rect 25962 10648 26018 10704
rect 25134 3984 25190 4040
rect 24950 3576 25006 3632
rect 24950 3168 25006 3224
rect 24858 2760 24914 2816
rect 24950 2372 25006 2408
rect 24950 2352 24952 2372
rect 24952 2352 25004 2372
rect 25004 2352 25006 2372
rect 25042 720 25098 776
rect 23386 312 23442 368
<< metal3 >>
rect 24945 26482 25011 26485
rect 26200 26482 27000 26512
rect 24945 26480 27000 26482
rect 24945 26424 24950 26480
rect 25006 26424 27000 26480
rect 24945 26422 27000 26424
rect 24945 26419 25011 26422
rect 26200 26392 27000 26422
rect 2262 26284 2268 26348
rect 2332 26346 2338 26348
rect 22185 26346 22251 26349
rect 2332 26344 22251 26346
rect 2332 26288 22190 26344
rect 22246 26288 22251 26344
rect 2332 26286 22251 26288
rect 2332 26284 2338 26286
rect 22185 26283 22251 26286
rect 4102 26148 4108 26212
rect 4172 26210 4178 26212
rect 21265 26210 21331 26213
rect 4172 26208 21331 26210
rect 4172 26152 21270 26208
rect 21326 26152 21331 26208
rect 4172 26150 21331 26152
rect 4172 26148 4178 26150
rect 21265 26147 21331 26150
rect 6177 26074 6243 26077
rect 20437 26074 20503 26077
rect 6177 26072 20503 26074
rect 6177 26016 6182 26072
rect 6238 26016 20442 26072
rect 20498 26016 20503 26072
rect 6177 26014 20503 26016
rect 6177 26011 6243 26014
rect 20437 26011 20503 26014
rect 24393 26074 24459 26077
rect 26200 26074 27000 26104
rect 24393 26072 27000 26074
rect 24393 26016 24398 26072
rect 24454 26016 27000 26072
rect 24393 26014 27000 26016
rect 24393 26011 24459 26014
rect 26200 25984 27000 26014
rect 0 25938 800 25968
rect 1577 25938 1643 25941
rect 0 25936 1643 25938
rect 0 25880 1582 25936
rect 1638 25880 1643 25936
rect 0 25878 1643 25880
rect 0 25848 800 25878
rect 1577 25875 1643 25878
rect 8661 25938 8727 25941
rect 21909 25938 21975 25941
rect 8661 25936 21975 25938
rect 8661 25880 8666 25936
rect 8722 25880 21914 25936
rect 21970 25880 21975 25936
rect 8661 25878 21975 25880
rect 8661 25875 8727 25878
rect 21909 25875 21975 25878
rect 10225 25802 10291 25805
rect 21173 25802 21239 25805
rect 10225 25800 21239 25802
rect 10225 25744 10230 25800
rect 10286 25744 21178 25800
rect 21234 25744 21239 25800
rect 10225 25742 21239 25744
rect 10225 25739 10291 25742
rect 21173 25739 21239 25742
rect 4797 25666 4863 25669
rect 19558 25666 19564 25668
rect 4797 25664 19564 25666
rect 4797 25608 4802 25664
rect 4858 25608 19564 25664
rect 4797 25606 19564 25608
rect 4797 25603 4863 25606
rect 19558 25604 19564 25606
rect 19628 25604 19634 25668
rect 20621 25666 20687 25669
rect 26200 25666 27000 25696
rect 20621 25664 27000 25666
rect 20621 25608 20626 25664
rect 20682 25608 27000 25664
rect 20621 25606 27000 25608
rect 20621 25603 20687 25606
rect 26200 25576 27000 25606
rect 5022 25468 5028 25532
rect 5092 25530 5098 25532
rect 24209 25530 24275 25533
rect 5092 25528 24275 25530
rect 5092 25472 24214 25528
rect 24270 25472 24275 25528
rect 5092 25470 24275 25472
rect 5092 25468 5098 25470
rect 24209 25467 24275 25470
rect 7782 25332 7788 25396
rect 7852 25394 7858 25396
rect 19425 25394 19491 25397
rect 7852 25392 19491 25394
rect 7852 25336 19430 25392
rect 19486 25336 19491 25392
rect 7852 25334 19491 25336
rect 7852 25332 7858 25334
rect 19425 25331 19491 25334
rect 4838 25196 4844 25260
rect 4908 25258 4914 25260
rect 19374 25258 19380 25260
rect 4908 25198 19380 25258
rect 4908 25196 4914 25198
rect 19374 25196 19380 25198
rect 19444 25196 19450 25260
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 10726 25060 10732 25124
rect 10796 25122 10802 25124
rect 23381 25122 23447 25125
rect 10796 25120 23447 25122
rect 10796 25064 23386 25120
rect 23442 25064 23447 25120
rect 10796 25062 23447 25064
rect 10796 25060 10802 25062
rect 23381 25059 23447 25062
rect 10317 24986 10383 24989
rect 24301 24986 24367 24989
rect 10317 24984 24367 24986
rect 10317 24928 10322 24984
rect 10378 24928 24306 24984
rect 24362 24928 24367 24984
rect 10317 24926 24367 24928
rect 10317 24923 10383 24926
rect 24301 24923 24367 24926
rect 0 24850 800 24880
rect 3601 24850 3667 24853
rect 0 24848 3667 24850
rect 0 24792 3606 24848
rect 3662 24792 3667 24848
rect 0 24790 3667 24792
rect 0 24760 800 24790
rect 3601 24787 3667 24790
rect 13486 24788 13492 24852
rect 13556 24850 13562 24852
rect 24761 24850 24827 24853
rect 26200 24850 27000 24880
rect 13556 24848 24827 24850
rect 13556 24792 24766 24848
rect 24822 24792 24827 24848
rect 13556 24790 24827 24792
rect 13556 24788 13562 24790
rect 24761 24787 24827 24790
rect 24902 24790 27000 24850
rect 9213 24714 9279 24717
rect 17861 24714 17927 24717
rect 9213 24712 17927 24714
rect 9213 24656 9218 24712
rect 9274 24656 17866 24712
rect 17922 24656 17927 24712
rect 9213 24654 17927 24656
rect 9213 24651 9279 24654
rect 17861 24651 17927 24654
rect 22093 24714 22159 24717
rect 24902 24714 24962 24790
rect 26200 24760 27000 24790
rect 22093 24712 24962 24714
rect 22093 24656 22098 24712
rect 22154 24656 24962 24712
rect 22093 24654 24962 24656
rect 22093 24651 22159 24654
rect 15561 24578 15627 24581
rect 18873 24578 18939 24581
rect 15561 24576 18939 24578
rect 15561 24520 15566 24576
rect 15622 24520 18878 24576
rect 18934 24520 18939 24576
rect 15561 24518 18939 24520
rect 15561 24515 15627 24518
rect 18873 24515 18939 24518
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 15193 24442 15259 24445
rect 16389 24442 16455 24445
rect 15193 24440 16455 24442
rect 15193 24384 15198 24440
rect 15254 24384 16394 24440
rect 16450 24384 16455 24440
rect 15193 24382 16455 24384
rect 15193 24379 15259 24382
rect 16389 24379 16455 24382
rect 16941 24442 17007 24445
rect 22737 24442 22803 24445
rect 16941 24440 22803 24442
rect 16941 24384 16946 24440
rect 17002 24384 22742 24440
rect 22798 24384 22803 24440
rect 16941 24382 22803 24384
rect 16941 24379 17007 24382
rect 22737 24379 22803 24382
rect 23381 24442 23447 24445
rect 26200 24442 27000 24472
rect 23381 24440 27000 24442
rect 23381 24384 23386 24440
rect 23442 24384 27000 24440
rect 23381 24382 27000 24384
rect 23381 24379 23447 24382
rect 26200 24352 27000 24382
rect 6269 24306 6335 24309
rect 21265 24306 21331 24309
rect 6269 24304 21331 24306
rect 6269 24248 6274 24304
rect 6330 24248 21270 24304
rect 21326 24248 21331 24304
rect 6269 24246 21331 24248
rect 6269 24243 6335 24246
rect 21265 24243 21331 24246
rect 6729 24172 6795 24173
rect 6678 24108 6684 24172
rect 6748 24170 6795 24172
rect 7005 24170 7071 24173
rect 15193 24170 15259 24173
rect 17953 24170 18019 24173
rect 6748 24168 6840 24170
rect 6790 24112 6840 24168
rect 6748 24110 6840 24112
rect 7005 24168 15259 24170
rect 7005 24112 7010 24168
rect 7066 24112 15198 24168
rect 15254 24112 15259 24168
rect 7005 24110 15259 24112
rect 6748 24108 6795 24110
rect 6729 24107 6795 24108
rect 7005 24107 7071 24110
rect 15193 24107 15259 24110
rect 15334 24168 18019 24170
rect 15334 24112 17958 24168
rect 18014 24112 18019 24168
rect 15334 24110 18019 24112
rect 8518 23972 8524 24036
rect 8588 24034 8594 24036
rect 15334 24034 15394 24110
rect 17953 24107 18019 24110
rect 8588 23974 15394 24034
rect 8588 23972 8594 23974
rect 21398 23972 21404 24036
rect 21468 24034 21474 24036
rect 26200 24034 27000 24064
rect 21468 23974 27000 24034
rect 21468 23972 21474 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 26200 23944 27000 23974
rect 17946 23903 18262 23904
rect 0 23762 800 23792
rect 1485 23762 1551 23765
rect 0 23760 1551 23762
rect 0 23704 1490 23760
rect 1546 23704 1551 23760
rect 0 23702 1551 23704
rect 0 23672 800 23702
rect 1485 23699 1551 23702
rect 1761 23762 1827 23765
rect 20621 23762 20687 23765
rect 1761 23760 20687 23762
rect 1761 23704 1766 23760
rect 1822 23704 20626 23760
rect 20682 23704 20687 23760
rect 1761 23702 20687 23704
rect 1761 23699 1827 23702
rect 20621 23699 20687 23702
rect 9070 23564 9076 23628
rect 9140 23626 9146 23628
rect 24577 23626 24643 23629
rect 9140 23624 24643 23626
rect 9140 23568 24582 23624
rect 24638 23568 24643 23624
rect 9140 23566 24643 23568
rect 9140 23564 9146 23566
rect 24577 23563 24643 23566
rect 24761 23626 24827 23629
rect 26200 23626 27000 23656
rect 24761 23624 27000 23626
rect 24761 23568 24766 23624
rect 24822 23568 27000 23624
rect 24761 23566 27000 23568
rect 24761 23563 24827 23566
rect 26200 23536 27000 23566
rect 6545 23492 6611 23493
rect 6494 23490 6500 23492
rect 6454 23430 6500 23490
rect 6564 23488 6611 23492
rect 6606 23432 6611 23488
rect 6494 23428 6500 23430
rect 6564 23428 6611 23432
rect 7414 23428 7420 23492
rect 7484 23490 7490 23492
rect 9765 23490 9831 23493
rect 7484 23488 9831 23490
rect 7484 23432 9770 23488
rect 9826 23432 9831 23488
rect 7484 23430 9831 23432
rect 7484 23428 7490 23430
rect 6545 23427 6611 23428
rect 9765 23427 9831 23430
rect 12566 23428 12572 23492
rect 12636 23490 12642 23492
rect 12709 23490 12775 23493
rect 12636 23488 12775 23490
rect 12636 23432 12714 23488
rect 12770 23432 12775 23488
rect 12636 23430 12775 23432
rect 12636 23428 12642 23430
rect 12709 23427 12775 23430
rect 16614 23428 16620 23492
rect 16684 23490 16690 23492
rect 17493 23490 17559 23493
rect 16684 23488 17559 23490
rect 16684 23432 17498 23488
rect 17554 23432 17559 23488
rect 16684 23430 17559 23432
rect 16684 23428 16690 23430
rect 17493 23427 17559 23430
rect 18137 23490 18203 23493
rect 19241 23490 19307 23493
rect 18137 23488 19307 23490
rect 18137 23432 18142 23488
rect 18198 23432 19246 23488
rect 19302 23432 19307 23488
rect 18137 23430 19307 23432
rect 18137 23427 18203 23430
rect 19241 23427 19307 23430
rect 19374 23428 19380 23492
rect 19444 23490 19450 23492
rect 19609 23490 19675 23493
rect 19444 23488 19675 23490
rect 19444 23432 19614 23488
rect 19670 23432 19675 23488
rect 19444 23430 19675 23432
rect 19444 23428 19450 23430
rect 19609 23427 19675 23430
rect 19885 23492 19951 23493
rect 19885 23488 19932 23492
rect 19996 23490 20002 23492
rect 20161 23490 20227 23493
rect 20294 23490 20300 23492
rect 19885 23432 19890 23488
rect 19885 23428 19932 23432
rect 19996 23430 20042 23490
rect 20161 23488 20300 23490
rect 20161 23432 20166 23488
rect 20222 23432 20300 23488
rect 20161 23430 20300 23432
rect 19996 23428 20002 23430
rect 19885 23427 19951 23428
rect 20161 23427 20227 23430
rect 20294 23428 20300 23430
rect 20364 23428 20370 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 14089 23354 14155 23357
rect 20805 23354 20871 23357
rect 14089 23352 20871 23354
rect 14089 23296 14094 23352
rect 14150 23296 20810 23352
rect 20866 23296 20871 23352
rect 14089 23294 20871 23296
rect 14089 23291 14155 23294
rect 20805 23291 20871 23294
rect 5441 23218 5507 23221
rect 15929 23218 15995 23221
rect 18137 23218 18203 23221
rect 5441 23216 15995 23218
rect 5441 23160 5446 23216
rect 5502 23160 15934 23216
rect 15990 23160 15995 23216
rect 5441 23158 15995 23160
rect 5441 23155 5507 23158
rect 15929 23155 15995 23158
rect 16070 23216 18203 23218
rect 16070 23160 18142 23216
rect 18198 23160 18203 23216
rect 16070 23158 18203 23160
rect 1853 23082 1919 23085
rect 2129 23082 2195 23085
rect 11053 23082 11119 23085
rect 1853 23080 11119 23082
rect 1853 23024 1858 23080
rect 1914 23024 2134 23080
rect 2190 23024 11058 23080
rect 11114 23024 11119 23080
rect 1853 23022 11119 23024
rect 1853 23019 1919 23022
rect 2129 23019 2195 23022
rect 11053 23019 11119 23022
rect 13629 23082 13695 23085
rect 16070 23082 16130 23158
rect 18137 23155 18203 23158
rect 22134 23156 22140 23220
rect 22204 23218 22210 23220
rect 23381 23218 23447 23221
rect 26200 23218 27000 23248
rect 22204 23216 23447 23218
rect 22204 23160 23386 23216
rect 23442 23160 23447 23216
rect 22204 23158 23447 23160
rect 22204 23156 22210 23158
rect 23381 23155 23447 23158
rect 23614 23158 27000 23218
rect 13629 23080 16130 23082
rect 13629 23024 13634 23080
rect 13690 23024 16130 23080
rect 13629 23022 16130 23024
rect 17309 23082 17375 23085
rect 21725 23082 21791 23085
rect 17309 23080 21791 23082
rect 17309 23024 17314 23080
rect 17370 23024 21730 23080
rect 21786 23024 21791 23080
rect 17309 23022 21791 23024
rect 13629 23019 13695 23022
rect 17309 23019 17375 23022
rect 21725 23019 21791 23022
rect 22461 23082 22527 23085
rect 23614 23082 23674 23158
rect 26200 23128 27000 23158
rect 22461 23080 23674 23082
rect 22461 23024 22466 23080
rect 22522 23024 23674 23080
rect 22461 23022 23674 23024
rect 22461 23019 22527 23022
rect 12341 22946 12407 22949
rect 15653 22946 15719 22949
rect 12341 22944 15719 22946
rect 12341 22888 12346 22944
rect 12402 22888 15658 22944
rect 15714 22888 15719 22944
rect 12341 22886 15719 22888
rect 12341 22883 12407 22886
rect 15653 22883 15719 22886
rect 16205 22946 16271 22949
rect 17677 22946 17743 22949
rect 16205 22944 17743 22946
rect 16205 22888 16210 22944
rect 16266 22888 17682 22944
rect 17738 22888 17743 22944
rect 16205 22886 17743 22888
rect 16205 22883 16271 22886
rect 17677 22883 17743 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 8334 22748 8340 22812
rect 8404 22810 8410 22812
rect 14089 22810 14155 22813
rect 8404 22808 14155 22810
rect 8404 22752 14094 22808
rect 14150 22752 14155 22808
rect 8404 22750 14155 22752
rect 8404 22748 8410 22750
rect 14089 22747 14155 22750
rect 14549 22810 14615 22813
rect 16757 22810 16823 22813
rect 26200 22810 27000 22840
rect 14549 22808 16823 22810
rect 14549 22752 14554 22808
rect 14610 22752 16762 22808
rect 16818 22752 16823 22808
rect 14549 22750 16823 22752
rect 14549 22747 14615 22750
rect 16757 22747 16823 22750
rect 22050 22750 27000 22810
rect 0 22674 800 22704
rect 1669 22674 1735 22677
rect 0 22672 1735 22674
rect 0 22616 1674 22672
rect 1730 22616 1735 22672
rect 0 22614 1735 22616
rect 0 22584 800 22614
rect 1669 22611 1735 22614
rect 9121 22674 9187 22677
rect 21357 22674 21423 22677
rect 9121 22672 21423 22674
rect 9121 22616 9126 22672
rect 9182 22616 21362 22672
rect 21418 22616 21423 22672
rect 9121 22614 21423 22616
rect 9121 22611 9187 22614
rect 21357 22611 21423 22614
rect 5533 22538 5599 22541
rect 14917 22538 14983 22541
rect 5533 22536 14983 22538
rect 5533 22480 5538 22536
rect 5594 22480 14922 22536
rect 14978 22480 14983 22536
rect 5533 22478 14983 22480
rect 5533 22475 5599 22478
rect 14917 22475 14983 22478
rect 16757 22538 16823 22541
rect 19425 22538 19491 22541
rect 19742 22538 19748 22540
rect 16757 22536 19748 22538
rect 16757 22480 16762 22536
rect 16818 22480 19430 22536
rect 19486 22480 19748 22536
rect 16757 22478 19748 22480
rect 16757 22475 16823 22478
rect 19425 22475 19491 22478
rect 19742 22476 19748 22478
rect 19812 22476 19818 22540
rect 9397 22402 9463 22405
rect 11513 22402 11579 22405
rect 9397 22400 11579 22402
rect 9397 22344 9402 22400
rect 9458 22344 11518 22400
rect 11574 22344 11579 22400
rect 9397 22342 11579 22344
rect 9397 22339 9463 22342
rect 11513 22339 11579 22342
rect 14549 22402 14615 22405
rect 15009 22402 15075 22405
rect 14549 22400 15075 22402
rect 14549 22344 14554 22400
rect 14610 22344 15014 22400
rect 15070 22344 15075 22400
rect 14549 22342 15075 22344
rect 14549 22339 14615 22342
rect 15009 22339 15075 22342
rect 16062 22340 16068 22404
rect 16132 22402 16138 22404
rect 22050 22402 22110 22750
rect 26200 22720 27000 22750
rect 16132 22342 22110 22402
rect 23381 22402 23447 22405
rect 26200 22402 27000 22432
rect 23381 22400 27000 22402
rect 23381 22344 23386 22400
rect 23442 22344 27000 22400
rect 23381 22342 27000 22344
rect 16132 22340 16138 22342
rect 23381 22339 23447 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 26200 22312 27000 22342
rect 22946 22271 23262 22272
rect 9765 22266 9831 22269
rect 12709 22266 12775 22269
rect 9765 22264 12775 22266
rect 9765 22208 9770 22264
rect 9826 22208 12714 22264
rect 12770 22208 12775 22264
rect 9765 22206 12775 22208
rect 9765 22203 9831 22206
rect 12709 22203 12775 22206
rect 13854 22204 13860 22268
rect 13924 22266 13930 22268
rect 18321 22266 18387 22269
rect 13924 22264 18387 22266
rect 13924 22208 18326 22264
rect 18382 22208 18387 22264
rect 13924 22206 18387 22208
rect 13924 22204 13930 22206
rect 18321 22203 18387 22206
rect 7238 22070 8402 22130
rect 1761 21994 1827 21997
rect 7238 21994 7298 22070
rect 1761 21992 7298 21994
rect 1761 21936 1766 21992
rect 1822 21936 7298 21992
rect 1761 21934 7298 21936
rect 1761 21931 1827 21934
rect 8342 21858 8402 22070
rect 10174 22068 10180 22132
rect 10244 22130 10250 22132
rect 21265 22130 21331 22133
rect 10244 22070 12266 22130
rect 10244 22068 10250 22070
rect 9397 21994 9463 21997
rect 11881 21994 11947 21997
rect 9397 21992 11947 21994
rect 9397 21936 9402 21992
rect 9458 21936 11886 21992
rect 11942 21936 11947 21992
rect 9397 21934 11947 21936
rect 12206 21994 12266 22070
rect 12942 22128 21331 22130
rect 12942 22072 21270 22128
rect 21326 22072 21331 22128
rect 12942 22070 21331 22072
rect 12942 21994 13002 22070
rect 21265 22067 21331 22070
rect 12206 21934 13002 21994
rect 13813 21994 13879 21997
rect 16757 21994 16823 21997
rect 24945 21994 25011 21997
rect 26200 21994 27000 22024
rect 13813 21992 16823 21994
rect 13813 21936 13818 21992
rect 13874 21936 16762 21992
rect 16818 21936 16823 21992
rect 13813 21934 16823 21936
rect 9397 21931 9463 21934
rect 11881 21931 11947 21934
rect 13813 21931 13879 21934
rect 16757 21931 16823 21934
rect 17174 21934 18476 21994
rect 10041 21858 10107 21861
rect 17174 21858 17234 21934
rect 8342 21856 17234 21858
rect 8342 21800 10046 21856
rect 10102 21800 17234 21856
rect 8342 21798 17234 21800
rect 18416 21858 18476 21934
rect 19750 21992 25011 21994
rect 19750 21936 24950 21992
rect 25006 21936 25011 21992
rect 19750 21934 25011 21936
rect 19750 21858 19810 21934
rect 24945 21931 25011 21934
rect 25086 21934 27000 21994
rect 18416 21798 19810 21858
rect 10041 21795 10107 21798
rect 21766 21796 21772 21860
rect 21836 21858 21842 21860
rect 25086 21858 25146 21934
rect 26200 21904 27000 21934
rect 21836 21798 25146 21858
rect 21836 21796 21842 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 9765 21722 9831 21725
rect 11145 21722 11211 21725
rect 17585 21722 17651 21725
rect 9765 21720 17651 21722
rect 9765 21664 9770 21720
rect 9826 21664 11150 21720
rect 11206 21664 17590 21720
rect 17646 21664 17651 21720
rect 9765 21662 17651 21664
rect 9765 21659 9831 21662
rect 11145 21659 11211 21662
rect 17585 21659 17651 21662
rect 19558 21660 19564 21724
rect 19628 21722 19634 21724
rect 19701 21722 19767 21725
rect 19628 21720 19767 21722
rect 19628 21664 19706 21720
rect 19762 21664 19767 21720
rect 19628 21662 19767 21664
rect 19628 21660 19634 21662
rect 19701 21659 19767 21662
rect 4797 21588 4863 21589
rect 4797 21586 4844 21588
rect 4752 21584 4844 21586
rect 4752 21528 4802 21584
rect 4752 21526 4844 21528
rect 4797 21524 4844 21526
rect 4908 21524 4914 21588
rect 17493 21586 17559 21589
rect 7606 21584 17559 21586
rect 7606 21528 17498 21584
rect 17554 21528 17559 21584
rect 7606 21526 17559 21528
rect 4797 21523 4863 21524
rect 1761 21450 1827 21453
rect 7606 21450 7666 21526
rect 17493 21523 17559 21526
rect 21950 21524 21956 21588
rect 22020 21586 22026 21588
rect 26200 21586 27000 21616
rect 22020 21526 27000 21586
rect 22020 21524 22026 21526
rect 26200 21496 27000 21526
rect 1761 21448 7666 21450
rect 1761 21392 1766 21448
rect 1822 21392 7666 21448
rect 1761 21390 7666 21392
rect 8753 21450 8819 21453
rect 15469 21450 15535 21453
rect 8753 21448 15535 21450
rect 8753 21392 8758 21448
rect 8814 21392 15474 21448
rect 15530 21392 15535 21448
rect 8753 21390 15535 21392
rect 1761 21387 1827 21390
rect 8753 21387 8819 21390
rect 15469 21387 15535 21390
rect 16297 21450 16363 21453
rect 22093 21450 22159 21453
rect 16297 21448 22159 21450
rect 16297 21392 16302 21448
rect 16358 21392 22098 21448
rect 22154 21392 22159 21448
rect 16297 21390 22159 21392
rect 16297 21387 16363 21390
rect 22093 21387 22159 21390
rect 22502 21388 22508 21452
rect 22572 21450 22578 21452
rect 23381 21450 23447 21453
rect 22572 21448 23447 21450
rect 22572 21392 23386 21448
rect 23442 21392 23447 21448
rect 22572 21390 23447 21392
rect 22572 21388 22578 21390
rect 23381 21387 23447 21390
rect 6361 21314 6427 21317
rect 11973 21314 12039 21317
rect 6361 21312 12039 21314
rect 6361 21256 6366 21312
rect 6422 21256 11978 21312
rect 12034 21256 12039 21312
rect 6361 21254 12039 21256
rect 6361 21251 6427 21254
rect 11973 21251 12039 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 14365 21178 14431 21181
rect 18689 21178 18755 21181
rect 14365 21176 18755 21178
rect 14365 21120 14370 21176
rect 14426 21120 18694 21176
rect 18750 21120 18755 21176
rect 14365 21118 18755 21120
rect 14365 21115 14431 21118
rect 18689 21115 18755 21118
rect 24117 21178 24183 21181
rect 24577 21178 24643 21181
rect 24117 21176 24643 21178
rect 24117 21120 24122 21176
rect 24178 21120 24582 21176
rect 24638 21120 24643 21176
rect 24117 21118 24643 21120
rect 24117 21115 24183 21118
rect 24577 21115 24643 21118
rect 26049 21178 26115 21181
rect 26200 21178 27000 21208
rect 26049 21176 27000 21178
rect 26049 21120 26054 21176
rect 26110 21120 27000 21176
rect 26049 21118 27000 21120
rect 26049 21115 26115 21118
rect 26200 21088 27000 21118
rect 8293 21042 8359 21045
rect 13629 21042 13695 21045
rect 8293 21040 13695 21042
rect 8293 20984 8298 21040
rect 8354 20984 13634 21040
rect 13690 20984 13695 21040
rect 8293 20982 13695 20984
rect 8293 20979 8359 20982
rect 13629 20979 13695 20982
rect 15009 21042 15075 21045
rect 15009 21040 24594 21042
rect 15009 20984 15014 21040
rect 15070 20984 24594 21040
rect 15009 20982 24594 20984
rect 15009 20979 15075 20982
rect 7833 20906 7899 20909
rect 11053 20906 11119 20909
rect 7833 20904 11119 20906
rect 7833 20848 7838 20904
rect 7894 20848 11058 20904
rect 11114 20848 11119 20904
rect 7833 20846 11119 20848
rect 7833 20843 7899 20846
rect 11053 20843 11119 20846
rect 11329 20906 11395 20909
rect 24117 20906 24183 20909
rect 11329 20904 24183 20906
rect 11329 20848 11334 20904
rect 11390 20848 24122 20904
rect 24178 20848 24183 20904
rect 11329 20846 24183 20848
rect 11329 20843 11395 20846
rect 24117 20843 24183 20846
rect 11094 20708 11100 20772
rect 11164 20770 11170 20772
rect 12249 20770 12315 20773
rect 11164 20768 12315 20770
rect 11164 20712 12254 20768
rect 12310 20712 12315 20768
rect 11164 20710 12315 20712
rect 11164 20708 11170 20710
rect 12249 20707 12315 20710
rect 15837 20772 15903 20773
rect 15837 20768 15884 20772
rect 15948 20770 15954 20772
rect 16481 20770 16547 20773
rect 15837 20712 15842 20768
rect 15837 20708 15884 20712
rect 15948 20710 15994 20770
rect 16438 20768 16547 20770
rect 16438 20712 16486 20768
rect 16542 20712 16547 20768
rect 15948 20708 15954 20710
rect 15837 20707 15903 20708
rect 16438 20707 16547 20712
rect 24534 20770 24594 20982
rect 26200 20770 27000 20800
rect 24534 20710 27000 20770
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 9397 20634 9463 20637
rect 12433 20634 12499 20637
rect 9397 20632 12499 20634
rect 9397 20576 9402 20632
rect 9458 20576 12438 20632
rect 12494 20576 12499 20632
rect 9397 20574 12499 20576
rect 16438 20634 16498 20707
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 26200 20680 27000 20710
rect 17946 20639 18262 20640
rect 17401 20634 17467 20637
rect 16438 20632 17467 20634
rect 16438 20576 17406 20632
rect 17462 20576 17467 20632
rect 16438 20574 17467 20576
rect 9397 20571 9463 20574
rect 12433 20571 12499 20574
rect 17401 20571 17467 20574
rect 19977 20634 20043 20637
rect 24669 20634 24735 20637
rect 19977 20632 24735 20634
rect 19977 20576 19982 20632
rect 20038 20576 24674 20632
rect 24730 20576 24735 20632
rect 19977 20574 24735 20576
rect 19977 20571 20043 20574
rect 24669 20571 24735 20574
rect 11329 20498 11395 20501
rect 2730 20496 11395 20498
rect 2730 20440 11334 20496
rect 11390 20440 11395 20496
rect 2730 20438 11395 20440
rect 2589 20362 2655 20365
rect 2730 20362 2790 20438
rect 11329 20435 11395 20438
rect 11513 20498 11579 20501
rect 15285 20498 15351 20501
rect 11513 20496 15351 20498
rect 11513 20440 11518 20496
rect 11574 20440 15290 20496
rect 15346 20440 15351 20496
rect 11513 20438 15351 20440
rect 11513 20435 11579 20438
rect 15285 20435 15351 20438
rect 2589 20360 2790 20362
rect 2589 20304 2594 20360
rect 2650 20304 2790 20360
rect 2589 20302 2790 20304
rect 6821 20362 6887 20365
rect 16205 20362 16271 20365
rect 6821 20360 16271 20362
rect 6821 20304 6826 20360
rect 6882 20304 16210 20360
rect 16266 20304 16271 20360
rect 6821 20302 16271 20304
rect 2589 20299 2655 20302
rect 6821 20299 6887 20302
rect 16205 20299 16271 20302
rect 17166 20300 17172 20364
rect 17236 20362 17242 20364
rect 19517 20362 19583 20365
rect 17236 20360 19583 20362
rect 17236 20304 19522 20360
rect 19578 20304 19583 20360
rect 17236 20302 19583 20304
rect 17236 20300 17242 20302
rect 19517 20299 19583 20302
rect 22277 20362 22343 20365
rect 26200 20362 27000 20392
rect 22277 20360 27000 20362
rect 22277 20304 22282 20360
rect 22338 20304 27000 20360
rect 22277 20302 27000 20304
rect 22277 20299 22343 20302
rect 26200 20272 27000 20302
rect 3601 20226 3667 20229
rect 10869 20226 10935 20229
rect 3601 20224 10935 20226
rect 3601 20168 3606 20224
rect 3662 20168 10874 20224
rect 10930 20168 10935 20224
rect 3601 20166 10935 20168
rect 3601 20163 3667 20166
rect 10869 20163 10935 20166
rect 13537 20226 13603 20229
rect 13813 20226 13879 20229
rect 14181 20226 14247 20229
rect 16665 20226 16731 20229
rect 13537 20224 16731 20226
rect 13537 20168 13542 20224
rect 13598 20168 13818 20224
rect 13874 20168 14186 20224
rect 14242 20168 16670 20224
rect 16726 20168 16731 20224
rect 13537 20166 16731 20168
rect 13537 20163 13603 20166
rect 13813 20163 13879 20166
rect 14181 20163 14247 20166
rect 16665 20163 16731 20166
rect 16849 20226 16915 20229
rect 18454 20226 18460 20228
rect 16849 20224 18460 20226
rect 16849 20168 16854 20224
rect 16910 20168 18460 20224
rect 16849 20166 18460 20168
rect 16849 20163 16915 20166
rect 18454 20164 18460 20166
rect 18524 20164 18530 20228
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 7281 20090 7347 20093
rect 7782 20090 7788 20092
rect 7281 20088 7788 20090
rect 7281 20032 7286 20088
rect 7342 20032 7788 20088
rect 7281 20030 7788 20032
rect 7281 20027 7347 20030
rect 7782 20028 7788 20030
rect 7852 20028 7858 20092
rect 22553 20090 22619 20093
rect 17174 20088 22619 20090
rect 17174 20032 22558 20088
rect 22614 20032 22619 20088
rect 17174 20030 22619 20032
rect 5349 19954 5415 19957
rect 10777 19954 10843 19957
rect 17174 19954 17234 20030
rect 22553 20027 22619 20030
rect 5349 19952 10610 19954
rect 5349 19896 5354 19952
rect 5410 19896 10610 19952
rect 5349 19894 10610 19896
rect 5349 19891 5415 19894
rect 7189 19818 7255 19821
rect 10409 19818 10475 19821
rect 7189 19816 10475 19818
rect 7189 19760 7194 19816
rect 7250 19760 10414 19816
rect 10470 19760 10475 19816
rect 7189 19758 10475 19760
rect 7189 19755 7255 19758
rect 10409 19755 10475 19758
rect 10550 19682 10610 19894
rect 10777 19952 17234 19954
rect 10777 19896 10782 19952
rect 10838 19896 17234 19952
rect 10777 19894 17234 19896
rect 17401 19954 17467 19957
rect 25037 19954 25103 19957
rect 26200 19954 27000 19984
rect 17401 19952 25103 19954
rect 17401 19896 17406 19952
rect 17462 19896 25042 19952
rect 25098 19896 25103 19952
rect 17401 19894 25103 19896
rect 10777 19891 10843 19894
rect 17401 19891 17467 19894
rect 25037 19891 25103 19894
rect 25270 19894 27000 19954
rect 10869 19818 10935 19821
rect 16757 19818 16823 19821
rect 19333 19818 19399 19821
rect 10869 19816 16823 19818
rect 10869 19760 10874 19816
rect 10930 19760 16762 19816
rect 16818 19760 16823 19816
rect 10869 19758 16823 19760
rect 10869 19755 10935 19758
rect 16757 19755 16823 19758
rect 17174 19816 19399 19818
rect 17174 19760 19338 19816
rect 19394 19760 19399 19816
rect 17174 19758 19399 19760
rect 13537 19682 13603 19685
rect 10550 19680 13603 19682
rect 10550 19624 13542 19680
rect 13598 19624 13603 19680
rect 10550 19622 13603 19624
rect 13537 19619 13603 19622
rect 13721 19682 13787 19685
rect 17174 19682 17234 19758
rect 19333 19755 19399 19758
rect 19517 19818 19583 19821
rect 23381 19818 23447 19821
rect 19517 19816 23447 19818
rect 19517 19760 19522 19816
rect 19578 19760 23386 19816
rect 23442 19760 23447 19816
rect 19517 19758 23447 19760
rect 19517 19755 19583 19758
rect 23381 19755 23447 19758
rect 13721 19680 17234 19682
rect 13721 19624 13726 19680
rect 13782 19624 17234 19680
rect 13721 19622 17234 19624
rect 20621 19682 20687 19685
rect 25270 19682 25330 19894
rect 26200 19864 27000 19894
rect 20621 19680 25330 19682
rect 20621 19624 20626 19680
rect 20682 19624 25330 19680
rect 20621 19622 25330 19624
rect 13721 19619 13787 19622
rect 20621 19619 20687 19622
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 7281 19548 7347 19549
rect 7230 19484 7236 19548
rect 7300 19546 7347 19548
rect 8385 19546 8451 19549
rect 15285 19546 15351 19549
rect 7300 19544 7392 19546
rect 7342 19488 7392 19544
rect 7300 19486 7392 19488
rect 8385 19544 15351 19546
rect 8385 19488 8390 19544
rect 8446 19488 15290 19544
rect 15346 19488 15351 19544
rect 8385 19486 15351 19488
rect 7300 19484 7347 19486
rect 7281 19483 7347 19484
rect 8385 19483 8451 19486
rect 15285 19483 15351 19486
rect 23749 19546 23815 19549
rect 26200 19546 27000 19576
rect 23749 19544 27000 19546
rect 23749 19488 23754 19544
rect 23810 19488 27000 19544
rect 23749 19486 27000 19488
rect 23749 19483 23815 19486
rect 26200 19456 27000 19486
rect 7005 19410 7071 19413
rect 8334 19410 8340 19412
rect 7005 19408 8340 19410
rect 7005 19352 7010 19408
rect 7066 19352 8340 19408
rect 7005 19350 8340 19352
rect 7005 19347 7071 19350
rect 8334 19348 8340 19350
rect 8404 19348 8410 19412
rect 13537 19410 13603 19413
rect 17401 19410 17467 19413
rect 13537 19408 17467 19410
rect 13537 19352 13542 19408
rect 13598 19352 17406 19408
rect 17462 19352 17467 19408
rect 13537 19350 17467 19352
rect 13537 19347 13603 19350
rect 17401 19347 17467 19350
rect 17534 19348 17540 19412
rect 17604 19410 17610 19412
rect 17769 19410 17835 19413
rect 17604 19408 17835 19410
rect 17604 19352 17774 19408
rect 17830 19352 17835 19408
rect 17604 19350 17835 19352
rect 17604 19348 17610 19350
rect 17769 19347 17835 19350
rect 19517 19410 19583 19413
rect 20110 19410 20116 19412
rect 19517 19408 20116 19410
rect 19517 19352 19522 19408
rect 19578 19352 20116 19408
rect 19517 19350 20116 19352
rect 19517 19347 19583 19350
rect 20110 19348 20116 19350
rect 20180 19348 20186 19412
rect 20713 19410 20779 19413
rect 22001 19410 22067 19413
rect 22185 19410 22251 19413
rect 20713 19408 22251 19410
rect 20713 19352 20718 19408
rect 20774 19352 22006 19408
rect 22062 19352 22190 19408
rect 22246 19352 22251 19408
rect 20713 19350 22251 19352
rect 20713 19347 20779 19350
rect 22001 19347 22067 19350
rect 22185 19347 22251 19350
rect 5625 19274 5691 19277
rect 21265 19274 21331 19277
rect 5625 19272 21331 19274
rect 5625 19216 5630 19272
rect 5686 19216 21270 19272
rect 21326 19216 21331 19272
rect 5625 19214 21331 19216
rect 5625 19211 5691 19214
rect 21265 19211 21331 19214
rect 14641 19138 14707 19141
rect 19057 19138 19123 19141
rect 14641 19136 19123 19138
rect 14641 19080 14646 19136
rect 14702 19080 19062 19136
rect 19118 19080 19123 19136
rect 14641 19078 19123 19080
rect 14641 19075 14707 19078
rect 19057 19075 19123 19078
rect 23381 19138 23447 19141
rect 26200 19138 27000 19168
rect 23381 19136 27000 19138
rect 23381 19080 23386 19136
rect 23442 19080 27000 19136
rect 23381 19078 27000 19080
rect 23381 19075 23447 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 26200 19048 27000 19078
rect 22946 19007 23262 19008
rect 3509 19002 3575 19005
rect 11421 19002 11487 19005
rect 3509 19000 11487 19002
rect 3509 18944 3514 19000
rect 3570 18944 11426 19000
rect 11482 18944 11487 19000
rect 3509 18942 11487 18944
rect 3509 18939 3575 18942
rect 11421 18939 11487 18942
rect 13353 19002 13419 19005
rect 13353 19000 22110 19002
rect 13353 18944 13358 19000
rect 13414 18944 22110 19000
rect 13353 18942 22110 18944
rect 13353 18939 13419 18942
rect 4981 18866 5047 18869
rect 9029 18866 9095 18869
rect 10225 18866 10291 18869
rect 4981 18864 10291 18866
rect 4981 18808 4986 18864
rect 5042 18808 9034 18864
rect 9090 18808 10230 18864
rect 10286 18808 10291 18864
rect 4981 18806 10291 18808
rect 4981 18803 5047 18806
rect 9029 18803 9095 18806
rect 10225 18803 10291 18806
rect 11053 18866 11119 18869
rect 16757 18866 16823 18869
rect 11053 18864 16823 18866
rect 11053 18808 11058 18864
rect 11114 18808 16762 18864
rect 16818 18808 16823 18864
rect 11053 18806 16823 18808
rect 22050 18866 22110 18942
rect 22318 18940 22324 19004
rect 22388 19002 22394 19004
rect 22461 19002 22527 19005
rect 22388 19000 22527 19002
rect 22388 18944 22466 19000
rect 22522 18944 22527 19000
rect 22388 18942 22527 18944
rect 22388 18940 22394 18942
rect 22461 18939 22527 18942
rect 23657 18866 23723 18869
rect 22050 18864 23723 18866
rect 22050 18808 23662 18864
rect 23718 18808 23723 18864
rect 22050 18806 23723 18808
rect 11053 18803 11119 18806
rect 16757 18803 16823 18806
rect 23657 18803 23723 18806
rect 5809 18730 5875 18733
rect 20897 18730 20963 18733
rect 5809 18728 20963 18730
rect 5809 18672 5814 18728
rect 5870 18672 20902 18728
rect 20958 18672 20963 18728
rect 5809 18670 20963 18672
rect 5809 18667 5875 18670
rect 20897 18667 20963 18670
rect 23381 18730 23447 18733
rect 26200 18730 27000 18760
rect 23381 18728 27000 18730
rect 23381 18672 23386 18728
rect 23442 18672 27000 18728
rect 23381 18670 27000 18672
rect 23381 18667 23447 18670
rect 26200 18640 27000 18670
rect 11605 18594 11671 18597
rect 15009 18594 15075 18597
rect 11605 18592 15075 18594
rect 11605 18536 11610 18592
rect 11666 18536 15014 18592
rect 15070 18536 15075 18592
rect 11605 18534 15075 18536
rect 11605 18531 11671 18534
rect 15009 18531 15075 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 9949 18458 10015 18461
rect 16481 18458 16547 18461
rect 9949 18456 16547 18458
rect 9949 18400 9954 18456
rect 10010 18400 16486 18456
rect 16542 18400 16547 18456
rect 9949 18398 16547 18400
rect 9949 18395 10015 18398
rect 16481 18395 16547 18398
rect 4061 18324 4127 18325
rect 4061 18322 4108 18324
rect 4016 18320 4108 18322
rect 4016 18264 4066 18320
rect 4016 18262 4108 18264
rect 4061 18260 4108 18262
rect 4172 18260 4178 18324
rect 9305 18322 9371 18325
rect 13854 18322 13860 18324
rect 9305 18320 13860 18322
rect 9305 18264 9310 18320
rect 9366 18264 13860 18320
rect 9305 18262 13860 18264
rect 4061 18259 4127 18260
rect 9305 18259 9371 18262
rect 13854 18260 13860 18262
rect 13924 18260 13930 18324
rect 14549 18322 14615 18325
rect 19701 18322 19767 18325
rect 14549 18320 19767 18322
rect 14549 18264 14554 18320
rect 14610 18264 19706 18320
rect 19762 18264 19767 18320
rect 14549 18262 19767 18264
rect 14549 18259 14615 18262
rect 19701 18259 19767 18262
rect 23381 18322 23447 18325
rect 26200 18322 27000 18352
rect 23381 18320 27000 18322
rect 23381 18264 23386 18320
rect 23442 18264 27000 18320
rect 23381 18262 27000 18264
rect 23381 18259 23447 18262
rect 26200 18232 27000 18262
rect 7649 18186 7715 18189
rect 23197 18186 23263 18189
rect 7649 18184 23263 18186
rect 7649 18128 7654 18184
rect 7710 18128 23202 18184
rect 23258 18128 23263 18184
rect 7649 18126 23263 18128
rect 7649 18123 7715 18126
rect 23197 18123 23263 18126
rect 4981 18050 5047 18053
rect 7414 18050 7420 18052
rect 4981 18048 7420 18050
rect 4981 17992 4986 18048
rect 5042 17992 7420 18048
rect 4981 17990 7420 17992
rect 4981 17987 5047 17990
rect 7414 17988 7420 17990
rect 7484 17988 7490 18052
rect 12525 18050 12591 18053
rect 7606 18048 12591 18050
rect 7606 17992 12530 18048
rect 12586 17992 12591 18048
rect 7606 17990 12591 17992
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 7606 17914 7666 17990
rect 12525 17987 12591 17990
rect 17677 18052 17743 18053
rect 17677 18048 17724 18052
rect 17788 18050 17794 18052
rect 24577 18050 24643 18053
rect 24710 18050 24716 18052
rect 17677 17992 17682 18048
rect 17677 17988 17724 17992
rect 17788 17990 17834 18050
rect 24577 18048 24716 18050
rect 24577 17992 24582 18048
rect 24638 17992 24716 18048
rect 24577 17990 24716 17992
rect 17788 17988 17794 17990
rect 17677 17987 17743 17988
rect 24577 17987 24643 17990
rect 24710 17988 24716 17990
rect 24780 17988 24786 18052
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 4662 17854 7666 17914
rect 7833 17914 7899 17917
rect 12617 17914 12683 17917
rect 7833 17912 12683 17914
rect 7833 17856 7838 17912
rect 7894 17856 12622 17912
rect 12678 17856 12683 17912
rect 7833 17854 12683 17856
rect 1945 17778 2011 17781
rect 4662 17778 4722 17854
rect 7833 17851 7899 17854
rect 12617 17851 12683 17854
rect 14457 17914 14523 17917
rect 20713 17914 20779 17917
rect 26200 17914 27000 17944
rect 14457 17912 20779 17914
rect 14457 17856 14462 17912
rect 14518 17856 20718 17912
rect 20774 17856 20779 17912
rect 14457 17854 20779 17856
rect 14457 17851 14523 17854
rect 20713 17851 20779 17854
rect 23384 17854 27000 17914
rect 1945 17776 4722 17778
rect 1945 17720 1950 17776
rect 2006 17720 4722 17776
rect 1945 17718 4722 17720
rect 4797 17778 4863 17781
rect 5022 17778 5028 17780
rect 4797 17776 5028 17778
rect 4797 17720 4802 17776
rect 4858 17720 5028 17776
rect 4797 17718 5028 17720
rect 1945 17715 2011 17718
rect 4797 17715 4863 17718
rect 5022 17716 5028 17718
rect 5092 17716 5098 17780
rect 7281 17778 7347 17781
rect 7465 17778 7531 17781
rect 7281 17776 7531 17778
rect 7281 17720 7286 17776
rect 7342 17720 7470 17776
rect 7526 17720 7531 17776
rect 7281 17718 7531 17720
rect 7281 17715 7347 17718
rect 7465 17715 7531 17718
rect 8293 17778 8359 17781
rect 22921 17778 22987 17781
rect 8293 17776 22987 17778
rect 8293 17720 8298 17776
rect 8354 17720 22926 17776
rect 22982 17720 22987 17776
rect 8293 17718 22987 17720
rect 8293 17715 8359 17718
rect 22921 17715 22987 17718
rect 23197 17778 23263 17781
rect 23384 17778 23444 17854
rect 26200 17824 27000 17854
rect 23197 17776 23444 17778
rect 23197 17720 23202 17776
rect 23258 17720 23444 17776
rect 23197 17718 23444 17720
rect 23197 17715 23263 17718
rect 3233 17642 3299 17645
rect 24025 17642 24091 17645
rect 3233 17640 24091 17642
rect 3233 17584 3238 17640
rect 3294 17584 24030 17640
rect 24086 17584 24091 17640
rect 3233 17582 24091 17584
rect 3233 17579 3299 17582
rect 24025 17579 24091 17582
rect 12433 17506 12499 17509
rect 26200 17506 27000 17536
rect 12433 17504 17418 17506
rect 12433 17448 12438 17504
rect 12494 17448 17418 17504
rect 12433 17446 17418 17448
rect 12433 17443 12499 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 8753 17370 8819 17373
rect 17217 17370 17283 17373
rect 8753 17368 17283 17370
rect 8753 17312 8758 17368
rect 8814 17312 17222 17368
rect 17278 17312 17283 17368
rect 8753 17310 17283 17312
rect 8753 17307 8819 17310
rect 17217 17307 17283 17310
rect 2129 17234 2195 17237
rect 12382 17234 12388 17236
rect 2129 17232 12388 17234
rect 2129 17176 2134 17232
rect 2190 17176 12388 17232
rect 2129 17174 12388 17176
rect 2129 17171 2195 17174
rect 12382 17172 12388 17174
rect 12452 17172 12458 17236
rect 15009 17234 15075 17237
rect 15653 17234 15719 17237
rect 16205 17234 16271 17237
rect 15009 17232 16271 17234
rect 15009 17176 15014 17232
rect 15070 17176 15658 17232
rect 15714 17176 16210 17232
rect 16266 17176 16271 17232
rect 15009 17174 16271 17176
rect 17358 17234 17418 17446
rect 22050 17446 27000 17506
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 18689 17234 18755 17237
rect 17358 17232 18755 17234
rect 17358 17176 18694 17232
rect 18750 17176 18755 17232
rect 17358 17174 18755 17176
rect 15009 17171 15075 17174
rect 15653 17171 15719 17174
rect 16205 17171 16271 17174
rect 18689 17171 18755 17174
rect 2773 17098 2839 17101
rect 11094 17098 11100 17100
rect 2773 17096 11100 17098
rect 2773 17040 2778 17096
rect 2834 17040 11100 17096
rect 2773 17038 11100 17040
rect 2773 17035 2839 17038
rect 11094 17036 11100 17038
rect 11164 17036 11170 17100
rect 11329 17098 11395 17101
rect 22050 17098 22110 17446
rect 26200 17416 27000 17446
rect 11329 17096 22110 17098
rect 11329 17040 11334 17096
rect 11390 17040 22110 17096
rect 11329 17038 22110 17040
rect 11329 17035 11395 17038
rect 22686 17036 22692 17100
rect 22756 17098 22762 17100
rect 23197 17098 23263 17101
rect 22756 17096 23263 17098
rect 22756 17040 23202 17096
rect 23258 17040 23263 17096
rect 22756 17038 23263 17040
rect 22756 17036 22762 17038
rect 23197 17035 23263 17038
rect 24669 17098 24735 17101
rect 26200 17098 27000 17128
rect 24669 17096 27000 17098
rect 24669 17040 24674 17096
rect 24730 17040 27000 17096
rect 24669 17038 27000 17040
rect 24669 17035 24735 17038
rect 26200 17008 27000 17038
rect 7281 16962 7347 16965
rect 8753 16962 8819 16965
rect 7281 16960 8819 16962
rect 7281 16904 7286 16960
rect 7342 16904 8758 16960
rect 8814 16904 8819 16960
rect 7281 16902 8819 16904
rect 7281 16899 7347 16902
rect 8753 16899 8819 16902
rect 19374 16900 19380 16964
rect 19444 16962 19450 16964
rect 19517 16962 19583 16965
rect 19444 16960 19583 16962
rect 19444 16904 19522 16960
rect 19578 16904 19583 16960
rect 19444 16902 19583 16904
rect 19444 16900 19450 16902
rect 19517 16899 19583 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 4245 16826 4311 16829
rect 5717 16826 5783 16829
rect 4245 16824 5783 16826
rect 4245 16768 4250 16824
rect 4306 16768 5722 16824
rect 5778 16768 5783 16824
rect 4245 16766 5783 16768
rect 4245 16763 4311 16766
rect 5717 16763 5783 16766
rect 6913 16826 6979 16829
rect 9029 16828 9095 16829
rect 8518 16826 8524 16828
rect 6913 16824 8524 16826
rect 6913 16768 6918 16824
rect 6974 16768 8524 16824
rect 6913 16766 8524 16768
rect 6913 16763 6979 16766
rect 8518 16764 8524 16766
rect 8588 16764 8594 16828
rect 9029 16826 9076 16828
rect 8984 16824 9076 16826
rect 8984 16768 9034 16824
rect 8984 16766 9076 16768
rect 9029 16764 9076 16766
rect 9140 16764 9146 16828
rect 10041 16826 10107 16829
rect 10174 16826 10180 16828
rect 10041 16824 10180 16826
rect 10041 16768 10046 16824
rect 10102 16768 10180 16824
rect 10041 16766 10180 16768
rect 9029 16763 9095 16764
rect 10041 16763 10107 16766
rect 10174 16764 10180 16766
rect 10244 16764 10250 16828
rect 17125 16826 17191 16829
rect 14966 16824 17191 16826
rect 14966 16768 17130 16824
rect 17186 16768 17191 16824
rect 14966 16766 17191 16768
rect 3877 16690 3943 16693
rect 14966 16690 15026 16766
rect 17125 16763 17191 16766
rect 3877 16688 15026 16690
rect 3877 16632 3882 16688
rect 3938 16632 15026 16688
rect 3877 16630 15026 16632
rect 23381 16690 23447 16693
rect 26200 16690 27000 16720
rect 23381 16688 27000 16690
rect 23381 16632 23386 16688
rect 23442 16632 27000 16688
rect 23381 16630 27000 16632
rect 3877 16627 3943 16630
rect 23381 16627 23447 16630
rect 26200 16600 27000 16630
rect 8293 16554 8359 16557
rect 9489 16554 9555 16557
rect 18781 16554 18847 16557
rect 8293 16552 8770 16554
rect 8293 16496 8298 16552
rect 8354 16496 8770 16552
rect 8293 16494 8770 16496
rect 8293 16491 8359 16494
rect 8710 16418 8770 16494
rect 9489 16552 18847 16554
rect 9489 16496 9494 16552
rect 9550 16496 18786 16552
rect 18842 16496 18847 16552
rect 9489 16494 18847 16496
rect 9489 16491 9555 16494
rect 18781 16491 18847 16494
rect 15837 16418 15903 16421
rect 8710 16416 15903 16418
rect 8710 16360 15842 16416
rect 15898 16360 15903 16416
rect 8710 16358 15903 16360
rect 15837 16355 15903 16358
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 14181 16282 14247 16285
rect 12390 16280 14247 16282
rect 12390 16224 14186 16280
rect 14242 16224 14247 16280
rect 12390 16222 14247 16224
rect 2129 16146 2195 16149
rect 2262 16146 2268 16148
rect 2129 16144 2268 16146
rect 2129 16088 2134 16144
rect 2190 16088 2268 16144
rect 2129 16086 2268 16088
rect 2129 16083 2195 16086
rect 2262 16084 2268 16086
rect 2332 16084 2338 16148
rect 8017 16146 8083 16149
rect 12390 16146 12450 16222
rect 14181 16219 14247 16222
rect 24853 16282 24919 16285
rect 25681 16282 25747 16285
rect 26200 16282 27000 16312
rect 24853 16280 27000 16282
rect 24853 16224 24858 16280
rect 24914 16224 25686 16280
rect 25742 16224 27000 16280
rect 24853 16222 27000 16224
rect 24853 16219 24919 16222
rect 25681 16219 25747 16222
rect 26200 16192 27000 16222
rect 8017 16144 12450 16146
rect 8017 16088 8022 16144
rect 8078 16088 12450 16144
rect 8017 16086 12450 16088
rect 8017 16083 8083 16086
rect 7281 16012 7347 16013
rect 7230 16010 7236 16012
rect 7190 15950 7236 16010
rect 7300 16008 7347 16012
rect 7342 15952 7347 16008
rect 7230 15948 7236 15950
rect 7300 15948 7347 15952
rect 7281 15947 7347 15948
rect 7833 16010 7899 16013
rect 20989 16010 21055 16013
rect 7833 16008 21055 16010
rect 7833 15952 7838 16008
rect 7894 15952 20994 16008
rect 21050 15952 21055 16008
rect 7833 15950 21055 15952
rect 7833 15947 7899 15950
rect 20989 15947 21055 15950
rect 8293 15874 8359 15877
rect 12341 15874 12407 15877
rect 8293 15872 12407 15874
rect 8293 15816 8298 15872
rect 8354 15816 12346 15872
rect 12402 15816 12407 15872
rect 8293 15814 12407 15816
rect 8293 15811 8359 15814
rect 12341 15811 12407 15814
rect 15745 15874 15811 15877
rect 22318 15874 22324 15876
rect 15745 15872 22324 15874
rect 15745 15816 15750 15872
rect 15806 15816 22324 15872
rect 15745 15814 22324 15816
rect 15745 15811 15811 15814
rect 22318 15812 22324 15814
rect 22388 15812 22394 15876
rect 25405 15874 25471 15877
rect 26200 15874 27000 15904
rect 25405 15872 27000 15874
rect 25405 15816 25410 15872
rect 25466 15816 27000 15872
rect 25405 15814 27000 15816
rect 25405 15811 25471 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 26200 15784 27000 15814
rect 22946 15743 23262 15744
rect 11513 15738 11579 15741
rect 11881 15738 11947 15741
rect 11513 15736 11947 15738
rect 11513 15680 11518 15736
rect 11574 15680 11886 15736
rect 11942 15680 11947 15736
rect 11513 15678 11947 15680
rect 11513 15675 11579 15678
rect 11881 15675 11947 15678
rect 14273 15738 14339 15741
rect 14641 15738 14707 15741
rect 19374 15738 19380 15740
rect 14273 15736 14707 15738
rect 14273 15680 14278 15736
rect 14334 15680 14646 15736
rect 14702 15680 14707 15736
rect 14273 15678 14707 15680
rect 14273 15675 14339 15678
rect 14641 15675 14707 15678
rect 16024 15678 19380 15738
rect 5257 15602 5323 15605
rect 11421 15602 11487 15605
rect 5257 15600 11487 15602
rect 5257 15544 5262 15600
rect 5318 15544 11426 15600
rect 11482 15544 11487 15600
rect 5257 15542 11487 15544
rect 5257 15539 5323 15542
rect 11421 15539 11487 15542
rect 4705 15466 4771 15469
rect 14457 15466 14523 15469
rect 4705 15464 14523 15466
rect 4705 15408 4710 15464
rect 4766 15408 14462 15464
rect 14518 15408 14523 15464
rect 4705 15406 14523 15408
rect 4705 15403 4771 15406
rect 14457 15403 14523 15406
rect 10777 15330 10843 15333
rect 13353 15330 13419 15333
rect 10777 15328 13419 15330
rect 10777 15272 10782 15328
rect 10838 15272 13358 15328
rect 13414 15272 13419 15328
rect 10777 15270 13419 15272
rect 10777 15267 10843 15270
rect 13353 15267 13419 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 10961 15194 11027 15197
rect 16024 15194 16084 15678
rect 19374 15676 19380 15678
rect 19444 15676 19450 15740
rect 16205 15602 16271 15605
rect 25221 15602 25287 15605
rect 16205 15600 25287 15602
rect 16205 15544 16210 15600
rect 16266 15544 25226 15600
rect 25282 15544 25287 15600
rect 16205 15542 25287 15544
rect 16205 15539 16271 15542
rect 25221 15539 25287 15542
rect 17585 15466 17651 15469
rect 21633 15466 21699 15469
rect 26200 15466 27000 15496
rect 17585 15464 18522 15466
rect 17585 15408 17590 15464
rect 17646 15408 18522 15464
rect 17585 15406 18522 15408
rect 17585 15403 17651 15406
rect 18462 15330 18522 15406
rect 21633 15464 27000 15466
rect 21633 15408 21638 15464
rect 21694 15408 27000 15464
rect 21633 15406 27000 15408
rect 21633 15403 21699 15406
rect 26200 15376 27000 15406
rect 23749 15330 23815 15333
rect 18462 15328 23815 15330
rect 18462 15272 23754 15328
rect 23810 15272 23815 15328
rect 18462 15270 23815 15272
rect 23749 15267 23815 15270
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 25129 15194 25195 15197
rect 10961 15192 16084 15194
rect 10961 15136 10966 15192
rect 11022 15136 16084 15192
rect 10961 15134 16084 15136
rect 22050 15192 25195 15194
rect 22050 15136 25134 15192
rect 25190 15136 25195 15192
rect 22050 15134 25195 15136
rect 10961 15131 11027 15134
rect 10501 15058 10567 15061
rect 10726 15058 10732 15060
rect 10501 15056 10732 15058
rect 10501 15000 10506 15056
rect 10562 15000 10732 15056
rect 10501 14998 10732 15000
rect 10501 14995 10567 14998
rect 10726 14996 10732 14998
rect 10796 14996 10802 15060
rect 22050 15058 22110 15134
rect 25129 15131 25195 15134
rect 26200 15058 27000 15088
rect 12390 14998 22110 15058
rect 24166 14998 27000 15058
rect 3877 14922 3943 14925
rect 12390 14922 12450 14998
rect 3877 14920 12450 14922
rect 3877 14864 3882 14920
rect 3938 14864 12450 14920
rect 3877 14862 12450 14864
rect 17217 14922 17283 14925
rect 24166 14922 24226 14998
rect 26200 14968 27000 14998
rect 17217 14920 24226 14922
rect 17217 14864 17222 14920
rect 17278 14864 24226 14920
rect 17217 14862 24226 14864
rect 3877 14859 3943 14862
rect 17217 14859 17283 14862
rect 11881 14786 11947 14789
rect 12617 14786 12683 14789
rect 11881 14784 12683 14786
rect 11881 14728 11886 14784
rect 11942 14728 12622 14784
rect 12678 14728 12683 14784
rect 11881 14726 12683 14728
rect 11881 14723 11947 14726
rect 12617 14723 12683 14726
rect 13905 14786 13971 14789
rect 22686 14786 22692 14788
rect 13905 14784 22692 14786
rect 13905 14728 13910 14784
rect 13966 14728 22692 14784
rect 13905 14726 22692 14728
rect 13905 14723 13971 14726
rect 22686 14724 22692 14726
rect 22756 14724 22762 14788
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 13813 14650 13879 14653
rect 20161 14650 20227 14653
rect 13813 14648 20227 14650
rect 13813 14592 13818 14648
rect 13874 14592 20166 14648
rect 20222 14592 20227 14648
rect 13813 14590 20227 14592
rect 13813 14587 13879 14590
rect 20161 14587 20227 14590
rect 24853 14650 24919 14653
rect 26200 14650 27000 14680
rect 24853 14648 27000 14650
rect 24853 14592 24858 14648
rect 24914 14592 27000 14648
rect 24853 14590 27000 14592
rect 24853 14587 24919 14590
rect 26200 14560 27000 14590
rect 5901 14514 5967 14517
rect 16614 14514 16620 14516
rect 5901 14512 16620 14514
rect 5901 14456 5906 14512
rect 5962 14456 16620 14512
rect 5901 14454 16620 14456
rect 5901 14451 5967 14454
rect 16614 14452 16620 14454
rect 16684 14452 16690 14516
rect 16757 14514 16823 14517
rect 20294 14514 20300 14516
rect 16757 14512 20300 14514
rect 16757 14456 16762 14512
rect 16818 14456 20300 14512
rect 16757 14454 20300 14456
rect 16757 14451 16823 14454
rect 20294 14452 20300 14454
rect 20364 14452 20370 14516
rect 21725 14514 21791 14517
rect 22645 14514 22711 14517
rect 21725 14512 22711 14514
rect 21725 14456 21730 14512
rect 21786 14456 22650 14512
rect 22706 14456 22711 14512
rect 21725 14454 22711 14456
rect 21725 14451 21791 14454
rect 22645 14451 22711 14454
rect 12065 14378 12131 14381
rect 20989 14378 21055 14381
rect 12065 14376 21055 14378
rect 12065 14320 12070 14376
rect 12126 14320 20994 14376
rect 21050 14320 21055 14376
rect 12065 14318 21055 14320
rect 12065 14315 12131 14318
rect 20989 14315 21055 14318
rect 22829 14242 22895 14245
rect 26200 14242 27000 14272
rect 22829 14240 27000 14242
rect 22829 14184 22834 14240
rect 22890 14184 27000 14240
rect 22829 14182 27000 14184
rect 22829 14179 22895 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 26200 14152 27000 14182
rect 17946 14111 18262 14112
rect 11605 14106 11671 14109
rect 13486 14106 13492 14108
rect 11605 14104 13492 14106
rect 11605 14048 11610 14104
rect 11666 14048 13492 14104
rect 11605 14046 13492 14048
rect 11605 14043 11671 14046
rect 13486 14044 13492 14046
rect 13556 14044 13562 14108
rect 6545 13970 6611 13973
rect 25129 13970 25195 13973
rect 6545 13968 25195 13970
rect 6545 13912 6550 13968
rect 6606 13912 25134 13968
rect 25190 13912 25195 13968
rect 6545 13910 25195 13912
rect 6545 13907 6611 13910
rect 25129 13907 25195 13910
rect 13721 13834 13787 13837
rect 14457 13834 14523 13837
rect 12758 13774 13554 13834
rect 7097 13698 7163 13701
rect 12758 13698 12818 13774
rect 7097 13696 12818 13698
rect 7097 13640 7102 13696
rect 7158 13640 12818 13696
rect 7097 13638 12818 13640
rect 13494 13698 13554 13774
rect 13721 13832 14523 13834
rect 13721 13776 13726 13832
rect 13782 13776 14462 13832
rect 14518 13776 14523 13832
rect 13721 13774 14523 13776
rect 13721 13771 13787 13774
rect 14457 13771 14523 13774
rect 24577 13834 24643 13837
rect 26200 13834 27000 13864
rect 24577 13832 27000 13834
rect 24577 13776 24582 13832
rect 24638 13776 27000 13832
rect 24577 13774 27000 13776
rect 24577 13771 24643 13774
rect 26200 13744 27000 13774
rect 17166 13698 17172 13700
rect 13494 13638 17172 13698
rect 7097 13635 7163 13638
rect 17166 13636 17172 13638
rect 17236 13636 17242 13700
rect 18597 13698 18663 13701
rect 22185 13698 22251 13701
rect 18597 13696 22251 13698
rect 18597 13640 18602 13696
rect 18658 13640 22190 13696
rect 22246 13640 22251 13696
rect 18597 13638 22251 13640
rect 18597 13635 18663 13638
rect 22185 13635 22251 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 16665 13562 16731 13565
rect 21398 13562 21404 13564
rect 16665 13560 21404 13562
rect 16665 13504 16670 13560
rect 16726 13504 21404 13560
rect 16665 13502 21404 13504
rect 16665 13499 16731 13502
rect 21398 13500 21404 13502
rect 21468 13500 21474 13564
rect 1945 13426 2011 13429
rect 22001 13426 22067 13429
rect 26200 13426 27000 13456
rect 1945 13424 17234 13426
rect 1945 13368 1950 13424
rect 2006 13368 17234 13424
rect 1945 13366 17234 13368
rect 1945 13363 2011 13366
rect 12341 13290 12407 13293
rect 16665 13290 16731 13293
rect 12341 13288 16731 13290
rect 12341 13232 12346 13288
rect 12402 13232 16670 13288
rect 16726 13232 16731 13288
rect 12341 13230 16731 13232
rect 17174 13290 17234 13366
rect 22001 13424 27000 13426
rect 22001 13368 22006 13424
rect 22062 13368 27000 13424
rect 22001 13366 27000 13368
rect 22001 13363 22067 13366
rect 26200 13336 27000 13366
rect 24393 13290 24459 13293
rect 17174 13288 24459 13290
rect 17174 13232 24398 13288
rect 24454 13232 24459 13288
rect 17174 13230 24459 13232
rect 12341 13227 12407 13230
rect 16665 13227 16731 13230
rect 24393 13227 24459 13230
rect 8661 13154 8727 13157
rect 15653 13154 15719 13157
rect 8661 13152 15719 13154
rect 8661 13096 8666 13152
rect 8722 13096 15658 13152
rect 15714 13096 15719 13152
rect 8661 13094 15719 13096
rect 8661 13091 8727 13094
rect 15653 13091 15719 13094
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 10409 13018 10475 13021
rect 16205 13018 16271 13021
rect 10409 13016 16271 13018
rect 10409 12960 10414 13016
rect 10470 12960 16210 13016
rect 16266 12960 16271 13016
rect 10409 12958 16271 12960
rect 10409 12955 10475 12958
rect 16205 12955 16271 12958
rect 24669 13018 24735 13021
rect 26200 13018 27000 13048
rect 24669 13016 27000 13018
rect 24669 12960 24674 13016
rect 24730 12960 27000 13016
rect 24669 12958 27000 12960
rect 24669 12955 24735 12958
rect 26200 12928 27000 12958
rect 16757 12882 16823 12885
rect 23565 12882 23631 12885
rect 16757 12880 23631 12882
rect 16757 12824 16762 12880
rect 16818 12824 23570 12880
rect 23626 12824 23631 12880
rect 16757 12822 23631 12824
rect 16757 12819 16823 12822
rect 23565 12819 23631 12822
rect 8385 12746 8451 12749
rect 19701 12746 19767 12749
rect 8385 12744 19767 12746
rect 8385 12688 8390 12744
rect 8446 12688 19706 12744
rect 19762 12688 19767 12744
rect 8385 12686 19767 12688
rect 8385 12683 8451 12686
rect 19701 12683 19767 12686
rect 25129 12610 25195 12613
rect 26200 12610 27000 12640
rect 25129 12608 27000 12610
rect 25129 12552 25134 12608
rect 25190 12552 27000 12608
rect 25129 12550 27000 12552
rect 25129 12547 25195 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 26200 12520 27000 12550
rect 22946 12479 23262 12480
rect 16665 12474 16731 12477
rect 22134 12474 22140 12476
rect 16665 12472 22140 12474
rect 16665 12416 16670 12472
rect 16726 12416 22140 12472
rect 16665 12414 22140 12416
rect 16665 12411 16731 12414
rect 22134 12412 22140 12414
rect 22204 12412 22210 12476
rect 15193 12338 15259 12341
rect 19241 12338 19307 12341
rect 15193 12336 19307 12338
rect 15193 12280 15198 12336
rect 15254 12280 19246 12336
rect 19302 12280 19307 12336
rect 15193 12278 19307 12280
rect 15193 12275 15259 12278
rect 19241 12275 19307 12278
rect 5533 12202 5599 12205
rect 18689 12202 18755 12205
rect 5533 12200 18755 12202
rect 5533 12144 5538 12200
rect 5594 12144 18694 12200
rect 18750 12144 18755 12200
rect 5533 12142 18755 12144
rect 5533 12139 5599 12142
rect 18689 12139 18755 12142
rect 24761 12202 24827 12205
rect 26200 12202 27000 12232
rect 24761 12200 27000 12202
rect 24761 12144 24766 12200
rect 24822 12144 27000 12200
rect 24761 12142 27000 12144
rect 24761 12139 24827 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 15837 11930 15903 11933
rect 16062 11930 16068 11932
rect 15837 11928 16068 11930
rect 15837 11872 15842 11928
rect 15898 11872 16068 11928
rect 15837 11870 16068 11872
rect 15837 11867 15903 11870
rect 16062 11868 16068 11870
rect 16132 11868 16138 11932
rect 7005 11794 7071 11797
rect 20069 11794 20135 11797
rect 7005 11792 20135 11794
rect 7005 11736 7010 11792
rect 7066 11736 20074 11792
rect 20130 11736 20135 11792
rect 7005 11734 20135 11736
rect 7005 11731 7071 11734
rect 20069 11731 20135 11734
rect 24853 11794 24919 11797
rect 26200 11794 27000 11824
rect 24853 11792 27000 11794
rect 24853 11736 24858 11792
rect 24914 11736 27000 11792
rect 24853 11734 27000 11736
rect 24853 11731 24919 11734
rect 26200 11704 27000 11734
rect 19425 11658 19491 11661
rect 23841 11658 23907 11661
rect 19425 11656 23907 11658
rect 19425 11600 19430 11656
rect 19486 11600 23846 11656
rect 23902 11600 23907 11656
rect 19425 11598 23907 11600
rect 19425 11595 19491 11598
rect 23841 11595 23907 11598
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 17401 11386 17467 11389
rect 17534 11386 17540 11388
rect 17401 11384 17540 11386
rect 17401 11328 17406 11384
rect 17462 11328 17540 11384
rect 17401 11326 17540 11328
rect 17401 11323 17467 11326
rect 17534 11324 17540 11326
rect 17604 11324 17610 11388
rect 20161 11386 20227 11389
rect 18462 11384 20227 11386
rect 18462 11328 20166 11384
rect 20222 11328 20227 11384
rect 18462 11326 20227 11328
rect 6494 11188 6500 11252
rect 6564 11250 6570 11252
rect 18462 11250 18522 11326
rect 20161 11323 20227 11326
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 6564 11190 18522 11250
rect 18689 11250 18755 11253
rect 19425 11250 19491 11253
rect 18689 11248 19491 11250
rect 18689 11192 18694 11248
rect 18750 11192 19430 11248
rect 19486 11192 19491 11248
rect 18689 11190 19491 11192
rect 6564 11188 6570 11190
rect 18689 11187 18755 11190
rect 19425 11187 19491 11190
rect 17718 11052 17724 11116
rect 17788 11114 17794 11116
rect 17861 11114 17927 11117
rect 17788 11112 17927 11114
rect 17788 11056 17866 11112
rect 17922 11056 17927 11112
rect 17788 11054 17927 11056
rect 17788 11052 17794 11054
rect 17861 11051 17927 11054
rect 18454 11052 18460 11116
rect 18524 11114 18530 11116
rect 18597 11114 18663 11117
rect 18524 11112 18663 11114
rect 18524 11056 18602 11112
rect 18658 11056 18663 11112
rect 18524 11054 18663 11056
rect 18524 11052 18530 11054
rect 18597 11051 18663 11054
rect 19609 10978 19675 10981
rect 19926 10978 19932 10980
rect 19609 10976 19932 10978
rect 19609 10920 19614 10976
rect 19670 10920 19932 10976
rect 19609 10918 19932 10920
rect 19609 10915 19675 10918
rect 19926 10916 19932 10918
rect 19996 10916 20002 10980
rect 24669 10978 24735 10981
rect 26200 10978 27000 11008
rect 24669 10976 27000 10978
rect 24669 10920 24674 10976
rect 24730 10920 27000 10976
rect 24669 10918 27000 10920
rect 24669 10915 24735 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 26200 10888 27000 10918
rect 17946 10847 18262 10848
rect 19333 10842 19399 10845
rect 20069 10842 20135 10845
rect 22502 10842 22508 10844
rect 19333 10840 22508 10842
rect 19333 10784 19338 10840
rect 19394 10784 20074 10840
rect 20130 10784 22508 10840
rect 19333 10782 22508 10784
rect 19333 10779 19399 10782
rect 20069 10779 20135 10782
rect 22502 10780 22508 10782
rect 22572 10780 22578 10844
rect 16297 10706 16363 10709
rect 25957 10706 26023 10709
rect 16297 10704 26023 10706
rect 16297 10648 16302 10704
rect 16358 10648 25962 10704
rect 26018 10648 26023 10704
rect 16297 10646 26023 10648
rect 16297 10643 16363 10646
rect 25957 10643 26023 10646
rect 12709 10570 12775 10573
rect 21265 10570 21331 10573
rect 12709 10568 21331 10570
rect 12709 10512 12714 10568
rect 12770 10512 21270 10568
rect 21326 10512 21331 10568
rect 12709 10510 21331 10512
rect 12709 10507 12775 10510
rect 21265 10507 21331 10510
rect 24853 10570 24919 10573
rect 26200 10570 27000 10600
rect 24853 10568 27000 10570
rect 24853 10512 24858 10568
rect 24914 10512 27000 10568
rect 24853 10510 27000 10512
rect 24853 10507 24919 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 19885 10298 19951 10301
rect 21081 10298 21147 10301
rect 21950 10298 21956 10300
rect 19885 10296 21956 10298
rect 19885 10240 19890 10296
rect 19946 10240 21086 10296
rect 21142 10240 21956 10296
rect 19885 10238 21956 10240
rect 19885 10235 19951 10238
rect 21081 10235 21147 10238
rect 21950 10236 21956 10238
rect 22020 10236 22026 10300
rect 24761 10162 24827 10165
rect 26200 10162 27000 10192
rect 24761 10160 27000 10162
rect 24761 10104 24766 10160
rect 24822 10104 27000 10160
rect 24761 10102 27000 10104
rect 24761 10099 24827 10102
rect 26200 10072 27000 10102
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 20897 9754 20963 9757
rect 21766 9754 21772 9756
rect 20897 9752 21772 9754
rect 20897 9696 20902 9752
rect 20958 9696 21772 9752
rect 20897 9694 21772 9696
rect 20897 9691 20963 9694
rect 21766 9692 21772 9694
rect 21836 9692 21842 9756
rect 23289 9754 23355 9757
rect 26200 9754 27000 9784
rect 23289 9752 27000 9754
rect 23289 9696 23294 9752
rect 23350 9696 27000 9752
rect 23289 9694 27000 9696
rect 23289 9691 23355 9694
rect 26200 9664 27000 9694
rect 20110 9556 20116 9620
rect 20180 9618 20186 9620
rect 21449 9618 21515 9621
rect 20180 9616 21515 9618
rect 20180 9560 21454 9616
rect 21510 9560 21515 9616
rect 20180 9558 21515 9560
rect 20180 9556 20186 9558
rect 21449 9555 21515 9558
rect 17585 9482 17651 9485
rect 24710 9482 24716 9484
rect 17585 9480 24716 9482
rect 17585 9424 17590 9480
rect 17646 9424 24716 9480
rect 17585 9422 24716 9424
rect 17585 9419 17651 9422
rect 24710 9420 24716 9422
rect 24780 9420 24786 9484
rect 24853 9346 24919 9349
rect 26200 9346 27000 9376
rect 24853 9344 27000 9346
rect 24853 9288 24858 9344
rect 24914 9288 27000 9344
rect 24853 9286 27000 9288
rect 24853 9283 24919 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 26200 9256 27000 9286
rect 22946 9215 23262 9216
rect 15878 9148 15884 9212
rect 15948 9210 15954 9212
rect 19425 9210 19491 9213
rect 15948 9208 19491 9210
rect 15948 9152 19430 9208
rect 19486 9152 19491 9208
rect 15948 9150 19491 9152
rect 15948 9148 15954 9150
rect 19425 9147 19491 9150
rect 6678 9012 6684 9076
rect 6748 9074 6754 9076
rect 22001 9074 22067 9077
rect 6748 9072 22067 9074
rect 6748 9016 22006 9072
rect 22062 9016 22067 9072
rect 6748 9014 22067 9016
rect 6748 9012 6754 9014
rect 22001 9011 22067 9014
rect 25129 8938 25195 8941
rect 26200 8938 27000 8968
rect 25129 8936 27000 8938
rect 25129 8880 25134 8936
rect 25190 8880 27000 8936
rect 25129 8878 27000 8880
rect 25129 8875 25195 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 24853 8530 24919 8533
rect 26200 8530 27000 8560
rect 24853 8528 27000 8530
rect 24853 8472 24858 8528
rect 24914 8472 27000 8528
rect 24853 8470 27000 8472
rect 24853 8467 24919 8470
rect 26200 8440 27000 8470
rect 19742 8332 19748 8396
rect 19812 8394 19818 8396
rect 20345 8394 20411 8397
rect 19812 8392 20411 8394
rect 19812 8336 20350 8392
rect 20406 8336 20411 8392
rect 19812 8334 20411 8336
rect 19812 8332 19818 8334
rect 20345 8331 20411 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24853 8122 24919 8125
rect 26200 8122 27000 8152
rect 24853 8120 27000 8122
rect 24853 8064 24858 8120
rect 24914 8064 27000 8120
rect 24853 8062 27000 8064
rect 24853 8059 24919 8062
rect 26200 8032 27000 8062
rect 24761 7714 24827 7717
rect 26200 7714 27000 7744
rect 24761 7712 27000 7714
rect 24761 7656 24766 7712
rect 24822 7656 27000 7712
rect 24761 7654 27000 7656
rect 24761 7651 24827 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 24945 6898 25011 6901
rect 26200 6898 27000 6928
rect 24945 6896 27000 6898
rect 24945 6840 24950 6896
rect 25006 6840 27000 6896
rect 24945 6838 27000 6840
rect 24945 6835 25011 6838
rect 26200 6808 27000 6838
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 24669 6490 24735 6493
rect 26200 6490 27000 6520
rect 24669 6488 27000 6490
rect 24669 6432 24674 6488
rect 24730 6432 27000 6488
rect 24669 6430 27000 6432
rect 24669 6427 24735 6430
rect 26200 6400 27000 6430
rect 24853 6082 24919 6085
rect 26200 6082 27000 6112
rect 24853 6080 27000 6082
rect 24853 6024 24858 6080
rect 24914 6024 27000 6080
rect 24853 6022 27000 6024
rect 24853 6019 24919 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 26200 5992 27000 6022
rect 22946 5951 23262 5952
rect 24945 5674 25011 5677
rect 26200 5674 27000 5704
rect 24945 5672 27000 5674
rect 24945 5616 24950 5672
rect 25006 5616 27000 5672
rect 24945 5614 27000 5616
rect 24945 5611 25011 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 24761 5266 24827 5269
rect 26200 5266 27000 5296
rect 24761 5264 27000 5266
rect 24761 5208 24766 5264
rect 24822 5208 27000 5264
rect 24761 5206 27000 5208
rect 24761 5203 24827 5206
rect 26200 5176 27000 5206
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24853 4858 24919 4861
rect 26200 4858 27000 4888
rect 24853 4856 27000 4858
rect 24853 4800 24858 4856
rect 24914 4800 27000 4856
rect 24853 4798 27000 4800
rect 24853 4795 24919 4798
rect 26200 4768 27000 4798
rect 24945 4450 25011 4453
rect 26200 4450 27000 4480
rect 24945 4448 27000 4450
rect 24945 4392 24950 4448
rect 25006 4392 27000 4448
rect 24945 4390 27000 4392
rect 24945 4387 25011 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 26200 4360 27000 4390
rect 17946 4319 18262 4320
rect 25129 4042 25195 4045
rect 26200 4042 27000 4072
rect 25129 4040 27000 4042
rect 25129 3984 25134 4040
rect 25190 3984 27000 4040
rect 25129 3982 27000 3984
rect 25129 3979 25195 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 24945 3634 25011 3637
rect 26200 3634 27000 3664
rect 24945 3632 27000 3634
rect 24945 3576 24950 3632
rect 25006 3576 27000 3632
rect 24945 3574 27000 3576
rect 24945 3571 25011 3574
rect 26200 3544 27000 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 24945 3226 25011 3229
rect 26200 3226 27000 3256
rect 24945 3224 27000 3226
rect 24945 3168 24950 3224
rect 25006 3168 27000 3224
rect 24945 3166 27000 3168
rect 24945 3163 25011 3166
rect 26200 3136 27000 3166
rect 24853 2818 24919 2821
rect 26200 2818 27000 2848
rect 24853 2816 27000 2818
rect 24853 2760 24858 2816
rect 24914 2760 27000 2816
rect 24853 2758 27000 2760
rect 24853 2755 24919 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 26200 2728 27000 2758
rect 22946 2687 23262 2688
rect 24945 2410 25011 2413
rect 26200 2410 27000 2440
rect 24945 2408 27000 2410
rect 24945 2352 24950 2408
rect 25006 2352 27000 2408
rect 24945 2350 27000 2352
rect 24945 2347 25011 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 22829 2002 22895 2005
rect 26200 2002 27000 2032
rect 22829 2000 27000 2002
rect 22829 1944 22834 2000
rect 22890 1944 27000 2000
rect 22829 1942 27000 1944
rect 22829 1939 22895 1942
rect 26200 1912 27000 1942
rect 22093 1594 22159 1597
rect 26200 1594 27000 1624
rect 22093 1592 27000 1594
rect 22093 1536 22098 1592
rect 22154 1536 27000 1592
rect 22093 1534 27000 1536
rect 22093 1531 22159 1534
rect 26200 1504 27000 1534
rect 22093 1186 22159 1189
rect 26200 1186 27000 1216
rect 22093 1184 27000 1186
rect 22093 1128 22098 1184
rect 22154 1128 27000 1184
rect 22093 1126 27000 1128
rect 22093 1123 22159 1126
rect 26200 1096 27000 1126
rect 25037 778 25103 781
rect 26200 778 27000 808
rect 25037 776 27000 778
rect 25037 720 25042 776
rect 25098 720 27000 776
rect 25037 718 27000 720
rect 25037 715 25103 718
rect 26200 688 27000 718
rect 23381 370 23447 373
rect 26200 370 27000 400
rect 23381 368 27000 370
rect 23381 312 23386 368
rect 23442 312 27000 368
rect 23381 310 27000 312
rect 23381 307 23447 310
rect 26200 280 27000 310
<< via3 >>
rect 2268 26284 2332 26348
rect 4108 26148 4172 26212
rect 19564 25604 19628 25668
rect 5028 25468 5092 25532
rect 7788 25332 7852 25396
rect 4844 25196 4908 25260
rect 19380 25196 19444 25260
rect 10732 25060 10796 25124
rect 13492 24788 13556 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 6684 24168 6748 24172
rect 6684 24112 6734 24168
rect 6734 24112 6748 24168
rect 6684 24108 6748 24112
rect 8524 23972 8588 24036
rect 21404 23972 21468 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 9076 23564 9140 23628
rect 6500 23488 6564 23492
rect 6500 23432 6550 23488
rect 6550 23432 6564 23488
rect 6500 23428 6564 23432
rect 7420 23428 7484 23492
rect 12572 23428 12636 23492
rect 16620 23428 16684 23492
rect 19380 23428 19444 23492
rect 19932 23488 19996 23492
rect 19932 23432 19946 23488
rect 19946 23432 19996 23488
rect 19932 23428 19996 23432
rect 20300 23428 20364 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 22140 23156 22204 23220
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 8340 22748 8404 22812
rect 19748 22476 19812 22540
rect 16068 22340 16132 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 13860 22204 13924 22268
rect 10180 22068 10244 22132
rect 21772 21796 21836 21860
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 19564 21660 19628 21724
rect 4844 21584 4908 21588
rect 4844 21528 4858 21584
rect 4858 21528 4908 21584
rect 4844 21524 4908 21528
rect 21956 21524 22020 21588
rect 22508 21388 22572 21452
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 11100 20708 11164 20772
rect 15884 20768 15948 20772
rect 15884 20712 15898 20768
rect 15898 20712 15948 20768
rect 15884 20708 15948 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 17172 20300 17236 20364
rect 18460 20164 18524 20228
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7788 20028 7852 20092
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 7236 19544 7300 19548
rect 7236 19488 7286 19544
rect 7286 19488 7300 19544
rect 7236 19484 7300 19488
rect 8340 19348 8404 19412
rect 17540 19348 17604 19412
rect 20116 19348 20180 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 22324 18940 22388 19004
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 4108 18320 4172 18324
rect 4108 18264 4122 18320
rect 4122 18264 4172 18320
rect 4108 18260 4172 18264
rect 13860 18260 13924 18324
rect 7420 17988 7484 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 17724 18048 17788 18052
rect 17724 17992 17738 18048
rect 17738 17992 17788 18048
rect 17724 17988 17788 17992
rect 24716 17988 24780 18052
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 5028 17716 5092 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 12388 17172 12452 17236
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 11100 17036 11164 17100
rect 22692 17036 22756 17100
rect 19380 16900 19444 16964
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 8524 16764 8588 16828
rect 9076 16824 9140 16828
rect 9076 16768 9090 16824
rect 9090 16768 9140 16824
rect 9076 16764 9140 16768
rect 10180 16764 10244 16828
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 2268 16084 2332 16148
rect 7236 16008 7300 16012
rect 7236 15952 7286 16008
rect 7286 15952 7300 16008
rect 7236 15948 7300 15952
rect 22324 15812 22388 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 19380 15676 19444 15740
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 10732 14996 10796 15060
rect 22692 14724 22756 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 16620 14452 16684 14516
rect 20300 14452 20364 14516
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 13492 14044 13556 14108
rect 17172 13636 17236 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 21404 13500 21468 13564
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 22140 12412 22204 12476
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 16068 11868 16132 11932
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 17540 11324 17604 11388
rect 6500 11188 6564 11252
rect 17724 11052 17788 11116
rect 18460 11052 18524 11116
rect 19932 10916 19996 10980
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 22508 10780 22572 10844
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 21956 10236 22020 10300
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 21772 9692 21836 9756
rect 20116 9556 20180 9620
rect 24716 9420 24780 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 15884 9148 15948 9212
rect 6684 9012 6748 9076
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 19748 8332 19812 8396
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2267 26348 2333 26349
rect 2267 26284 2268 26348
rect 2332 26284 2333 26348
rect 2267 26283 2333 26284
rect 2270 16149 2330 26283
rect 4107 26212 4173 26213
rect 4107 26148 4108 26212
rect 4172 26148 4173 26212
rect 4107 26147 4173 26148
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 4110 18325 4170 26147
rect 19563 25668 19629 25669
rect 19563 25604 19564 25668
rect 19628 25604 19629 25668
rect 19563 25603 19629 25604
rect 5027 25532 5093 25533
rect 5027 25468 5028 25532
rect 5092 25468 5093 25532
rect 5027 25467 5093 25468
rect 4843 25260 4909 25261
rect 4843 25196 4844 25260
rect 4908 25196 4909 25260
rect 4843 25195 4909 25196
rect 4846 21589 4906 25195
rect 4843 21588 4909 21589
rect 4843 21524 4844 21588
rect 4908 21524 4909 21588
rect 4843 21523 4909 21524
rect 4107 18324 4173 18325
rect 4107 18260 4108 18324
rect 4172 18260 4173 18324
rect 4107 18259 4173 18260
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 5030 17781 5090 25467
rect 7787 25396 7853 25397
rect 7787 25332 7788 25396
rect 7852 25332 7853 25396
rect 7787 25331 7853 25332
rect 6683 24172 6749 24173
rect 6683 24108 6684 24172
rect 6748 24108 6749 24172
rect 6683 24107 6749 24108
rect 6499 23492 6565 23493
rect 6499 23428 6500 23492
rect 6564 23428 6565 23492
rect 6499 23427 6565 23428
rect 5027 17780 5093 17781
rect 5027 17716 5028 17780
rect 5092 17716 5093 17780
rect 5027 17715 5093 17716
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2267 16148 2333 16149
rect 2267 16084 2268 16148
rect 2332 16084 2333 16148
rect 2267 16083 2333 16084
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 6502 11253 6562 23427
rect 6499 11252 6565 11253
rect 6499 11188 6500 11252
rect 6564 11188 6565 11252
rect 6499 11187 6565 11188
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 6686 9077 6746 24107
rect 7419 23492 7485 23493
rect 7419 23428 7420 23492
rect 7484 23428 7485 23492
rect 7419 23427 7485 23428
rect 7235 19548 7301 19549
rect 7235 19484 7236 19548
rect 7300 19484 7301 19548
rect 7235 19483 7301 19484
rect 7238 16013 7298 19483
rect 7422 18053 7482 23427
rect 7790 20093 7850 25331
rect 19379 25260 19445 25261
rect 19379 25196 19380 25260
rect 19444 25196 19445 25260
rect 19379 25195 19445 25196
rect 10731 25124 10797 25125
rect 10731 25060 10732 25124
rect 10796 25060 10797 25124
rect 10731 25059 10797 25060
rect 7944 23968 8264 24528
rect 8523 24036 8589 24037
rect 8523 23972 8524 24036
rect 8588 23972 8589 24036
rect 8523 23971 8589 23972
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 8339 22812 8405 22813
rect 8339 22748 8340 22812
rect 8404 22748 8405 22812
rect 8339 22747 8405 22748
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7787 20092 7853 20093
rect 7787 20028 7788 20092
rect 7852 20028 7853 20092
rect 7787 20027 7853 20028
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 8342 19413 8402 22747
rect 8339 19412 8405 19413
rect 8339 19348 8340 19412
rect 8404 19348 8405 19412
rect 8339 19347 8405 19348
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7419 18052 7485 18053
rect 7419 17988 7420 18052
rect 7484 17988 7485 18052
rect 7419 17987 7485 17988
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 8526 16829 8586 23971
rect 9075 23628 9141 23629
rect 9075 23564 9076 23628
rect 9140 23564 9141 23628
rect 9075 23563 9141 23564
rect 9078 16829 9138 23563
rect 10179 22132 10245 22133
rect 10179 22068 10180 22132
rect 10244 22068 10245 22132
rect 10179 22067 10245 22068
rect 10182 16829 10242 22067
rect 8523 16828 8589 16829
rect 8523 16764 8524 16828
rect 8588 16764 8589 16828
rect 8523 16763 8589 16764
rect 9075 16828 9141 16829
rect 9075 16764 9076 16828
rect 9140 16764 9141 16828
rect 9075 16763 9141 16764
rect 10179 16828 10245 16829
rect 10179 16764 10180 16828
rect 10244 16764 10245 16828
rect 10179 16763 10245 16764
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7235 16012 7301 16013
rect 7235 15948 7236 16012
rect 7300 15948 7301 16012
rect 7235 15947 7301 15948
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 10734 15061 10794 25059
rect 13491 24852 13557 24853
rect 13491 24788 13492 24852
rect 13556 24788 13557 24852
rect 13491 24787 13557 24788
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23428 12637 23492
rect 12571 23427 12637 23428
rect 11099 20772 11165 20773
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 11102 17101 11162 20707
rect 12574 17370 12634 23427
rect 12390 17310 12634 17370
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12390 17237 12450 17310
rect 12387 17236 12453 17237
rect 12387 17172 12388 17236
rect 12452 17172 12453 17236
rect 12387 17171 12453 17172
rect 11099 17100 11165 17101
rect 11099 17036 11100 17100
rect 11164 17036 11165 17100
rect 11099 17035 11165 17036
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 10731 15060 10797 15061
rect 10731 14996 10732 15060
rect 10796 14996 10797 15060
rect 10731 14995 10797 14996
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 6683 9076 6749 9077
rect 6683 9012 6684 9076
rect 6748 9012 6749 9076
rect 6683 9011 6749 9012
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 13494 14109 13554 24787
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 16619 23492 16685 23493
rect 16619 23428 16620 23492
rect 16684 23428 16685 23492
rect 16619 23427 16685 23428
rect 16067 22404 16133 22405
rect 16067 22340 16068 22404
rect 16132 22340 16133 22404
rect 16067 22339 16133 22340
rect 13859 22268 13925 22269
rect 13859 22204 13860 22268
rect 13924 22204 13925 22268
rect 13859 22203 13925 22204
rect 13862 18325 13922 22203
rect 15883 20772 15949 20773
rect 15883 20708 15884 20772
rect 15948 20708 15949 20772
rect 15883 20707 15949 20708
rect 13859 18324 13925 18325
rect 13859 18260 13860 18324
rect 13924 18260 13925 18324
rect 13859 18259 13925 18260
rect 13491 14108 13557 14109
rect 13491 14044 13492 14108
rect 13556 14044 13557 14108
rect 13491 14043 13557 14044
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 15886 9213 15946 20707
rect 16070 11933 16130 22339
rect 16622 14517 16682 23427
rect 17944 22880 18264 23904
rect 19382 23493 19442 25195
rect 19379 23492 19445 23493
rect 19379 23428 19380 23492
rect 19444 23428 19445 23492
rect 19379 23427 19445 23428
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 19566 21725 19626 25603
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 21403 24036 21469 24037
rect 21403 23972 21404 24036
rect 21468 23972 21469 24036
rect 21403 23971 21469 23972
rect 19931 23492 19997 23493
rect 19931 23428 19932 23492
rect 19996 23428 19997 23492
rect 19931 23427 19997 23428
rect 20299 23492 20365 23493
rect 20299 23428 20300 23492
rect 20364 23428 20365 23492
rect 20299 23427 20365 23428
rect 19747 22540 19813 22541
rect 19747 22476 19748 22540
rect 19812 22476 19813 22540
rect 19747 22475 19813 22476
rect 19563 21724 19629 21725
rect 19563 21660 19564 21724
rect 19628 21660 19629 21724
rect 19563 21659 19629 21660
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17171 20364 17237 20365
rect 17171 20300 17172 20364
rect 17236 20300 17237 20364
rect 17171 20299 17237 20300
rect 16619 14516 16685 14517
rect 16619 14452 16620 14516
rect 16684 14452 16685 14516
rect 16619 14451 16685 14452
rect 17174 13701 17234 20299
rect 17944 19616 18264 20640
rect 18459 20228 18525 20229
rect 18459 20164 18460 20228
rect 18524 20164 18525 20228
rect 18459 20163 18525 20164
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 17171 13700 17237 13701
rect 17171 13636 17172 13700
rect 17236 13636 17237 13700
rect 17171 13635 17237 13636
rect 16067 11932 16133 11933
rect 16067 11868 16068 11932
rect 16132 11868 16133 11932
rect 16067 11867 16133 11868
rect 17542 11389 17602 19347
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17723 18052 17789 18053
rect 17723 17988 17724 18052
rect 17788 17988 17789 18052
rect 17723 17987 17789 17988
rect 17539 11388 17605 11389
rect 17539 11324 17540 11388
rect 17604 11324 17605 11388
rect 17539 11323 17605 11324
rect 17726 11117 17786 17987
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17723 11116 17789 11117
rect 17723 11052 17724 11116
rect 17788 11052 17789 11116
rect 17723 11051 17789 11052
rect 17944 10912 18264 11936
rect 18462 11117 18522 20163
rect 19379 16964 19445 16965
rect 19379 16900 19380 16964
rect 19444 16900 19445 16964
rect 19379 16899 19445 16900
rect 19382 15741 19442 16899
rect 19379 15740 19445 15741
rect 19379 15676 19380 15740
rect 19444 15676 19445 15740
rect 19379 15675 19445 15676
rect 18459 11116 18525 11117
rect 18459 11052 18460 11116
rect 18524 11052 18525 11116
rect 18459 11051 18525 11052
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 15883 9212 15949 9213
rect 15883 9148 15884 9212
rect 15948 9148 15949 9212
rect 15883 9147 15949 9148
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 19750 8397 19810 22475
rect 19934 10981 19994 23427
rect 20115 19412 20181 19413
rect 20115 19348 20116 19412
rect 20180 19348 20181 19412
rect 20115 19347 20181 19348
rect 19931 10980 19997 10981
rect 19931 10916 19932 10980
rect 19996 10916 19997 10980
rect 19931 10915 19997 10916
rect 20118 9621 20178 19347
rect 20302 14517 20362 23427
rect 20299 14516 20365 14517
rect 20299 14452 20300 14516
rect 20364 14452 20365 14516
rect 20299 14451 20365 14452
rect 21406 13565 21466 23971
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22139 23220 22205 23221
rect 22139 23156 22140 23220
rect 22204 23156 22205 23220
rect 22139 23155 22205 23156
rect 21771 21860 21837 21861
rect 21771 21796 21772 21860
rect 21836 21796 21837 21860
rect 21771 21795 21837 21796
rect 21403 13564 21469 13565
rect 21403 13500 21404 13564
rect 21468 13500 21469 13564
rect 21403 13499 21469 13500
rect 21774 9757 21834 21795
rect 21955 21588 22021 21589
rect 21955 21524 21956 21588
rect 22020 21524 22021 21588
rect 21955 21523 22021 21524
rect 21958 10301 22018 21523
rect 22142 12477 22202 23155
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22507 21452 22573 21453
rect 22507 21388 22508 21452
rect 22572 21388 22573 21452
rect 22507 21387 22573 21388
rect 22323 19004 22389 19005
rect 22323 18940 22324 19004
rect 22388 18940 22389 19004
rect 22323 18939 22389 18940
rect 22326 15877 22386 18939
rect 22323 15876 22389 15877
rect 22323 15812 22324 15876
rect 22388 15812 22389 15876
rect 22323 15811 22389 15812
rect 22139 12476 22205 12477
rect 22139 12412 22140 12476
rect 22204 12412 22205 12476
rect 22139 12411 22205 12412
rect 22510 10845 22570 21387
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 24715 18052 24781 18053
rect 24715 17988 24716 18052
rect 24780 17988 24781 18052
rect 24715 17987 24781 17988
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22691 17100 22757 17101
rect 22691 17036 22692 17100
rect 22756 17036 22757 17100
rect 22691 17035 22757 17036
rect 22694 14789 22754 17035
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22691 14788 22757 14789
rect 22691 14724 22692 14788
rect 22756 14724 22757 14788
rect 22691 14723 22757 14724
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22507 10844 22573 10845
rect 22507 10780 22508 10844
rect 22572 10780 22573 10844
rect 22507 10779 22573 10780
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 21955 10300 22021 10301
rect 21955 10236 21956 10300
rect 22020 10236 22021 10300
rect 21955 10235 22021 10236
rect 21771 9756 21837 9757
rect 21771 9692 21772 9756
rect 21836 9692 21837 9756
rect 21771 9691 21837 9692
rect 20115 9620 20181 9621
rect 20115 9556 20116 9620
rect 20180 9556 20181 9620
rect 20115 9555 20181 9556
rect 22944 9280 23264 10304
rect 24718 9485 24778 17987
rect 24715 9484 24781 9485
rect 24715 9420 24716 9484
rect 24780 9420 24781 9484
rect 24715 9419 24781 9420
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 19747 8396 19813 8397
rect 19747 8332 19748 8396
rect 19812 8332 19813 8396
rect 19747 8331 19813 8332
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1679235063
transform 1 0 19596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1679235063
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1679235063
transform 1 0 25024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1679235063
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1679235063
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1679235063
transform 1 0 23736 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1679235063
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1679235063
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1679235063
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18032 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1679235063
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1679235063
transform 1 0 21160 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1679235063
transform 1 0 23736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1679235063
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1679235063
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1679235063
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1679235063
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1679235063
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _096_
timestamp 1679235063
transform 1 0 14444 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1679235063
transform 1 0 20056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1679235063
transform 1 0 18032 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1679235063
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_
timestamp 1679235063
transform 1 0 12880 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _101_
timestamp 1679235063
transform 1 0 21252 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1679235063
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1679235063
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1679235063
transform 1 0 4508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1679235063
transform 1 0 5244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1679235063
transform 1 0 2576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform 1 0 6808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1679235063
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _115_
timestamp 1679235063
transform 1 0 4508 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1679235063
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1679235063
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 18400 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _122_
timestamp 1679235063
transform 1 0 3220 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _123_
timestamp 1679235063
transform 1 0 4508 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _124_
timestamp 1679235063
transform 1 0 5152 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1679235063
transform 1 0 4508 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_
timestamp 1679235063
transform 1 0 6440 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1679235063
transform 1 0 2576 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1679235063
transform 1 0 5152 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _129_
timestamp 1679235063
transform 1 0 3956 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1679235063
transform 1 0 5152 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1679235063
transform 1 0 4508 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 8188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 13892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 9476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 20240 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 20240 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 2392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 20148 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1679235063
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1679235063
transform 1 0 20148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1679235063
transform 1 0 24932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1679235063
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1679235063
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1679235063
transform 1 0 25300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1679235063
transform 1 0 20608 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1679235063
transform 1 0 25300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1679235063
transform 1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1679235063
transform 1 0 20240 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1679235063
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform 1 0 19596 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 6440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform 1 0 15088 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1679235063
transform 1 0 21252 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1679235063
transform 1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_prog_clk_A
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_prog_clk_A
timestamp 1679235063
transform 1 0 14996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_prog_clk_A
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_prog_clk_A
timestamp 1679235063
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_prog_clk_A
timestamp 1679235063
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_prog_clk_A
timestamp 1679235063
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold1_A
timestamp 1679235063
transform 1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1679235063
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold5_A
timestamp 1679235063
transform 1 0 6440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold7_A
timestamp 1679235063
transform 1 0 19596 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold10_A
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold11_A
timestamp 1679235063
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold13_A
timestamp 1679235063
transform 1 0 20792 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold14_A
timestamp 1679235063
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold15_A
timestamp 1679235063
transform 1 0 25300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold16_A
timestamp 1679235063
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold17_A
timestamp 1679235063
transform 1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold18_A
timestamp 1679235063
transform 1 0 16192 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold19_A
timestamp 1679235063
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold20_A
timestamp 1679235063
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold21_A
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold22_A
timestamp 1679235063
transform 1 0 25300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold23_A
timestamp 1679235063
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold24_A
timestamp 1679235063
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold25_A
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold26_A
timestamp 1679235063
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold27_A
timestamp 1679235063
transform 1 0 1472 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold28_A
timestamp 1679235063
transform 1 0 1472 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold29_A
timestamp 1679235063
transform 1 0 24656 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold30_A
timestamp 1679235063
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold31_A
timestamp 1679235063
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold32_A
timestamp 1679235063
transform 1 0 2392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold33_A
timestamp 1679235063
transform 1 0 1564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold34_A
timestamp 1679235063
transform 1 0 24472 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold35_A
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold36_A
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold37_A
timestamp 1679235063
transform 1 0 6440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 7820 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 19872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 20884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 19964 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 10580 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 20240 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 2024 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 5796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 6624 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 20056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 8004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 1656 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 24564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 9016 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 1656 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 2116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output102_A
timestamp 1679235063
transform 1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output110_A
timestamp 1679235063
transform 1 0 1472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20424 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 1472 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 1656 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24196 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23000 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 13984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9200 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21068 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16008 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12696 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 23368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 17664 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22816 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23184 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 20608 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 2208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 6808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13248 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21436 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4232 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17112 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1679235063
transform 1 0 9568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1679235063
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1679235063
transform 1 0 10396 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1679235063
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1679235063
transform 1 0 18216 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1679235063
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1679235063
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1679235063
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1679235063
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1679235063
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1679235063
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1679235063
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1679235063
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1679235063
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1679235063
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1679235063
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1679235063
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1679235063
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1679235063
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1679235063
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1679235063
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1679235063
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1679235063
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_60
timestamp 1679235063
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_70
timestamp 1679235063
transform 1 0 7544 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_82
timestamp 1679235063
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1679235063
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1679235063
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1679235063
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1679235063
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1679235063
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1679235063
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1679235063
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1679235063
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1679235063
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1679235063
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_53
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1679235063
transform 1 0 6716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_70
timestamp 1679235063
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1679235063
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1679235063
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1679235063
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1679235063
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1679235063
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1679235063
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1679235063
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1679235063
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_259
timestamp 1679235063
transform 1 0 24932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_265
timestamp 1679235063
transform 1 0 25484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1679235063
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1679235063
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1679235063
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1679235063
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1679235063
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1679235063
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1679235063
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1679235063
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1679235063
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1679235063
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_205
timestamp 1679235063
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1679235063
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1679235063
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp 1679235063
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1679235063
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1679235063
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_209
timestamp 1679235063
transform 1 0 20332 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_217
timestamp 1679235063
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1679235063
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1679235063
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_259
timestamp 1679235063
transform 1 0 24932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_263
timestamp 1679235063
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1679235063
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1679235063
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp 1679235063
transform 1 0 21068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1679235063
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1679235063
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1679235063
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1679235063
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1679235063
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_222
timestamp 1679235063
transform 1 0 21528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_226
timestamp 1679235063
transform 1 0 21896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1679235063
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1679235063
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_259
timestamp 1679235063
transform 1 0 24932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_90
timestamp 1679235063
transform 1 0 9384 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1679235063
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1679235063
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_205
timestamp 1679235063
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1679235063
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1679235063
transform 1 0 20884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1679235063
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1679235063
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_208
timestamp 1679235063
transform 1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1679235063
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1679235063
transform 1 0 22172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_233
timestamp 1679235063
transform 1 0 22540 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_259
timestamp 1679235063
transform 1 0 24932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1679235063
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1679235063
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1679235063
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_208
timestamp 1679235063
transform 1 0 20240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1679235063
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1679235063
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1679235063
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1679235063
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1679235063
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1679235063
transform 1 0 19780 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_208
timestamp 1679235063
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_212
timestamp 1679235063
transform 1 0 20608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_216
timestamp 1679235063
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1679235063
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1679235063
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_258
timestamp 1679235063
transform 1 0 24840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_264
timestamp 1679235063
transform 1 0 25392 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1679235063
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1679235063
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1679235063
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1679235063
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1679235063
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_189
timestamp 1679235063
transform 1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_195
timestamp 1679235063
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_202
timestamp 1679235063
transform 1 0 19688 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_210
timestamp 1679235063
transform 1 0 20424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1679235063
transform 1 0 20884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1679235063
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1679235063
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1679235063
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1679235063
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1679235063
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1679235063
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1679235063
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1679235063
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_177
timestamp 1679235063
transform 1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1679235063
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1679235063
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_209
timestamp 1679235063
transform 1 0 20332 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_218
timestamp 1679235063
transform 1 0 21160 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1679235063
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1679235063
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1679235063
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1679235063
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1679235063
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1679235063
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1679235063
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1679235063
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1679235063
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1679235063
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_180
timestamp 1679235063
transform 1 0 17664 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1679235063
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1679235063
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_198
timestamp 1679235063
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_202
timestamp 1679235063
transform 1 0 19688 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1679235063
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1679235063
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1679235063
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1679235063
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1679235063
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1679235063
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1679235063
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1679235063
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1679235063
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_173
timestamp 1679235063
transform 1 0 17020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1679235063
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1679235063
transform 1 0 18308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1679235063
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1679235063
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1679235063
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_241
timestamp 1679235063
transform 1 0 23276 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_245
timestamp 1679235063
transform 1 0 23644 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1679235063
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1679235063
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1679235063
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1679235063
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1679235063
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1679235063
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1679235063
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1679235063
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_180
timestamp 1679235063
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1679235063
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1679235063
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_201
timestamp 1679235063
transform 1 0 19596 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_209
timestamp 1679235063
transform 1 0 20332 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1679235063
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1679235063
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1679235063
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1679235063
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1679235063
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1679235063
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1679235063
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1679235063
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1679235063
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1679235063
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1679235063
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_205
timestamp 1679235063
transform 1 0 19964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1679235063
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1679235063
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_233
timestamp 1679235063
transform 1 0 22540 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1679235063
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1679235063
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1679235063
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1679235063
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1679235063
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1679235063
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1679235063
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_151
timestamp 1679235063
transform 1 0 14996 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1679235063
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1679235063
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_171
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1679235063
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_198
timestamp 1679235063
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_219
timestamp 1679235063
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1679235063
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1679235063
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1679235063
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1679235063
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_121
timestamp 1679235063
transform 1 0 12236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_127
timestamp 1679235063
transform 1 0 12788 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1679235063
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1679235063
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1679235063
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1679235063
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1679235063
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_263
timestamp 1679235063
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1679235063
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1679235063
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1679235063
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1679235063
transform 1 0 10764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1679235063
transform 1 0 11132 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_119
timestamp 1679235063
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1679235063
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1679235063
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1679235063
transform 1 0 14812 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_153
timestamp 1679235063
transform 1 0 15180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1679235063
transform 1 0 15732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1679235063
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1679235063
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1679235063
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1679235063
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1679235063
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_259
timestamp 1679235063
transform 1 0 24932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1679235063
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1679235063
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1679235063
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1679235063
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1679235063
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1679235063
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1679235063
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1679235063
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1679235063
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_199
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1679235063
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_246
timestamp 1679235063
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_264
timestamp 1679235063
transform 1 0 25392 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1679235063
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1679235063
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1679235063
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1679235063
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1679235063
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1679235063
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1679235063
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_93
timestamp 1679235063
transform 1 0 9660 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_99
timestamp 1679235063
transform 1 0 10212 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1679235063
transform 1 0 10488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1679235063
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_119
timestamp 1679235063
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1679235063
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1679235063
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_135
timestamp 1679235063
transform 1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1679235063
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_161
timestamp 1679235063
transform 1 0 15916 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1679235063
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1679235063
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_210
timestamp 1679235063
transform 1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_231
timestamp 1679235063
transform 1 0 22356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_235
timestamp 1679235063
transform 1 0 22724 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1679235063
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1679235063
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1679235063
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1679235063
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_100
timestamp 1679235063
transform 1 0 10304 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1679235063
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1679235063
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1679235063
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1679235063
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1679235063
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1679235063
transform 1 0 22632 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_238
timestamp 1679235063
transform 1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_263
timestamp 1679235063
transform 1 0 25300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1679235063
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_27
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_33
timestamp 1679235063
transform 1 0 4140 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_36
timestamp 1679235063
transform 1 0 4416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_48
timestamp 1679235063
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1679235063
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_64
timestamp 1679235063
transform 1 0 6992 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_76
timestamp 1679235063
transform 1 0 8096 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_88
timestamp 1679235063
transform 1 0 9200 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1679235063
transform 1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1679235063
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1679235063
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_154
timestamp 1679235063
transform 1 0 15272 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1679235063
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_195
timestamp 1679235063
transform 1 0 19044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1679235063
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1679235063
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_235
timestamp 1679235063
transform 1 0 22724 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1679235063
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1679235063
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_14
timestamp 1679235063
transform 1 0 2392 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1679235063
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1679235063
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1679235063
transform 1 0 4968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_49
timestamp 1679235063
transform 1 0 5612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_62
timestamp 1679235063
transform 1 0 6808 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_69
timestamp 1679235063
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_91
timestamp 1679235063
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1679235063
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1679235063
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_135
timestamp 1679235063
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1679235063
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_169
timestamp 1679235063
transform 1 0 16652 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1679235063
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1679235063
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1679235063
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_246
timestamp 1679235063
transform 1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_264
timestamp 1679235063
transform 1 0 25392 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1679235063
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_19
timestamp 1679235063
transform 1 0 2852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1679235063
transform 1 0 3496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_33
timestamp 1679235063
transform 1 0 4140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_40
timestamp 1679235063
transform 1 0 4784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1679235063
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1679235063
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1679235063
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_90
timestamp 1679235063
transform 1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1679235063
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1679235063
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1679235063
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1679235063
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1679235063
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_171
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1679235063
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1679235063
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1679235063
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1679235063
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_263
timestamp 1679235063
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1679235063
transform 1 0 2208 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_19
timestamp 1679235063
transform 1 0 2852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_31
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1679235063
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1679235063
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_58
timestamp 1679235063
transform 1 0 6440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1679235063
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1679235063
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1679235063
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1679235063
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1679235063
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1679235063
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1679235063
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1679235063
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1679235063
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1679235063
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1679235063
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1679235063
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1679235063
transform 1 0 1840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 1679235063
transform 1 0 2392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_19
timestamp 1679235063
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1679235063
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_47
timestamp 1679235063
transform 1 0 5428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1679235063
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1679235063
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1679235063
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1679235063
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1679235063
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1679235063
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1679235063
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1679235063
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1679235063
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1679235063
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1679235063
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1679235063
transform 1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_184
timestamp 1679235063
transform 1 0 18032 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1679235063
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_219
timestamp 1679235063
transform 1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1679235063
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1679235063
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1679235063
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_261
timestamp 1679235063
transform 1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1679235063
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_12
timestamp 1679235063
transform 1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 1679235063
transform 1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_35
timestamp 1679235063
transform 1 0 4324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1679235063
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1679235063
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1679235063
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1679235063
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1679235063
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1679235063
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1679235063
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1679235063
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1679235063
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_187
timestamp 1679235063
transform 1 0 18308 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_192
timestamp 1679235063
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1679235063
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1679235063
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_233
timestamp 1679235063
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_239
timestamp 1679235063
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1679235063
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1679235063
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_12
timestamp 1679235063
transform 1 0 2208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1679235063
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_26
timestamp 1679235063
transform 1 0 3496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1679235063
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1679235063
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_59
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1679235063
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_67
timestamp 1679235063
transform 1 0 7268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_74
timestamp 1679235063
transform 1 0 7912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1679235063
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1679235063
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1679235063
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1679235063
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1679235063
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1679235063
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1679235063
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_219
timestamp 1679235063
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_247
timestamp 1679235063
transform 1 0 23828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_253
timestamp 1679235063
transform 1 0 24380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1679235063
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_9
timestamp 1679235063
transform 1 0 1932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_13
timestamp 1679235063
transform 1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1679235063
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_47
timestamp 1679235063
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1679235063
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1679235063
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1679235063
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1679235063
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1679235063
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1679235063
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1679235063
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1679235063
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1679235063
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1679235063
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1679235063
transform 1 0 19780 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_207
timestamp 1679235063
transform 1 0 20148 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1679235063
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1679235063
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_5
timestamp 1679235063
transform 1 0 1564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1679235063
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_27
timestamp 1679235063
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_33
timestamp 1679235063
transform 1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1679235063
transform 1 0 4784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1679235063
transform 1 0 6808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_66
timestamp 1679235063
transform 1 0 7176 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_70
timestamp 1679235063
transform 1 0 7544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1679235063
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1679235063
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_117
timestamp 1679235063
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1679235063
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1679235063
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1679235063
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1679235063
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1679235063
transform 1 0 20056 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_219
timestamp 1679235063
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1679235063
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1679235063
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1679235063
transform 1 0 25116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1679235063
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_8
timestamp 1679235063
transform 1 0 1840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1679235063
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_48
timestamp 1679235063
transform 1 0 5520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_52
timestamp 1679235063
transform 1 0 5888 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_56
timestamp 1679235063
transform 1 0 6256 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1679235063
transform 1 0 6900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1679235063
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_87
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1679235063
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1679235063
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1679235063
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1679235063
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1679235063
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1679235063
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_175
timestamp 1679235063
transform 1 0 17204 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1679235063
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1679235063
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1679235063
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1679235063
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_214
timestamp 1679235063
transform 1 0 20792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1679235063
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1679235063
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1679235063
transform 1 0 1932 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_17
timestamp 1679235063
transform 1 0 2668 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_35
timestamp 1679235063
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_43
timestamp 1679235063
transform 1 0 5060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_47
timestamp 1679235063
transform 1 0 5428 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_51
timestamp 1679235063
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_60
timestamp 1679235063
transform 1 0 6624 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_70
timestamp 1679235063
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1679235063
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1679235063
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1679235063
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_128
timestamp 1679235063
transform 1 0 12880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1679235063
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_155
timestamp 1679235063
transform 1 0 15364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_159
timestamp 1679235063
transform 1 0 15732 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1679235063
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1679235063
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1679235063
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_217
timestamp 1679235063
transform 1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1679235063
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1679235063
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_241
timestamp 1679235063
transform 1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1679235063
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_8
timestamp 1679235063
transform 1 0 1840 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_59
timestamp 1679235063
transform 1 0 6532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_79
timestamp 1679235063
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_91
timestamp 1679235063
transform 1 0 9476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_95
timestamp 1679235063
transform 1 0 9844 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1679235063
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1679235063
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1679235063
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1679235063
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1679235063
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1679235063
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_191
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1679235063
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1679235063
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_232
timestamp 1679235063
transform 1 0 22448 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_244
timestamp 1679235063
transform 1 0 23552 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1679235063
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_9
timestamp 1679235063
transform 1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_16
timestamp 1679235063
transform 1 0 2576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1679235063
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1679235063
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1679235063
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1679235063
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_119
timestamp 1679235063
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_130
timestamp 1679235063
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1679235063
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1679235063
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_160
timestamp 1679235063
transform 1 0 15824 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_171
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1679235063
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_206
timestamp 1679235063
transform 1 0 20056 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1679235063
transform 1 0 21252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1679235063
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_8
timestamp 1679235063
transform 1 0 1840 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1679235063
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1679235063
transform 1 0 4048 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_42
timestamp 1679235063
transform 1 0 4968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_90
timestamp 1679235063
transform 1 0 9384 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1679235063
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_124
timestamp 1679235063
transform 1 0 12512 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_128
timestamp 1679235063
transform 1 0 12880 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1679235063
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1679235063
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_189
timestamp 1679235063
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1679235063
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1679235063
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1679235063
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1679235063
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_233
timestamp 1679235063
transform 1 0 22540 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1679235063
transform 1 0 2392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_59
timestamp 1679235063
transform 1 0 6532 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_66
timestamp 1679235063
transform 1 0 7176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1679235063
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1679235063
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1679235063
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1679235063
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1679235063
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_199
timestamp 1679235063
transform 1 0 19412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_203
timestamp 1679235063
transform 1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_215
timestamp 1679235063
transform 1 0 20884 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1679235063
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1679235063
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_261
timestamp 1679235063
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1679235063
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_8
timestamp 1679235063
transform 1 0 1840 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1679235063
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1679235063
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1679235063
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1679235063
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_131
timestamp 1679235063
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1679235063
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1679235063
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1679235063
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_192
timestamp 1679235063
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1679235063
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1679235063
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_60
timestamp 1679235063
transform 1 0 6624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1679235063
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_117
timestamp 1679235063
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_135
timestamp 1679235063
transform 1 0 13524 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_150
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_154
timestamp 1679235063
transform 1 0 15272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1679235063
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1679235063
transform 1 0 19872 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1679235063
transform 1 0 20424 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_227
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_250
timestamp 1679235063
transform 1 0 24104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_257
timestamp 1679235063
transform 1 0 24748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1679235063
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1679235063
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1679235063
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1679235063
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1679235063
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_227
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  hold2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20056 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  hold3
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14536 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold5
timestamp 1679235063
transform 1 0 7268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  hold6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22632 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold7
timestamp 1679235063
transform 1 0 21344 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold10
timestamp 1679235063
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold11
timestamp 1679235063
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold12
timestamp 1679235063
transform 1 0 24564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold13
timestamp 1679235063
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold14
timestamp 1679235063
transform 1 0 23000 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold15
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold16
timestamp 1679235063
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold17
timestamp 1679235063
transform 1 0 20516 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold18
timestamp 1679235063
transform 1 0 14352 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold19
timestamp 1679235063
transform 1 0 21896 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold20
timestamp 1679235063
transform 1 0 14352 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold21
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold22
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 9568 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold24
timestamp 1679235063
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 6808 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold26
timestamp 1679235063
transform 1 0 24656 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 1656 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 4232 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold29
timestamp 1679235063
transform 1 0 24196 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold30
timestamp 1679235063
transform 1 0 6808 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold31
timestamp 1679235063
transform 1 0 7912 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold32
timestamp 1679235063
transform 1 0 5796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold33
timestamp 1679235063
transform 1 0 1656 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold34
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold35
timestamp 1679235063
transform 1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold36
timestamp 1679235063
transform 1 0 9292 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 6808 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 7176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 12880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1679235063
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1679235063
transform 1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1679235063
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1679235063
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1679235063
transform 1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1679235063
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 16100 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 1564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 3864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1679235063
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1679235063
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 4692 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1679235063
transform 1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1679235063
transform 1 0 7636 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1679235063
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1679235063
transform 1 0 2576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 9752 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1679235063
transform 1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1679235063
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 19412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1679235063
transform 1 0 6532 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 7820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input62
timestamp 1679235063
transform 1 0 20056 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1679235063
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1679235063
transform 1 0 20608 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1679235063
transform 1 0 23736 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1679235063
transform 1 0 4692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1679235063
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1679235063
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1679235063
transform 1 0 20056 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1679235063
transform 1 0 22080 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1679235063
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1679235063
transform 1 0 22632 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1679235063
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1679235063
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1679235063
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 22080 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 1748 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 7176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 9844 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 11684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 12052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 2852 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 2760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 2024 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14904 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17020 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21620 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23276 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23276 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22540 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20700 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22816 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21896 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18308 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21344 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15456 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18032 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14996 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13616 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11592 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10672 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9016 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9016 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8924 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9200 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10488 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10672 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11776 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13708 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20424 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_0.mux_l1_in_1__159 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_2.mux_l2_in_0__165
timestamp 1679235063
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_4.mux_l2_in_0__134
timestamp 1679235063
transform 1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_6.mux_l1_in_1__139
timestamp 1679235063
transform 1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_8.mux_l2_in_0__140
timestamp 1679235063
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_10.mux_l2_in_0__160
timestamp 1679235063
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21620 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_12.mux_l2_in_0__161
timestamp 1679235063
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_14.mux_l2_in_0__162
timestamp 1679235063
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_16.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_18.mux_l2_in_0__164
timestamp 1679235063
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_28.mux_l2_in_0__166
timestamp 1679235063
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_30.mux_l2_in_0__167
timestamp 1679235063
transform 1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_32.mux_l2_in_0__132
timestamp 1679235063
transform 1 0 20516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18768 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_34.mux_l2_in_0__133
timestamp 1679235063
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_44.mux_l2_in_0__135
timestamp 1679235063
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_46.mux_l2_in_0__136
timestamp 1679235063
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_48.mux_l2_in_0__137
timestamp 1679235063
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_50.mux_l2_in_0__138
timestamp 1679235063
transform 1 0 20056 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_0.mux_l1_in_1__141
timestamp 1679235063
transform 1 0 21620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_2.mux_l2_in_0__147
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17848 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_4.mux_l2_in_0__152
timestamp 1679235063
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14352 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_6.mux_l1_in_1__157
timestamp 1679235063
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17204 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14076 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_8.mux_l2_in_0__158
timestamp 1679235063
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13800 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_10.mux_l2_in_0__142
timestamp 1679235063
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_12.mux_l2_in_0__143
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_14.mux_l2_in_0__144
timestamp 1679235063
transform 1 0 4508 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15456 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_16.mux_l2_in_0__145
timestamp 1679235063
transform 1 0 5336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_18.mux_l2_in_0__146
timestamp 1679235063
transform 1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_28.mux_l2_in_0__148
timestamp 1679235063
transform 1 0 5980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2576 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_30.mux_l2_in_0__149
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_32.mux_l2_in_0__150
timestamp 1679235063
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15456 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_34.mux_l2_in_0__151
timestamp 1679235063
transform 1 0 7268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10764 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_44.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_46.mux_l2_in_0__154
timestamp 1679235063
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_48.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17112 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_50.mux_l2_in_0__156
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 26200 280 27000 400 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 26200 17416 27000 17536 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 26200 18232 27000 18352 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 26200 19048 27000 19168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 26200 20680 27000 20800 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 26200 13336 27000 13456 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 16 nsew signal input
flabel metal3 s 26200 21496 27000 21616 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 17 nsew signal input
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 18 nsew signal input
flabel metal3 s 26200 22312 27000 22432 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 19 nsew signal input
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 20 nsew signal input
flabel metal3 s 26200 23128 27000 23248 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 21 nsew signal input
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 22 nsew signal input
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 23 nsew signal input
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 24 nsew signal input
flabel metal3 s 26200 24760 27000 24880 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 25 nsew signal input
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 26 nsew signal input
flabel metal3 s 26200 14152 27000 14272 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 27 nsew signal input
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 28 nsew signal input
flabel metal3 s 26200 14968 27000 15088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 29 nsew signal input
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 30 nsew signal input
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 31 nsew signal input
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 32 nsew signal input
flabel metal3 s 26200 16600 27000 16720 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 33 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 34 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 35 nsew signal tristate
flabel metal3 s 26200 5176 27000 5296 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 36 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 37 nsew signal tristate
flabel metal3 s 26200 5992 27000 6112 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 38 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 39 nsew signal tristate
flabel metal3 s 26200 6808 27000 6928 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 40 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 41 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 42 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 43 nsew signal tristate
flabel metal3 s 26200 8440 27000 8560 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 44 nsew signal tristate
flabel metal3 s 26200 1096 27000 1216 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 45 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 46 nsew signal tristate
flabel metal3 s 26200 9256 27000 9376 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 47 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 48 nsew signal tristate
flabel metal3 s 26200 10072 27000 10192 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 49 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 50 nsew signal tristate
flabel metal3 s 26200 10888 27000 11008 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 51 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 52 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 53 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 54 nsew signal tristate
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 55 nsew signal tristate
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 56 nsew signal tristate
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 57 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 58 nsew signal tristate
flabel metal3 s 26200 2728 27000 2848 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 59 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 60 nsew signal tristate
flabel metal3 s 26200 3544 27000 3664 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 61 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 62 nsew signal tristate
flabel metal3 s 26200 4360 27000 4480 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 63 nsew signal tristate
flabel metal2 s 12714 26200 12770 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 64 nsew signal input
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 65 nsew signal input
flabel metal2 s 16762 26200 16818 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 66 nsew signal input
flabel metal2 s 17130 26200 17186 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 67 nsew signal input
flabel metal2 s 17498 26200 17554 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 68 nsew signal input
flabel metal2 s 17866 26200 17922 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 69 nsew signal input
flabel metal2 s 18234 26200 18290 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 70 nsew signal input
flabel metal2 s 18602 26200 18658 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 71 nsew signal input
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 72 nsew signal input
flabel metal2 s 19338 26200 19394 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 73 nsew signal input
flabel metal2 s 19706 26200 19762 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 74 nsew signal input
flabel metal2 s 13082 26200 13138 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 75 nsew signal input
flabel metal2 s 20074 26200 20130 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 76 nsew signal input
flabel metal2 s 20442 26200 20498 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 77 nsew signal input
flabel metal2 s 20810 26200 20866 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 78 nsew signal input
flabel metal2 s 21178 26200 21234 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 79 nsew signal input
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 80 nsew signal input
flabel metal2 s 21914 26200 21970 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 81 nsew signal input
flabel metal2 s 22282 26200 22338 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 82 nsew signal input
flabel metal2 s 22650 26200 22706 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 83 nsew signal input
flabel metal2 s 23018 26200 23074 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 84 nsew signal input
flabel metal2 s 23386 26200 23442 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 85 nsew signal input
flabel metal2 s 13450 26200 13506 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 86 nsew signal input
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 87 nsew signal input
flabel metal2 s 14186 26200 14242 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 88 nsew signal input
flabel metal2 s 14554 26200 14610 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 89 nsew signal input
flabel metal2 s 14922 26200 14978 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 90 nsew signal input
flabel metal2 s 15290 26200 15346 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 91 nsew signal input
flabel metal2 s 15658 26200 15714 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 92 nsew signal input
flabel metal2 s 16026 26200 16082 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 93 nsew signal input
flabel metal2 s 1674 26200 1730 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 94 nsew signal tristate
flabel metal2 s 5354 26200 5410 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 95 nsew signal tristate
flabel metal2 s 5722 26200 5778 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 96 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 97 nsew signal tristate
flabel metal2 s 6458 26200 6514 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 98 nsew signal tristate
flabel metal2 s 6826 26200 6882 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 99 nsew signal tristate
flabel metal2 s 7194 26200 7250 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 100 nsew signal tristate
flabel metal2 s 7562 26200 7618 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 101 nsew signal tristate
flabel metal2 s 7930 26200 7986 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 102 nsew signal tristate
flabel metal2 s 8298 26200 8354 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 103 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 104 nsew signal tristate
flabel metal2 s 2042 26200 2098 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 105 nsew signal tristate
flabel metal2 s 9034 26200 9090 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 106 nsew signal tristate
flabel metal2 s 9402 26200 9458 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 107 nsew signal tristate
flabel metal2 s 9770 26200 9826 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 108 nsew signal tristate
flabel metal2 s 10138 26200 10194 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 109 nsew signal tristate
flabel metal2 s 10506 26200 10562 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 110 nsew signal tristate
flabel metal2 s 10874 26200 10930 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 111 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 112 nsew signal tristate
flabel metal2 s 11610 26200 11666 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 113 nsew signal tristate
flabel metal2 s 11978 26200 12034 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 114 nsew signal tristate
flabel metal2 s 12346 26200 12402 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 115 nsew signal tristate
flabel metal2 s 2410 26200 2466 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 116 nsew signal tristate
flabel metal2 s 2778 26200 2834 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 117 nsew signal tristate
flabel metal2 s 3146 26200 3202 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 118 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 119 nsew signal tristate
flabel metal2 s 3882 26200 3938 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 120 nsew signal tristate
flabel metal2 s 4250 26200 4306 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 121 nsew signal tristate
flabel metal2 s 4618 26200 4674 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 122 nsew signal tristate
flabel metal2 s 4986 26200 5042 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 123 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 prog_clk
port 124 nsew signal input
flabel metal2 s 24490 26200 24546 27000 0 FreeSans 224 90 0 0 prog_reset
port 125 nsew signal input
flabel metal2 s 24858 26200 24914 27000 0 FreeSans 224 90 0 0 reset
port 126 nsew signal input
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 26200 25576 27000 25696 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 26200 26392 27000 26512 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 25226 26200 25282 27000 0 FreeSans 224 90 0 0 test_enable
port 131 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
rlabel metal1 13478 23936 13478 23936 0 VGND
rlabel metal1 13478 24480 13478 24480 0 VPWR
rlabel metal1 6670 2822 6670 2822 0 ccff_head
rlabel metal3 24894 340 24894 340 0 ccff_tail
rlabel metal1 24656 11118 24656 11118 0 chanx_right_in[0]
rlabel metal1 24472 8058 24472 8058 0 chanx_right_in[10]
rlabel metal2 11362 18105 11362 18105 0 chanx_right_in[11]
rlabel metal2 13938 14127 13938 14127 0 chanx_right_in[12]
rlabel metal2 12834 18105 12834 18105 0 chanx_right_in[13]
rlabel metal1 19734 18870 19734 18870 0 chanx_right_in[14]
rlabel metal1 19550 19822 19550 19822 0 chanx_right_in[15]
rlabel metal1 23184 16082 23184 16082 0 chanx_right_in[16]
rlabel metal1 15640 17170 15640 17170 0 chanx_right_in[17]
rlabel metal2 22310 18819 22310 18819 0 chanx_right_in[18]
rlabel metal2 15042 19788 15042 19788 0 chanx_right_in[19]
rlabel metal1 21252 11118 21252 11118 0 chanx_right_in[1]
rlabel metal1 19918 8942 19918 8942 0 chanx_right_in[20]
rlabel metal1 21068 9554 21068 9554 0 chanx_right_in[21]
rlabel metal1 20884 9554 20884 9554 0 chanx_right_in[22]
rlabel metal3 22977 21420 22977 21420 0 chanx_right_in[23]
rlabel metal2 15870 11849 15870 11849 0 chanx_right_in[24]
rlabel metal1 15732 11118 15732 11118 0 chanx_right_in[25]
rlabel metal4 13524 19448 13524 19448 0 chanx_right_in[26]
rlabel metal2 16698 13396 16698 13396 0 chanx_right_in[27]
rlabel via2 10534 15011 10534 15011 0 chanx_right_in[28]
rlabel via2 16330 21403 16330 21403 0 chanx_right_in[29]
rlabel metal2 24610 10676 24610 10676 0 chanx_right_in[2]
rlabel metal1 22862 6732 22862 6732 0 chanx_right_in[3]
rlabel metal1 24748 14382 24748 14382 0 chanx_right_in[4]
rlabel metal2 17204 14450 17204 14450 0 chanx_right_in[5]
rlabel metal1 21022 8398 21022 8398 0 chanx_right_in[6]
rlabel metal1 25070 15470 25070 15470 0 chanx_right_in[7]
rlabel metal1 25576 6698 25576 6698 0 chanx_right_in[8]
rlabel metal1 23690 15674 23690 15674 0 chanx_right_in[9]
rlabel metal2 25070 1853 25070 1853 0 chanx_right_out[0]
rlabel metal1 24104 5270 24104 5270 0 chanx_right_out[10]
rlabel metal2 24794 4641 24794 4641 0 chanx_right_out[11]
rlabel metal3 25676 5644 25676 5644 0 chanx_right_out[12]
rlabel metal1 24104 6358 24104 6358 0 chanx_right_out[13]
rlabel metal2 24702 5797 24702 5797 0 chanx_right_out[14]
rlabel metal1 24426 6834 24426 6834 0 chanx_right_out[15]
rlabel metal1 24104 7446 24104 7446 0 chanx_right_out[16]
rlabel metal3 25584 7684 25584 7684 0 chanx_right_out[17]
rlabel metal1 24380 7922 24380 7922 0 chanx_right_out[18]
rlabel metal1 24104 8534 24104 8534 0 chanx_right_out[19]
rlabel metal3 24250 1156 24250 1156 0 chanx_right_out[1]
rlabel metal2 25162 8177 25162 8177 0 chanx_right_out[20]
rlabel metal1 24380 9010 24380 9010 0 chanx_right_out[21]
rlabel metal2 23322 9673 23322 9673 0 chanx_right_out[22]
rlabel metal2 24794 9265 24794 9265 0 chanx_right_out[23]
rlabel metal1 24104 10710 24104 10710 0 chanx_right_out[24]
rlabel metal2 24702 10217 24702 10217 0 chanx_right_out[25]
rlabel metal1 24380 11186 24380 11186 0 chanx_right_out[26]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[27]
rlabel metal2 24794 11373 24794 11373 0 chanx_right_out[28]
rlabel metal3 25768 12580 25768 12580 0 chanx_right_out[29]
rlabel metal2 22126 2805 22126 2805 0 chanx_right_out[2]
rlabel metal1 21114 2618 21114 2618 0 chanx_right_out[3]
rlabel metal3 25676 2380 25676 2380 0 chanx_right_out[4]
rlabel metal1 24104 3094 24104 3094 0 chanx_right_out[5]
rlabel metal3 25676 3196 25676 3196 0 chanx_right_out[6]
rlabel metal1 23322 4012 23322 4012 0 chanx_right_out[7]
rlabel metal2 25162 3553 25162 3553 0 chanx_right_out[8]
rlabel metal3 25676 4420 25676 4420 0 chanx_right_out[9]
rlabel via2 2162 17187 2162 17187 0 chany_top_in[0]
rlabel metal2 15226 24276 15226 24276 0 chany_top_in[10]
rlabel metal1 16146 14994 16146 14994 0 chany_top_in[11]
rlabel metal1 16054 22950 16054 22950 0 chany_top_in[12]
rlabel metal3 17089 23460 17089 23460 0 chany_top_in[13]
rlabel metal2 17894 25493 17894 25493 0 chany_top_in[14]
rlabel metal2 18814 24684 18814 24684 0 chany_top_in[15]
rlabel metal1 12650 22644 12650 22644 0 chany_top_in[16]
rlabel metal1 1840 22610 1840 22610 0 chany_top_in[17]
rlabel metal2 19366 24881 19366 24881 0 chany_top_in[18]
rlabel metal2 19734 24388 19734 24388 0 chany_top_in[19]
rlabel metal2 8878 19652 8878 19652 0 chany_top_in[1]
rlabel metal2 13662 23936 13662 23936 0 chany_top_in[20]
rlabel metal2 20470 26173 20470 26173 0 chany_top_in[21]
rlabel metal2 14122 23052 14122 23052 0 chany_top_in[22]
rlabel metal2 21206 26037 21206 26037 0 chany_top_in[23]
rlabel metal2 21298 26248 21298 26248 0 chany_top_in[24]
rlabel metal2 21942 26105 21942 26105 0 chany_top_in[25]
rlabel via2 2162 16099 2162 16099 0 chany_top_in[26]
rlabel metal3 17135 22100 17135 22100 0 chany_top_in[27]
rlabel metal1 25806 21862 25806 21862 0 chany_top_in[28]
rlabel metal1 16514 11118 16514 11118 0 chany_top_in[29]
rlabel metal2 13386 24803 13386 24803 0 chany_top_in[2]
rlabel metal2 13938 24735 13938 24735 0 chany_top_in[3]
rlabel metal1 1794 23698 1794 23698 0 chany_top_in[4]
rlabel metal2 14214 17884 14214 17884 0 chany_top_in[5]
rlabel metal2 7774 15963 7774 15963 0 chany_top_in[6]
rlabel metal2 15318 23385 15318 23385 0 chany_top_in[7]
rlabel metal2 15686 24609 15686 24609 0 chany_top_in[8]
rlabel metal1 16422 16626 16422 16626 0 chany_top_in[9]
rlabel metal1 2070 19278 2070 19278 0 chany_top_out[0]
rlabel metal1 4600 23766 4600 23766 0 chany_top_out[10]
rlabel metal2 5750 24490 5750 24490 0 chany_top_out[11]
rlabel metal2 6118 24184 6118 24184 0 chany_top_out[12]
rlabel metal1 4876 24242 4876 24242 0 chany_top_out[13]
rlabel metal1 7176 20978 7176 20978 0 chany_top_out[14]
rlabel metal1 7498 21454 7498 21454 0 chany_top_out[15]
rlabel metal1 6624 23766 6624 23766 0 chany_top_out[16]
rlabel metal1 7130 23018 7130 23018 0 chany_top_out[17]
rlabel metal2 8326 24184 8326 24184 0 chany_top_out[18]
rlabel metal1 7130 24106 7130 24106 0 chany_top_out[19]
rlabel metal2 2070 23028 2070 23028 0 chany_top_out[1]
rlabel metal2 8786 24497 8786 24497 0 chany_top_out[20]
rlabel metal1 8832 23086 8832 23086 0 chany_top_out[21]
rlabel metal1 8970 24242 8970 24242 0 chany_top_out[22]
rlabel metal1 9338 23766 9338 23766 0 chany_top_out[23]
rlabel metal2 10534 24728 10534 24728 0 chany_top_out[24]
rlabel metal2 10902 25034 10902 25034 0 chany_top_out[25]
rlabel metal1 11132 24242 11132 24242 0 chany_top_out[26]
rlabel metal1 12144 23154 12144 23154 0 chany_top_out[27]
rlabel metal2 12006 24966 12006 24966 0 chany_top_out[28]
rlabel metal2 12374 25272 12374 25272 0 chany_top_out[29]
rlabel metal2 2438 24252 2438 24252 0 chany_top_out[2]
rlabel metal1 3266 26418 3266 26418 0 chany_top_out[3]
rlabel metal2 3029 26316 3029 26316 0 chany_top_out[4]
rlabel metal2 3542 23878 3542 23878 0 chany_top_out[5]
rlabel metal1 4416 20978 4416 20978 0 chany_top_out[6]
rlabel metal1 4140 22678 4140 22678 0 chany_top_out[7]
rlabel metal1 3956 23018 3956 23018 0 chany_top_out[8]
rlabel metal2 5067 26316 5067 26316 0 chany_top_out[9]
rlabel metal1 21804 18326 21804 18326 0 clknet_0_prog_clk
rlabel metal1 10488 13158 10488 13158 0 clknet_3_0__leaf_prog_clk
rlabel metal1 15640 15538 15640 15538 0 clknet_3_1__leaf_prog_clk
rlabel metal2 9062 20978 9062 20978 0 clknet_3_2__leaf_prog_clk
rlabel metal1 14076 18394 14076 18394 0 clknet_3_3__leaf_prog_clk
rlabel metal1 19458 14042 19458 14042 0 clknet_3_4__leaf_prog_clk
rlabel metal1 20884 16626 20884 16626 0 clknet_3_5__leaf_prog_clk
rlabel metal1 19412 20910 19412 20910 0 clknet_3_6__leaf_prog_clk
rlabel metal1 23368 21522 23368 21522 0 clknet_3_7__leaf_prog_clk
rlabel metal2 7038 3604 7038 3604 0 net1
rlabel metal3 16054 15436 16054 15436 0 net10
rlabel metal2 24058 6494 24058 6494 0 net100
rlabel metal1 22862 4624 22862 4624 0 net101
rlabel metal2 18446 23902 18446 23902 0 net102
rlabel metal1 3588 23698 3588 23698 0 net103
rlabel metal1 13478 22984 13478 22984 0 net104
rlabel metal1 6026 17850 6026 17850 0 net105
rlabel metal1 4784 16626 4784 16626 0 net106
rlabel metal1 7452 17850 7452 17850 0 net107
rlabel metal1 7636 17306 7636 17306 0 net108
rlabel metal1 4830 23664 4830 23664 0 net109
rlabel metal2 19688 17238 19688 17238 0 net11
rlabel metal1 16100 17714 16100 17714 0 net110
rlabel metal2 16790 18887 16790 18887 0 net111
rlabel metal3 19665 21692 19665 21692 0 net112
rlabel metal1 2254 19856 2254 19856 0 net113
rlabel metal1 4094 17170 4094 17170 0 net114
rlabel metal1 4876 18802 4876 18802 0 net115
rlabel metal1 5382 16082 5382 16082 0 net116
rlabel metal1 6210 17238 6210 17238 0 net117
rlabel metal2 9476 20434 9476 20434 0 net118
rlabel metal1 3358 18802 3358 18802 0 net119
rlabel metal2 15318 19601 15318 19601 0 net12
rlabel metal1 6624 19414 6624 19414 0 net120
rlabel metal1 10856 23086 10856 23086 0 net121
rlabel metal2 5474 19897 5474 19897 0 net122
rlabel metal2 6394 19737 6394 19737 0 net123
rlabel metal1 2254 20944 2254 20944 0 net124
rlabel metal2 3082 20604 3082 20604 0 net125
rlabel metal1 2254 21964 2254 21964 0 net126
rlabel metal1 3174 21522 3174 21522 0 net127
rlabel metal1 4738 20026 4738 20026 0 net128
rlabel metal2 2898 18887 2898 18887 0 net129
rlabel metal2 12788 17748 12788 17748 0 net13
rlabel metal1 2300 23086 2300 23086 0 net130
rlabel metal4 19412 24344 19412 24344 0 net131
rlabel metal1 20470 10778 20470 10778 0 net132
rlabel metal1 19573 14382 19573 14382 0 net133
rlabel via2 1978 17731 1978 17731 0 net134
rlabel metal1 17664 13906 17664 13906 0 net135
rlabel metal2 19734 10761 19734 10761 0 net136
rlabel metal1 20608 12818 20608 12818 0 net137
rlabel metal2 24978 9486 24978 9486 0 net138
rlabel metal2 17572 12852 17572 12852 0 net139
rlabel via3 15893 20740 15893 20740 0 net14
rlabel metal1 13340 14246 13340 14246 0 net140
rlabel metal1 20930 16762 20930 16762 0 net141
rlabel metal1 15640 19346 15640 19346 0 net142
rlabel metal1 11822 21658 11822 21658 0 net143
rlabel metal1 5106 16218 5106 16218 0 net144
rlabel metal1 6624 15538 6624 15538 0 net145
rlabel metal1 10810 19856 10810 19856 0 net146
rlabel metal1 18354 20910 18354 20910 0 net147
rlabel metal1 9568 18666 9568 18666 0 net148
rlabel via2 12466 20587 12466 20587 0 net149
rlabel metal3 17687 20196 17687 20196 0 net15
rlabel metal1 10304 18394 10304 18394 0 net150
rlabel metal1 11132 16558 11132 16558 0 net151
rlabel metal1 14950 12818 14950 12818 0 net152
rlabel metal1 10580 16218 10580 16218 0 net153
rlabel metal1 13478 15470 13478 15470 0 net154
rlabel metal2 13570 15266 13570 15266 0 net155
rlabel metal1 13662 18666 13662 18666 0 net156
rlabel metal2 14766 23902 14766 23902 0 net157
rlabel metal1 14214 23698 14214 23698 0 net158
rlabel metal1 19872 19142 19872 19142 0 net159
rlabel via3 17733 18020 17733 18020 0 net16
rlabel metal1 20562 14552 20562 14552 0 net160
rlabel metal1 22425 11594 22425 11594 0 net161
rlabel metal1 20240 13838 20240 13838 0 net162
rlabel metal1 22494 6426 22494 6426 0 net163
rlabel metal1 24058 4454 24058 4454 0 net164
rlabel metal2 1978 14909 1978 14909 0 net165
rlabel metal1 21482 13906 21482 13906 0 net166
rlabel metal1 21022 15334 21022 15334 0 net167
rlabel metal2 14766 12954 14766 12954 0 net168
rlabel metal1 21712 22610 21712 22610 0 net169
rlabel metal3 17687 19380 17687 19380 0 net17
rlabel metal2 20194 11237 20194 11237 0 net170
rlabel metal1 16008 14926 16008 14926 0 net171
rlabel metal2 19458 23987 19458 23987 0 net172
rlabel metal1 2116 20774 2116 20774 0 net173
rlabel via2 22034 9027 22034 9027 0 net174
rlabel metal2 7222 2890 7222 2890 0 net175
rlabel metal1 9844 8874 9844 8874 0 net176
rlabel metal1 10787 11254 10787 11254 0 net177
rlabel metal2 14490 14586 14490 14586 0 net178
rlabel metal2 16238 14280 16238 14280 0 net179
rlabel metal2 18354 21250 18354 21250 0 net18
rlabel metal2 19182 11424 19182 11424 0 net180
rlabel via2 16790 12835 16790 12835 0 net181
rlabel metal1 25392 16558 25392 16558 0 net182
rlabel via2 16790 19805 16790 19805 0 net183
rlabel metal2 15686 14909 15686 14909 0 net184
rlabel metal1 14536 20774 14536 20774 0 net185
rlabel metal2 20746 14654 20746 14654 0 net186
rlabel metal2 11178 16014 11178 16014 0 net187
rlabel metal2 25254 10200 25254 10200 0 net188
rlabel metal2 25438 9282 25438 9282 0 net189
rlabel metal1 15180 11322 15180 11322 0 net19
rlabel metal1 7222 18224 7222 18224 0 net190
rlabel metal2 7866 18564 7866 18564 0 net191
rlabel metal1 6854 17170 6854 17170 0 net192
rlabel via2 16330 10659 16330 10659 0 net193
rlabel metal2 2714 20536 2714 20536 0 net194
rlabel metal1 4232 19890 4232 19890 0 net195
rlabel metal1 18998 12784 18998 12784 0 net196
rlabel metal2 5152 19924 5152 19924 0 net197
rlabel metal1 2806 17612 2806 17612 0 net198
rlabel metal1 4094 16116 4094 16116 0 net199
rlabel metal1 18906 19686 18906 19686 0 net2
rlabel via2 1794 21947 1794 21947 0 net20
rlabel metal1 2300 23494 2300 23494 0 net200
rlabel metal1 18906 11220 18906 11220 0 net201
rlabel metal1 8970 20502 8970 20502 0 net202
rlabel metal2 16514 17187 16514 17187 0 net203
rlabel metal2 7498 3332 7498 3332 0 net204
rlabel metal1 6831 2414 6831 2414 0 net205
rlabel metal1 8648 4794 8648 4794 0 net206
rlabel via2 2622 20349 2622 20349 0 net21
rlabel metal2 19366 19737 19366 19737 0 net22
rlabel metal1 18446 23018 18446 23018 0 net23
rlabel metal1 20562 7718 20562 7718 0 net24
rlabel metal1 17296 17578 17296 17578 0 net25
rlabel metal1 19274 16150 19274 16150 0 net26
rlabel metal1 17112 17170 17112 17170 0 net27
rlabel metal1 18124 9418 18124 9418 0 net28
rlabel metal2 13524 19108 13524 19108 0 net29
rlabel metal1 17066 8058 17066 8058 0 net3
rlabel metal2 22954 22814 22954 22814 0 net30
rlabel metal2 7176 21012 7176 21012 0 net31
rlabel metal1 1702 17306 1702 17306 0 net32
rlabel metal3 12420 14960 12420 14960 0 net33
rlabel metal2 21022 14195 21022 14195 0 net34
rlabel metal1 22310 11832 22310 11832 0 net35
rlabel metal2 19734 18241 19734 18241 0 net36
rlabel metal1 21712 16422 21712 16422 0 net37
rlabel metal1 21988 19142 21988 19142 0 net38
rlabel metal2 20930 18445 20930 18445 0 net39
rlabel metal2 8418 17408 8418 17408 0 net4
rlabel metal2 21298 10591 21298 10591 0 net40
rlabel via2 7682 18139 7682 18139 0 net41
rlabel metal1 13662 14008 13662 14008 0 net42
rlabel metal1 2668 17510 2668 17510 0 net43
rlabel metal2 3266 17561 3266 17561 0 net44
rlabel metal1 7084 17034 7084 17034 0 net45
rlabel metal3 12788 13736 12788 13736 0 net46
rlabel metal3 17204 19992 17204 19992 0 net47
rlabel metal2 21298 20043 21298 20043 0 net48
rlabel metal2 10258 20400 10258 20400 0 net49
rlabel metal1 13156 14042 13156 14042 0 net5
rlabel metal1 14214 24072 14214 24072 0 net50
rlabel metal1 17020 23766 17020 23766 0 net51
rlabel metal1 19550 9418 19550 9418 0 net52
rlabel metal1 16100 23766 16100 23766 0 net53
rlabel metal1 5704 15130 5704 15130 0 net54
rlabel metal1 25116 9146 25116 9146 0 net55
rlabel via1 6877 7514 6877 7514 0 net56
rlabel via2 21022 15997 21022 15997 0 net57
rlabel metal2 13386 13566 13386 13566 0 net58
rlabel metal1 17756 18802 17756 18802 0 net59
rlabel metal2 18814 18241 18814 18241 0 net6
rlabel metal2 15870 17357 15870 17357 0 net60
rlabel metal1 22954 9928 22954 9928 0 net61
rlabel metal2 20562 24446 20562 24446 0 net62
rlabel metal1 17250 21522 17250 21522 0 net63
rlabel metal2 20746 19023 20746 19023 0 net64
rlabel metal1 20930 17544 20930 17544 0 net65
rlabel metal1 20976 19482 20976 19482 0 net66
rlabel metal1 8694 20264 8694 20264 0 net67
rlabel metal1 17618 17170 17618 17170 0 net68
rlabel metal1 20700 16150 20700 16150 0 net69
rlabel metal2 14030 18054 14030 18054 0 net7
rlabel metal1 13110 20570 13110 20570 0 net70
rlabel metal1 20746 2414 20746 2414 0 net71
rlabel metal1 19504 3026 19504 3026 0 net72
rlabel metal1 22402 5202 22402 5202 0 net73
rlabel metal1 23966 4148 23966 4148 0 net74
rlabel metal1 23782 6630 23782 6630 0 net75
rlabel metal2 22034 7004 22034 7004 0 net76
rlabel metal1 22586 5236 22586 5236 0 net77
rlabel metal2 22678 6324 22678 6324 0 net78
rlabel metal2 21942 8942 21942 8942 0 net79
rlabel metal2 6578 17527 6578 17527 0 net8
rlabel metal1 25024 6290 25024 6290 0 net80
rlabel metal1 22678 7922 22678 7922 0 net81
rlabel metal1 22126 8534 22126 8534 0 net82
rlabel metal1 20332 3502 20332 3502 0 net83
rlabel metal1 23966 7344 23966 7344 0 net84
rlabel metal1 21390 5338 21390 5338 0 net85
rlabel metal1 22126 9588 22126 9588 0 net86
rlabel metal2 22218 8262 22218 8262 0 net87
rlabel metal2 22126 11526 22126 11526 0 net88
rlabel metal1 23966 9486 23966 9486 0 net89
rlabel metal2 12742 14212 12742 14212 0 net9
rlabel metal2 22678 10676 22678 10676 0 net90
rlabel metal2 22310 10064 22310 10064 0 net91
rlabel metal1 22218 10676 22218 10676 0 net92
rlabel metal1 23874 6766 23874 6766 0 net93
rlabel metal1 22218 4080 22218 4080 0 net94
rlabel metal1 25668 7786 25668 7786 0 net95
rlabel metal1 22862 2346 22862 2346 0 net96
rlabel metal2 22310 3196 22310 3196 0 net97
rlabel metal1 23782 3502 23782 3502 0 net98
rlabel metal1 22862 4114 22862 4114 0 net99
rlabel metal1 20056 14586 20056 14586 0 prog_clk
rlabel metal2 21390 8466 21390 8466 0 prog_reset
rlabel metal1 25530 5814 25530 5814 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 1794 23511 1794 23511 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 23966 20910 23966 20910 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 21390 22593 21390 22593 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 15410 17714 15410 17714 0 sb_0__0_.mem_right_track_0.ccff_head
rlabel metal2 19918 19822 19918 19822 0 sb_0__0_.mem_right_track_0.ccff_tail
rlabel metal2 17342 18394 17342 18394 0 sb_0__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 25254 19516 25254 19516 0 sb_0__0_.mem_right_track_10.ccff_head
rlabel metal1 23736 17714 23736 17714 0 sb_0__0_.mem_right_track_10.ccff_tail
rlabel metal1 25392 19482 25392 19482 0 sb_0__0_.mem_right_track_10.mem_out\[0\]
rlabel metal2 22218 16932 22218 16932 0 sb_0__0_.mem_right_track_12.ccff_tail
rlabel metal2 21666 19244 21666 19244 0 sb_0__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 23966 15572 23966 15572 0 sb_0__0_.mem_right_track_14.ccff_tail
rlabel metal1 22586 17850 22586 17850 0 sb_0__0_.mem_right_track_14.mem_out\[0\]
rlabel metal1 23460 12274 23460 12274 0 sb_0__0_.mem_right_track_16.ccff_tail
rlabel metal1 24702 15130 24702 15130 0 sb_0__0_.mem_right_track_16.mem_out\[0\]
rlabel metal1 23000 12954 23000 12954 0 sb_0__0_.mem_right_track_18.ccff_tail
rlabel metal1 23230 12410 23230 12410 0 sb_0__0_.mem_right_track_18.mem_out\[0\]
rlabel metal1 22264 21862 22264 21862 0 sb_0__0_.mem_right_track_2.ccff_tail
rlabel metal1 20746 20570 20746 20570 0 sb_0__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 21298 13804 21298 13804 0 sb_0__0_.mem_right_track_28.ccff_tail
rlabel metal1 20095 13498 20095 13498 0 sb_0__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 20194 16422 20194 16422 0 sb_0__0_.mem_right_track_30.ccff_tail
rlabel metal1 19957 16762 19957 16762 0 sb_0__0_.mem_right_track_30.mem_out\[0\]
rlabel metal1 18078 16422 18078 16422 0 sb_0__0_.mem_right_track_32.ccff_tail
rlabel metal1 20194 17306 20194 17306 0 sb_0__0_.mem_right_track_32.mem_out\[0\]
rlabel metal1 18492 14790 18492 14790 0 sb_0__0_.mem_right_track_34.ccff_tail
rlabel metal1 19320 15674 19320 15674 0 sb_0__0_.mem_right_track_34.mem_out\[0\]
rlabel metal1 25300 18190 25300 18190 0 sb_0__0_.mem_right_track_4.ccff_tail
rlabel metal2 22586 23460 22586 23460 0 sb_0__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 17296 13158 17296 13158 0 sb_0__0_.mem_right_track_44.ccff_tail
rlabel metal1 18400 14518 18400 14518 0 sb_0__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 19136 12682 19136 12682 0 sb_0__0_.mem_right_track_46.ccff_tail
rlabel metal1 17756 12750 17756 12750 0 sb_0__0_.mem_right_track_46.mem_out\[0\]
rlabel metal1 20746 12682 20746 12682 0 sb_0__0_.mem_right_track_48.ccff_tail
rlabel metal2 20102 15067 20102 15067 0 sb_0__0_.mem_right_track_48.mem_out\[0\]
rlabel metal1 21252 16014 21252 16014 0 sb_0__0_.mem_right_track_50.mem_out\[0\]
rlabel metal1 24288 21454 24288 21454 0 sb_0__0_.mem_right_track_6.ccff_tail
rlabel metal1 17572 23630 17572 23630 0 sb_0__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 24472 21318 24472 21318 0 sb_0__0_.mem_right_track_8.mem_out\[0\]
rlabel metal1 15916 18666 15916 18666 0 sb_0__0_.mem_top_track_0.ccff_tail
rlabel metal1 20332 19890 20332 19890 0 sb_0__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 15088 22746 15088 22746 0 sb_0__0_.mem_top_track_10.ccff_head
rlabel metal1 14398 20366 14398 20366 0 sb_0__0_.mem_top_track_10.ccff_tail
rlabel metal1 15088 21862 15088 21862 0 sb_0__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 12144 20978 12144 20978 0 sb_0__0_.mem_top_track_12.ccff_tail
rlabel metal2 14490 19720 14490 19720 0 sb_0__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 12374 22066 12374 22066 0 sb_0__0_.mem_top_track_14.ccff_tail
rlabel metal1 13248 21114 13248 21114 0 sb_0__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 10534 20672 10534 20672 0 sb_0__0_.mem_top_track_16.ccff_tail
rlabel metal1 11224 22406 11224 22406 0 sb_0__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 10028 19482 10028 19482 0 sb_0__0_.mem_top_track_18.ccff_tail
rlabel metal2 10810 20128 10810 20128 0 sb_0__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 19136 20978 19136 20978 0 sb_0__0_.mem_top_track_2.ccff_tail
rlabel metal1 18032 20366 18032 20366 0 sb_0__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 10074 17340 10074 17340 0 sb_0__0_.mem_top_track_28.ccff_tail
rlabel metal1 15778 18258 15778 18258 0 sb_0__0_.mem_top_track_28.mem_out\[0\]
rlabel via1 12650 17731 12650 17731 0 sb_0__0_.mem_top_track_30.ccff_tail
rlabel via2 12466 17493 12466 17493 0 sb_0__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 12374 17306 12374 17306 0 sb_0__0_.mem_top_track_32.ccff_tail
rlabel metal1 13754 17544 13754 17544 0 sb_0__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 11960 15334 11960 15334 0 sb_0__0_.mem_top_track_34.ccff_tail
rlabel metal1 13800 15878 13800 15878 0 sb_0__0_.mem_top_track_34.mem_out\[0\]
rlabel metal2 18354 23460 18354 23460 0 sb_0__0_.mem_top_track_4.ccff_tail
rlabel metal1 20470 23154 20470 23154 0 sb_0__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 12006 15402 12006 15402 0 sb_0__0_.mem_top_track_44.ccff_tail
rlabel metal1 12558 14450 12558 14450 0 sb_0__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 14398 13226 14398 13226 0 sb_0__0_.mem_top_track_46.ccff_tail
rlabel metal1 14720 13158 14720 13158 0 sb_0__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14582 15232 14582 15232 0 sb_0__0_.mem_top_track_48.ccff_tail
rlabel metal1 15035 13702 15035 13702 0 sb_0__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16376 14246 16376 14246 0 sb_0__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 16560 23154 16560 23154 0 sb_0__0_.mem_top_track_6.ccff_tail
rlabel metal2 19826 22814 19826 22814 0 sb_0__0_.mem_top_track_6.mem_out\[0\]
rlabel metal2 21022 22202 21022 22202 0 sb_0__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 21298 8092 21298 8092 0 sb_0__0_.mux_right_track_0.out
rlabel metal1 19182 19346 19182 19346 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 19482 20056 19482 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 19849 19380 19849 19380 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16238 10234 16238 10234 0 sb_0__0_.mux_right_track_10.out
rlabel metal1 23874 17646 23874 17646 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18538 12818 18538 12818 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19780 7854 19780 7854 0 sb_0__0_.mux_right_track_12.out
rlabel metal2 21942 18496 21942 18496 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18538 12784 18538 12784 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20700 7174 20700 7174 0 sb_0__0_.mux_right_track_14.out
rlabel metal2 23874 18224 23874 18224 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21620 7378 21620 7378 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20700 5202 20700 5202 0 sb_0__0_.mux_right_track_16.out
rlabel metal1 23644 14450 23644 14450 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 10132 21482 10132 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20838 8636 20838 8636 0 sb_0__0_.mux_right_track_18.out
rlabel metal1 25070 13396 25070 13396 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20838 10608 20838 10608 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9200 12206 9200 12206 0 sb_0__0_.mux_right_track_2.out
rlabel metal2 16468 21318 16468 21318 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4784 17646 4784 17646 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 5678 20746 5678 0 sb_0__0_.mux_right_track_28.out
rlabel metal1 20838 13974 20838 13974 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20792 8466 20792 8466 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20516 5814 20516 5814 0 sb_0__0_.mux_right_track_30.out
rlabel metal2 21206 17510 21206 17510 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22034 5678 22034 5678 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21666 8058 21666 8058 0 sb_0__0_.mux_right_track_32.out
rlabel metal1 20286 15470 20286 15470 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19274 8466 19274 8466 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24932 7140 24932 7140 0 sb_0__0_.mux_right_track_34.out
rlabel metal1 19596 14246 19596 14246 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21574 8330 21574 8330 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14168 17510 14168 17510 0 sb_0__0_.mux_right_track_4.out
rlabel via2 16974 24395 16974 24395 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20746 18003 20746 18003 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19642 7378 19642 7378 0 sb_0__0_.mux_right_track_44.out
rlabel metal2 17526 16048 17526 16048 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17756 12716 17756 12716 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23920 4590 23920 4590 0 sb_0__0_.mux_right_track_46.out
rlabel metal1 19228 12954 19228 12954 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20010 7786 20010 7786 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24886 3536 24886 3536 0 sb_0__0_.mux_right_track_48.out
rlabel metal1 20286 12954 20286 12954 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20332 12614 20332 12614 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 2414 24702 2414 0 sb_0__0_.mux_right_track_50.out
rlabel metal1 25024 10030 25024 10030 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23690 10166 23690 10166 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10603 10778 10603 10778 0 sb_0__0_.mux_right_track_6.out
rlabel metal2 24702 23936 24702 23936 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24794 17850 24794 17850 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 9062 16779 9062 16779 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17434 9452 17434 9452 0 sb_0__0_.mux_right_track_8.out
rlabel metal1 20056 18326 20056 18326 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17618 9503 17618 9503 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21298 24157 21298 24157 0 sb_0__0_.mux_top_track_0.out
rlabel metal2 14306 19176 14306 19176 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15410 19482 15410 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14766 19482 14766 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 5336 19210 5336 19210 0 sb_0__0_.mux_top_track_10.out
rlabel metal2 17710 21726 17710 21726 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13800 21658 13800 21658 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2622 16456 2622 16456 0 sb_0__0_.mux_top_track_12.out
rlabel metal2 16698 21386 16698 21386 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 2645 16626 2645 16626 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5290 16014 5290 16014 0 sb_0__0_.mux_top_track_14.out
rlabel metal1 15410 22066 15410 22066 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9522 17646 9522 17646 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8326 18530 8326 18530 0 sb_0__0_.mux_top_track_16.out
rlabel metal1 14168 21046 14168 21046 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8510 19652 8510 19652 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3312 17170 3312 17170 0 sb_0__0_.mux_top_track_18.out
rlabel metal1 11040 19754 11040 19754 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 3450 18190 3450 18190 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5106 17646 5106 17646 0 sb_0__0_.mux_top_track_2.out
rlabel metal2 20010 20723 20010 20723 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17572 21114 17572 21114 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 5566 16490 5566 16490 0 sb_0__0_.mux_top_track_28.out
rlabel metal1 14858 18394 14858 18394 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 3128 16082 3128 16082 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7038 16694 7038 16694 0 sb_0__0_.mux_top_track_30.out
rlabel metal1 16882 20026 16882 20026 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 6762 16388 6762 16388 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4554 16660 4554 16660 0 sb_0__0_.mux_top_track_32.out
rlabel metal1 12926 18088 12926 18088 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11040 18122 11040 18122 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6256 16762 6256 16762 0 sb_0__0_.mux_top_track_34.out
rlabel metal2 15134 16864 15134 16864 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6026 16524 6026 16524 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5336 15674 5336 15674 0 sb_0__0_.mux_top_track_4.out
rlabel metal1 19366 24174 19366 24174 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 15364 24072 15364 24072 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2806 18734 2806 18734 0 sb_0__0_.mux_top_track_44.out
rlabel metal1 14766 15946 14766 15946 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9844 15878 9844 15878 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6578 19652 6578 19652 0 sb_0__0_.mux_top_track_46.out
rlabel metal1 13202 15606 13202 15606 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11914 15657 11914 15657 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6670 20434 6670 20434 0 sb_0__0_.mux_top_track_48.out
rlabel metal1 16882 16218 16882 16218 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13202 15912 13202 15912 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1978 18360 1978 18360 0 sb_0__0_.mux_top_track_50.out
rlabel metal1 16100 17850 16100 17850 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7406 18904 7406 18904 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4232 16422 4232 16422 0 sb_0__0_.mux_top_track_6.out
rlabel metal1 14996 21318 14996 21318 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17250 23086 17250 23086 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 14996 16728 14996 16728 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 2622 17204 2622 17204 0 sb_0__0_.mux_top_track_8.out
rlabel metal1 19504 21658 19504 21658 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14122 23596 14122 23596 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 1702 21573 1702 21573 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1610 18734 1610 18734 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 2507 20570 2507 20570 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 1656 21590 1656 21590 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 27000
<< end >>
