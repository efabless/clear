* NGSPICE file created from fpga_core.ext - technology: sky130A

* Black-box entry subcircuit for cbx_1__1_ abstract view
.subckt cbx_1__1_ REGIN_FEEDTHROUGH REGOUT_FEEDTHROUGH SC_IN_BOT SC_IN_TOP SC_OUT_BOT
+ SC_OUT_TOP VGND VPWR bottom_grid_pin_0_ bottom_grid_pin_10_ bottom_grid_pin_11_
+ bottom_grid_pin_12_ bottom_grid_pin_13_ bottom_grid_pin_14_ bottom_grid_pin_15_
+ bottom_grid_pin_1_ bottom_grid_pin_2_ bottom_grid_pin_3_ bottom_grid_pin_4_ bottom_grid_pin_5_
+ bottom_grid_pin_6_ bottom_grid_pin_7_ bottom_grid_pin_8_ bottom_grid_pin_9_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] clk_1_N_out clk_1_S_out clk_1_W_in clk_2_E_out
+ clk_2_W_in clk_2_W_out clk_3_E_out clk_3_W_in clk_3_W_out prog_clk_0_N_in prog_clk_0_W_out
+ prog_clk_1_N_out prog_clk_1_S_out prog_clk_1_W_in prog_clk_2_E_out prog_clk_2_W_in
+ prog_clk_2_W_out prog_clk_3_E_out prog_clk_3_W_in prog_clk_3_W_out
.ends

* Black-box entry subcircuit for cby_1__1_ abstract view
.subckt cby_1__1_ Test_en_E_in Test_en_E_out Test_en_N_out Test_en_S_in Test_en_W_in
+ Test_en_W_out VGND VPWR ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9]
+ chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ clk_2_N_out clk_2_S_in clk_2_S_out clk_3_N_out clk_3_S_in clk_3_S_out left_grid_pin_16_
+ left_grid_pin_17_ left_grid_pin_18_ left_grid_pin_19_ left_grid_pin_20_ left_grid_pin_21_
+ left_grid_pin_22_ left_grid_pin_23_ left_grid_pin_24_ left_grid_pin_25_ left_grid_pin_26_
+ left_grid_pin_27_ left_grid_pin_28_ left_grid_pin_29_ left_grid_pin_30_ left_grid_pin_31_
+ prog_clk_0_N_out prog_clk_0_S_out prog_clk_0_W_in prog_clk_2_N_out prog_clk_2_S_in
+ prog_clk_2_S_out prog_clk_3_N_out prog_clk_3_S_in prog_clk_3_S_out
.ends

* Black-box entry subcircuit for sb_1__2_ abstract view
.subckt sb_1__2_ SC_IN_BOT SC_OUT_BOT VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ left_top_grid_pin_1_ prog_clk_0_S_in right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ right_top_grid_pin_1_
.ends

* Black-box entry subcircuit for grid_clb abstract view
.subckt grid_clb SC_IN_TOP SC_OUT_BOT SC_OUT_TOP Test_en_E_in Test_en_E_out Test_en_W_in
+ Test_en_W_out VGND VPWR bottom_width_0_height_0__pin_50_ bottom_width_0_height_0__pin_51_
+ ccff_head ccff_tail clk_0_N_in clk_0_S_in prog_clk_0_E_out prog_clk_0_N_in prog_clk_0_N_out
+ prog_clk_0_S_in prog_clk_0_S_out prog_clk_0_W_out right_width_0_height_0__pin_16_
+ right_width_0_height_0__pin_17_ right_width_0_height_0__pin_18_ right_width_0_height_0__pin_19_
+ right_width_0_height_0__pin_20_ right_width_0_height_0__pin_21_ right_width_0_height_0__pin_22_
+ right_width_0_height_0__pin_23_ right_width_0_height_0__pin_24_ right_width_0_height_0__pin_25_
+ right_width_0_height_0__pin_26_ right_width_0_height_0__pin_27_ right_width_0_height_0__pin_28_
+ right_width_0_height_0__pin_29_ right_width_0_height_0__pin_30_ right_width_0_height_0__pin_31_
+ right_width_0_height_0__pin_42_lower right_width_0_height_0__pin_42_upper right_width_0_height_0__pin_43_lower
+ right_width_0_height_0__pin_43_upper right_width_0_height_0__pin_44_lower right_width_0_height_0__pin_44_upper
+ right_width_0_height_0__pin_45_lower right_width_0_height_0__pin_45_upper right_width_0_height_0__pin_46_lower
+ right_width_0_height_0__pin_46_upper right_width_0_height_0__pin_47_lower right_width_0_height_0__pin_47_upper
+ right_width_0_height_0__pin_48_lower right_width_0_height_0__pin_48_upper right_width_0_height_0__pin_49_lower
+ right_width_0_height_0__pin_49_upper top_width_0_height_0__pin_0_ top_width_0_height_0__pin_10_
+ top_width_0_height_0__pin_11_ top_width_0_height_0__pin_12_ top_width_0_height_0__pin_13_
+ top_width_0_height_0__pin_14_ top_width_0_height_0__pin_15_ top_width_0_height_0__pin_1_
+ top_width_0_height_0__pin_2_ top_width_0_height_0__pin_32_ top_width_0_height_0__pin_33_
+ top_width_0_height_0__pin_34_lower top_width_0_height_0__pin_34_upper top_width_0_height_0__pin_35_lower
+ top_width_0_height_0__pin_35_upper top_width_0_height_0__pin_36_lower top_width_0_height_0__pin_36_upper
+ top_width_0_height_0__pin_37_lower top_width_0_height_0__pin_37_upper top_width_0_height_0__pin_38_lower
+ top_width_0_height_0__pin_38_upper top_width_0_height_0__pin_39_lower top_width_0_height_0__pin_39_upper
+ top_width_0_height_0__pin_3_ top_width_0_height_0__pin_40_lower top_width_0_height_0__pin_40_upper
+ top_width_0_height_0__pin_41_lower top_width_0_height_0__pin_41_upper top_width_0_height_0__pin_4_
+ top_width_0_height_0__pin_5_ top_width_0_height_0__pin_6_ top_width_0_height_0__pin_7_
+ top_width_0_height_0__pin_8_ top_width_0_height_0__pin_9_
.ends

* Black-box entry subcircuit for sb_1__0_ abstract view
.subckt sb_1__0_ SC_IN_TOP SC_OUT_TOP Test_en_N_out Test_en_S_in VGND VPWR ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11]
+ chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16]
+ chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11]
+ chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16]
+ chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] chany_top_out[9] clk_3_N_out clk_3_S_in left_bottom_grid_pin_11_
+ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ prog_clk_0_N_in prog_clk_3_N_out prog_clk_3_S_in right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_17_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_
+ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ top_left_grid_pin_42_
+ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_
+ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
.ends

* Black-box entry subcircuit for cby_2__1_ abstract view
.subckt cby_2__1_ IO_ISOL_N VGND VPWR ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9]
+ chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ left_grid_pin_16_ left_grid_pin_17_ left_grid_pin_18_ left_grid_pin_19_ left_grid_pin_20_
+ left_grid_pin_21_ left_grid_pin_22_ left_grid_pin_23_ left_grid_pin_24_ left_grid_pin_25_
+ left_grid_pin_26_ left_grid_pin_27_ left_grid_pin_28_ left_grid_pin_29_ left_grid_pin_30_
+ left_grid_pin_31_ left_width_0_height_0__pin_0_ left_width_0_height_0__pin_1_lower
+ left_width_0_height_0__pin_1_upper prog_clk_0_N_out prog_clk_0_S_out prog_clk_0_W_in
+ right_grid_pin_0_
.ends

* Black-box entry subcircuit for cbx_1__2_ abstract view
.subckt cbx_1__2_ IO_ISOL_N SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP VGND VPWR bottom_grid_pin_0_
+ bottom_grid_pin_10_ bottom_grid_pin_11_ bottom_grid_pin_12_ bottom_grid_pin_13_
+ bottom_grid_pin_14_ bottom_grid_pin_15_ bottom_grid_pin_1_ bottom_grid_pin_2_ bottom_grid_pin_3_
+ bottom_grid_pin_4_ bottom_grid_pin_5_ bottom_grid_pin_6_ bottom_grid_pin_7_ bottom_grid_pin_8_
+ bottom_grid_pin_9_ bottom_width_0_height_0__pin_0_ bottom_width_0_height_0__pin_1_lower
+ bottom_width_0_height_0__pin_1_upper ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ prog_clk_0_S_in prog_clk_0_W_out top_grid_pin_0_
.ends

* Black-box entry subcircuit for sb_1__1_ abstract view
.subckt sb_1__1_ Test_en_N_out Test_en_S_in VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] clk_1_E_out clk_1_N_in clk_1_W_out clk_2_E_out clk_2_N_in clk_2_N_out
+ clk_2_S_out clk_2_W_out clk_3_E_out clk_3_N_in clk_3_N_out clk_3_S_out clk_3_W_out
+ left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_ left_bottom_grid_pin_37_
+ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_ left_bottom_grid_pin_41_
+ prog_clk_0_N_in prog_clk_1_E_out prog_clk_1_N_in prog_clk_1_W_out prog_clk_2_E_out
+ prog_clk_2_N_in prog_clk_2_N_out prog_clk_2_S_out prog_clk_2_W_out prog_clk_3_E_out
+ prog_clk_3_N_in prog_clk_3_N_out prog_clk_3_S_out prog_clk_3_W_out right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ top_left_grid_pin_42_
+ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_
+ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
.ends

* Black-box entry subcircuit for cbx_1__0_ abstract view
.subckt cbx_1__0_ IO_ISOL_N SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP VGND VPWR bottom_grid_pin_0_
+ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_ bottom_grid_pin_16_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] prog_clk_0_N_in prog_clk_0_W_out top_width_0_height_0__pin_0_
+ top_width_0_height_0__pin_10_ top_width_0_height_0__pin_11_lower top_width_0_height_0__pin_11_upper
+ top_width_0_height_0__pin_12_ top_width_0_height_0__pin_13_lower top_width_0_height_0__pin_13_upper
+ top_width_0_height_0__pin_14_ top_width_0_height_0__pin_15_lower top_width_0_height_0__pin_15_upper
+ top_width_0_height_0__pin_16_ top_width_0_height_0__pin_17_lower top_width_0_height_0__pin_17_upper
+ top_width_0_height_0__pin_1_lower top_width_0_height_0__pin_1_upper top_width_0_height_0__pin_2_
+ top_width_0_height_0__pin_3_lower top_width_0_height_0__pin_3_upper top_width_0_height_0__pin_4_
+ top_width_0_height_0__pin_5_lower top_width_0_height_0__pin_5_upper top_width_0_height_0__pin_6_
+ top_width_0_height_0__pin_7_lower top_width_0_height_0__pin_7_upper top_width_0_height_0__pin_8_
+ top_width_0_height_0__pin_9_lower top_width_0_height_0__pin_9_upper
.ends

* Black-box entry subcircuit for sb_2__2_ abstract view
.subckt sb_2__2_ SC_IN_BOT SC_OUT_BOT VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ left_top_grid_pin_1_ prog_clk_0_S_in
.ends

* Black-box entry subcircuit for sb_2__1_ abstract view
.subckt sb_2__1_ VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_ bottom_left_grid_pin_44_
+ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_ bottom_left_grid_pin_48_
+ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ prog_clk_0_N_in top_left_grid_pin_42_ top_left_grid_pin_43_
+ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_ top_left_grid_pin_47_
+ top_left_grid_pin_48_ top_left_grid_pin_49_ top_right_grid_pin_1_
.ends

* Black-box entry subcircuit for sb_2__0_ abstract view
.subckt sb_2__0_ VGND VPWR ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_11_ left_bottom_grid_pin_13_
+ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_
+ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ prog_clk_0_N_in
+ top_left_grid_pin_42_ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_
+ top_left_grid_pin_46_ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
+ top_right_grid_pin_1_
.ends

* Black-box entry subcircuit for cby_0__1_ abstract view
.subckt cby_0__1_ IO_ISOL_N VGND VPWR ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9]
+ chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ left_grid_pin_0_ prog_clk_0_E_in right_width_0_height_0__pin_0_ right_width_0_height_0__pin_1_lower
+ right_width_0_height_0__pin_1_upper
.ends

* Black-box entry subcircuit for sb_0__2_ abstract view
.subckt sb_0__2_ SC_IN_TOP SC_OUT_BOT VGND VPWR bottom_left_grid_pin_1_ ccff_head
+ ccff_tail chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] prog_clk_0_E_in right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ right_top_grid_pin_1_
.ends

* Black-box entry subcircuit for sb_0__1_ abstract view
.subckt sb_0__1_ VGND VPWR bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk_0_E_in right_bottom_grid_pin_34_ right_bottom_grid_pin_35_
+ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_
+ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ top_left_grid_pin_1_
.ends

* Black-box entry subcircuit for tie_array abstract view
.subckt tie_array VGND VPWR x[0] x[1] x[2] x[3] x[4] x[5] x[6] x[7]
.ends

* Black-box entry subcircuit for sb_0__0_ abstract view
.subckt sb_0__0_ VGND VPWR ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9]
+ chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ prog_clk_0_E_in right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_
+ right_bottom_grid_pin_17_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ top_left_grid_pin_1_
.ends

.subckt fpga_core IO_ISOL_N Test_en VGND VPWR ccff_head ccff_tail clk gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9] prog_clk
+ sc_head sc_tail
Xcbx_5__6_ cbx_5__6_/REGIN_FEEDTHROUGH cbx_5__6_/REGOUT_FEEDTHROUGH cbx_5__6_/SC_IN_BOT
+ cbx_5__6_/SC_IN_TOP cbx_5__6_/SC_OUT_BOT cbx_5__6_/SC_OUT_TOP VGND VPWR cbx_5__6_/bottom_grid_pin_0_
+ cbx_5__6_/bottom_grid_pin_10_ cbx_5__6_/bottom_grid_pin_11_ cbx_5__6_/bottom_grid_pin_12_
+ cbx_5__6_/bottom_grid_pin_13_ cbx_5__6_/bottom_grid_pin_14_ cbx_5__6_/bottom_grid_pin_15_
+ cbx_5__6_/bottom_grid_pin_1_ cbx_5__6_/bottom_grid_pin_2_ cbx_5__6_/bottom_grid_pin_3_
+ cbx_5__6_/bottom_grid_pin_4_ cbx_5__6_/bottom_grid_pin_5_ cbx_5__6_/bottom_grid_pin_6_
+ cbx_5__6_/bottom_grid_pin_7_ cbx_5__6_/bottom_grid_pin_8_ cbx_5__6_/bottom_grid_pin_9_
+ sb_5__6_/ccff_tail sb_4__6_/ccff_head cbx_5__6_/chanx_left_in[0] cbx_5__6_/chanx_left_in[10]
+ cbx_5__6_/chanx_left_in[11] cbx_5__6_/chanx_left_in[12] cbx_5__6_/chanx_left_in[13]
+ cbx_5__6_/chanx_left_in[14] cbx_5__6_/chanx_left_in[15] cbx_5__6_/chanx_left_in[16]
+ cbx_5__6_/chanx_left_in[17] cbx_5__6_/chanx_left_in[18] cbx_5__6_/chanx_left_in[19]
+ cbx_5__6_/chanx_left_in[1] cbx_5__6_/chanx_left_in[2] cbx_5__6_/chanx_left_in[3]
+ cbx_5__6_/chanx_left_in[4] cbx_5__6_/chanx_left_in[5] cbx_5__6_/chanx_left_in[6]
+ cbx_5__6_/chanx_left_in[7] cbx_5__6_/chanx_left_in[8] cbx_5__6_/chanx_left_in[9]
+ sb_4__6_/chanx_right_in[0] sb_4__6_/chanx_right_in[10] sb_4__6_/chanx_right_in[11]
+ sb_4__6_/chanx_right_in[12] sb_4__6_/chanx_right_in[13] sb_4__6_/chanx_right_in[14]
+ sb_4__6_/chanx_right_in[15] sb_4__6_/chanx_right_in[16] sb_4__6_/chanx_right_in[17]
+ sb_4__6_/chanx_right_in[18] sb_4__6_/chanx_right_in[19] sb_4__6_/chanx_right_in[1]
+ sb_4__6_/chanx_right_in[2] sb_4__6_/chanx_right_in[3] sb_4__6_/chanx_right_in[4]
+ sb_4__6_/chanx_right_in[5] sb_4__6_/chanx_right_in[6] sb_4__6_/chanx_right_in[7]
+ sb_4__6_/chanx_right_in[8] sb_4__6_/chanx_right_in[9] sb_5__6_/chanx_left_out[0]
+ sb_5__6_/chanx_left_out[10] sb_5__6_/chanx_left_out[11] sb_5__6_/chanx_left_out[12]
+ sb_5__6_/chanx_left_out[13] sb_5__6_/chanx_left_out[14] sb_5__6_/chanx_left_out[15]
+ sb_5__6_/chanx_left_out[16] sb_5__6_/chanx_left_out[17] sb_5__6_/chanx_left_out[18]
+ sb_5__6_/chanx_left_out[19] sb_5__6_/chanx_left_out[1] sb_5__6_/chanx_left_out[2]
+ sb_5__6_/chanx_left_out[3] sb_5__6_/chanx_left_out[4] sb_5__6_/chanx_left_out[5]
+ sb_5__6_/chanx_left_out[6] sb_5__6_/chanx_left_out[7] sb_5__6_/chanx_left_out[8]
+ sb_5__6_/chanx_left_out[9] sb_5__6_/chanx_left_in[0] sb_5__6_/chanx_left_in[10]
+ sb_5__6_/chanx_left_in[11] sb_5__6_/chanx_left_in[12] sb_5__6_/chanx_left_in[13]
+ sb_5__6_/chanx_left_in[14] sb_5__6_/chanx_left_in[15] sb_5__6_/chanx_left_in[16]
+ sb_5__6_/chanx_left_in[17] sb_5__6_/chanx_left_in[18] sb_5__6_/chanx_left_in[19]
+ sb_5__6_/chanx_left_in[1] sb_5__6_/chanx_left_in[2] sb_5__6_/chanx_left_in[3] sb_5__6_/chanx_left_in[4]
+ sb_5__6_/chanx_left_in[5] sb_5__6_/chanx_left_in[6] sb_5__6_/chanx_left_in[7] sb_5__6_/chanx_left_in[8]
+ sb_5__6_/chanx_left_in[9] cbx_5__6_/clk_1_N_out cbx_5__6_/clk_1_S_out cbx_5__6_/clk_1_W_in
+ cbx_5__6_/clk_2_E_out cbx_5__6_/clk_2_W_in cbx_5__6_/clk_2_W_out cbx_5__6_/clk_3_E_out
+ cbx_5__6_/clk_3_W_in cbx_5__6_/clk_3_W_out cbx_5__6_/prog_clk_0_N_in cbx_5__6_/prog_clk_0_W_out
+ cbx_5__6_/prog_clk_1_N_out cbx_5__6_/prog_clk_1_S_out cbx_5__6_/prog_clk_1_W_in
+ cbx_5__6_/prog_clk_2_E_out cbx_5__6_/prog_clk_2_W_in cbx_5__6_/prog_clk_2_W_out
+ cbx_5__6_/prog_clk_3_E_out cbx_5__6_/prog_clk_3_W_in cbx_5__6_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_2__2_ cby_2__2_/Test_en_W_in cby_2__2_/Test_en_E_out cby_2__2_/Test_en_N_out
+ cby_2__2_/Test_en_W_in cby_2__2_/Test_en_W_in cby_2__2_/Test_en_W_out VGND VPWR
+ cby_2__2_/ccff_head cby_2__2_/ccff_tail sb_2__1_/chany_top_out[0] sb_2__1_/chany_top_out[10]
+ sb_2__1_/chany_top_out[11] sb_2__1_/chany_top_out[12] sb_2__1_/chany_top_out[13]
+ sb_2__1_/chany_top_out[14] sb_2__1_/chany_top_out[15] sb_2__1_/chany_top_out[16]
+ sb_2__1_/chany_top_out[17] sb_2__1_/chany_top_out[18] sb_2__1_/chany_top_out[19]
+ sb_2__1_/chany_top_out[1] sb_2__1_/chany_top_out[2] sb_2__1_/chany_top_out[3] sb_2__1_/chany_top_out[4]
+ sb_2__1_/chany_top_out[5] sb_2__1_/chany_top_out[6] sb_2__1_/chany_top_out[7] sb_2__1_/chany_top_out[8]
+ sb_2__1_/chany_top_out[9] sb_2__1_/chany_top_in[0] sb_2__1_/chany_top_in[10] sb_2__1_/chany_top_in[11]
+ sb_2__1_/chany_top_in[12] sb_2__1_/chany_top_in[13] sb_2__1_/chany_top_in[14] sb_2__1_/chany_top_in[15]
+ sb_2__1_/chany_top_in[16] sb_2__1_/chany_top_in[17] sb_2__1_/chany_top_in[18] sb_2__1_/chany_top_in[19]
+ sb_2__1_/chany_top_in[1] sb_2__1_/chany_top_in[2] sb_2__1_/chany_top_in[3] sb_2__1_/chany_top_in[4]
+ sb_2__1_/chany_top_in[5] sb_2__1_/chany_top_in[6] sb_2__1_/chany_top_in[7] sb_2__1_/chany_top_in[8]
+ sb_2__1_/chany_top_in[9] cby_2__2_/chany_top_in[0] cby_2__2_/chany_top_in[10] cby_2__2_/chany_top_in[11]
+ cby_2__2_/chany_top_in[12] cby_2__2_/chany_top_in[13] cby_2__2_/chany_top_in[14]
+ cby_2__2_/chany_top_in[15] cby_2__2_/chany_top_in[16] cby_2__2_/chany_top_in[17]
+ cby_2__2_/chany_top_in[18] cby_2__2_/chany_top_in[19] cby_2__2_/chany_top_in[1]
+ cby_2__2_/chany_top_in[2] cby_2__2_/chany_top_in[3] cby_2__2_/chany_top_in[4] cby_2__2_/chany_top_in[5]
+ cby_2__2_/chany_top_in[6] cby_2__2_/chany_top_in[7] cby_2__2_/chany_top_in[8] cby_2__2_/chany_top_in[9]
+ cby_2__2_/chany_top_out[0] cby_2__2_/chany_top_out[10] cby_2__2_/chany_top_out[11]
+ cby_2__2_/chany_top_out[12] cby_2__2_/chany_top_out[13] cby_2__2_/chany_top_out[14]
+ cby_2__2_/chany_top_out[15] cby_2__2_/chany_top_out[16] cby_2__2_/chany_top_out[17]
+ cby_2__2_/chany_top_out[18] cby_2__2_/chany_top_out[19] cby_2__2_/chany_top_out[1]
+ cby_2__2_/chany_top_out[2] cby_2__2_/chany_top_out[3] cby_2__2_/chany_top_out[4]
+ cby_2__2_/chany_top_out[5] cby_2__2_/chany_top_out[6] cby_2__2_/chany_top_out[7]
+ cby_2__2_/chany_top_out[8] cby_2__2_/chany_top_out[9] cby_2__2_/clk_2_N_out cby_2__2_/clk_2_S_in
+ cby_2__2_/clk_2_S_out cby_2__2_/clk_3_N_out cby_2__2_/clk_3_S_in cby_2__2_/clk_3_S_out
+ cby_2__2_/left_grid_pin_16_ cby_2__2_/left_grid_pin_17_ cby_2__2_/left_grid_pin_18_
+ cby_2__2_/left_grid_pin_19_ cby_2__2_/left_grid_pin_20_ cby_2__2_/left_grid_pin_21_
+ cby_2__2_/left_grid_pin_22_ cby_2__2_/left_grid_pin_23_ cby_2__2_/left_grid_pin_24_
+ cby_2__2_/left_grid_pin_25_ cby_2__2_/left_grid_pin_26_ cby_2__2_/left_grid_pin_27_
+ cby_2__2_/left_grid_pin_28_ cby_2__2_/left_grid_pin_29_ cby_2__2_/left_grid_pin_30_
+ cby_2__2_/left_grid_pin_31_ cby_2__2_/prog_clk_0_N_out sb_2__1_/prog_clk_0_N_in
+ cby_2__2_/prog_clk_0_W_in cby_2__2_/prog_clk_2_N_out cby_2__2_/prog_clk_2_S_in cby_2__2_/prog_clk_2_S_out
+ cby_2__2_/prog_clk_3_N_out cby_2__2_/prog_clk_3_S_in cby_2__2_/prog_clk_3_S_out
+ cby_1__1_
Xsb_2__8_ sb_2__8_/SC_IN_BOT sb_2__8_/SC_OUT_BOT VGND VPWR sb_2__8_/bottom_left_grid_pin_42_
+ sb_2__8_/bottom_left_grid_pin_43_ sb_2__8_/bottom_left_grid_pin_44_ sb_2__8_/bottom_left_grid_pin_45_
+ sb_2__8_/bottom_left_grid_pin_46_ sb_2__8_/bottom_left_grid_pin_47_ sb_2__8_/bottom_left_grid_pin_48_
+ sb_2__8_/bottom_left_grid_pin_49_ sb_2__8_/ccff_head sb_2__8_/ccff_tail sb_2__8_/chanx_left_in[0]
+ sb_2__8_/chanx_left_in[10] sb_2__8_/chanx_left_in[11] sb_2__8_/chanx_left_in[12]
+ sb_2__8_/chanx_left_in[13] sb_2__8_/chanx_left_in[14] sb_2__8_/chanx_left_in[15]
+ sb_2__8_/chanx_left_in[16] sb_2__8_/chanx_left_in[17] sb_2__8_/chanx_left_in[18]
+ sb_2__8_/chanx_left_in[19] sb_2__8_/chanx_left_in[1] sb_2__8_/chanx_left_in[2] sb_2__8_/chanx_left_in[3]
+ sb_2__8_/chanx_left_in[4] sb_2__8_/chanx_left_in[5] sb_2__8_/chanx_left_in[6] sb_2__8_/chanx_left_in[7]
+ sb_2__8_/chanx_left_in[8] sb_2__8_/chanx_left_in[9] sb_2__8_/chanx_left_out[0] sb_2__8_/chanx_left_out[10]
+ sb_2__8_/chanx_left_out[11] sb_2__8_/chanx_left_out[12] sb_2__8_/chanx_left_out[13]
+ sb_2__8_/chanx_left_out[14] sb_2__8_/chanx_left_out[15] sb_2__8_/chanx_left_out[16]
+ sb_2__8_/chanx_left_out[17] sb_2__8_/chanx_left_out[18] sb_2__8_/chanx_left_out[19]
+ sb_2__8_/chanx_left_out[1] sb_2__8_/chanx_left_out[2] sb_2__8_/chanx_left_out[3]
+ sb_2__8_/chanx_left_out[4] sb_2__8_/chanx_left_out[5] sb_2__8_/chanx_left_out[6]
+ sb_2__8_/chanx_left_out[7] sb_2__8_/chanx_left_out[8] sb_2__8_/chanx_left_out[9]
+ sb_2__8_/chanx_right_in[0] sb_2__8_/chanx_right_in[10] sb_2__8_/chanx_right_in[11]
+ sb_2__8_/chanx_right_in[12] sb_2__8_/chanx_right_in[13] sb_2__8_/chanx_right_in[14]
+ sb_2__8_/chanx_right_in[15] sb_2__8_/chanx_right_in[16] sb_2__8_/chanx_right_in[17]
+ sb_2__8_/chanx_right_in[18] sb_2__8_/chanx_right_in[19] sb_2__8_/chanx_right_in[1]
+ sb_2__8_/chanx_right_in[2] sb_2__8_/chanx_right_in[3] sb_2__8_/chanx_right_in[4]
+ sb_2__8_/chanx_right_in[5] sb_2__8_/chanx_right_in[6] sb_2__8_/chanx_right_in[7]
+ sb_2__8_/chanx_right_in[8] sb_2__8_/chanx_right_in[9] cbx_3__8_/chanx_left_in[0]
+ cbx_3__8_/chanx_left_in[10] cbx_3__8_/chanx_left_in[11] cbx_3__8_/chanx_left_in[12]
+ cbx_3__8_/chanx_left_in[13] cbx_3__8_/chanx_left_in[14] cbx_3__8_/chanx_left_in[15]
+ cbx_3__8_/chanx_left_in[16] cbx_3__8_/chanx_left_in[17] cbx_3__8_/chanx_left_in[18]
+ cbx_3__8_/chanx_left_in[19] cbx_3__8_/chanx_left_in[1] cbx_3__8_/chanx_left_in[2]
+ cbx_3__8_/chanx_left_in[3] cbx_3__8_/chanx_left_in[4] cbx_3__8_/chanx_left_in[5]
+ cbx_3__8_/chanx_left_in[6] cbx_3__8_/chanx_left_in[7] cbx_3__8_/chanx_left_in[8]
+ cbx_3__8_/chanx_left_in[9] cby_2__8_/chany_top_out[0] cby_2__8_/chany_top_out[10]
+ cby_2__8_/chany_top_out[11] cby_2__8_/chany_top_out[12] cby_2__8_/chany_top_out[13]
+ cby_2__8_/chany_top_out[14] cby_2__8_/chany_top_out[15] cby_2__8_/chany_top_out[16]
+ cby_2__8_/chany_top_out[17] cby_2__8_/chany_top_out[18] cby_2__8_/chany_top_out[19]
+ cby_2__8_/chany_top_out[1] cby_2__8_/chany_top_out[2] cby_2__8_/chany_top_out[3]
+ cby_2__8_/chany_top_out[4] cby_2__8_/chany_top_out[5] cby_2__8_/chany_top_out[6]
+ cby_2__8_/chany_top_out[7] cby_2__8_/chany_top_out[8] cby_2__8_/chany_top_out[9]
+ cby_2__8_/chany_top_in[0] cby_2__8_/chany_top_in[10] cby_2__8_/chany_top_in[11]
+ cby_2__8_/chany_top_in[12] cby_2__8_/chany_top_in[13] cby_2__8_/chany_top_in[14]
+ cby_2__8_/chany_top_in[15] cby_2__8_/chany_top_in[16] cby_2__8_/chany_top_in[17]
+ cby_2__8_/chany_top_in[18] cby_2__8_/chany_top_in[19] cby_2__8_/chany_top_in[1]
+ cby_2__8_/chany_top_in[2] cby_2__8_/chany_top_in[3] cby_2__8_/chany_top_in[4] cby_2__8_/chany_top_in[5]
+ cby_2__8_/chany_top_in[6] cby_2__8_/chany_top_in[7] cby_2__8_/chany_top_in[8] cby_2__8_/chany_top_in[9]
+ sb_2__8_/left_bottom_grid_pin_34_ sb_2__8_/left_bottom_grid_pin_35_ sb_2__8_/left_bottom_grid_pin_36_
+ sb_2__8_/left_bottom_grid_pin_37_ sb_2__8_/left_bottom_grid_pin_38_ sb_2__8_/left_bottom_grid_pin_39_
+ sb_2__8_/left_bottom_grid_pin_40_ sb_2__8_/left_bottom_grid_pin_41_ sb_2__8_/left_top_grid_pin_1_
+ sb_2__8_/prog_clk_0_S_in sb_2__8_/right_bottom_grid_pin_34_ sb_2__8_/right_bottom_grid_pin_35_
+ sb_2__8_/right_bottom_grid_pin_36_ sb_2__8_/right_bottom_grid_pin_37_ sb_2__8_/right_bottom_grid_pin_38_
+ sb_2__8_/right_bottom_grid_pin_39_ sb_2__8_/right_bottom_grid_pin_40_ sb_2__8_/right_bottom_grid_pin_41_
+ sb_2__8_/right_top_grid_pin_1_ sb_1__2_
Xgrid_clb_4__6_ cbx_4__5_/SC_OUT_TOP grid_clb_4__6_/SC_OUT_BOT cbx_4__6_/SC_IN_BOT
+ cby_4__6_/Test_en_W_out grid_clb_4__6_/Test_en_E_out cby_4__6_/Test_en_W_out cby_3__6_/Test_en_W_in
+ VGND VPWR cbx_4__5_/REGIN_FEEDTHROUGH grid_clb_4__6_/bottom_width_0_height_0__pin_51_
+ cby_3__6_/ccff_tail cby_4__6_/ccff_head cbx_4__5_/clk_1_N_out cbx_4__5_/clk_1_N_out
+ cby_4__6_/prog_clk_0_W_in cbx_4__5_/prog_clk_1_N_out grid_clb_4__6_/prog_clk_0_N_out
+ cbx_4__5_/prog_clk_1_N_out cbx_4__5_/prog_clk_0_N_in grid_clb_4__6_/prog_clk_0_W_out
+ cby_4__6_/left_grid_pin_16_ cby_4__6_/left_grid_pin_17_ cby_4__6_/left_grid_pin_18_
+ cby_4__6_/left_grid_pin_19_ cby_4__6_/left_grid_pin_20_ cby_4__6_/left_grid_pin_21_
+ cby_4__6_/left_grid_pin_22_ cby_4__6_/left_grid_pin_23_ cby_4__6_/left_grid_pin_24_
+ cby_4__6_/left_grid_pin_25_ cby_4__6_/left_grid_pin_26_ cby_4__6_/left_grid_pin_27_
+ cby_4__6_/left_grid_pin_28_ cby_4__6_/left_grid_pin_29_ cby_4__6_/left_grid_pin_30_
+ cby_4__6_/left_grid_pin_31_ sb_4__5_/top_left_grid_pin_42_ sb_4__6_/bottom_left_grid_pin_42_
+ sb_4__5_/top_left_grid_pin_43_ sb_4__6_/bottom_left_grid_pin_43_ sb_4__5_/top_left_grid_pin_44_
+ sb_4__6_/bottom_left_grid_pin_44_ sb_4__5_/top_left_grid_pin_45_ sb_4__6_/bottom_left_grid_pin_45_
+ sb_4__5_/top_left_grid_pin_46_ sb_4__6_/bottom_left_grid_pin_46_ sb_4__5_/top_left_grid_pin_47_
+ sb_4__6_/bottom_left_grid_pin_47_ sb_4__5_/top_left_grid_pin_48_ sb_4__6_/bottom_left_grid_pin_48_
+ sb_4__5_/top_left_grid_pin_49_ sb_4__6_/bottom_left_grid_pin_49_ cbx_4__6_/bottom_grid_pin_0_
+ cbx_4__6_/bottom_grid_pin_10_ cbx_4__6_/bottom_grid_pin_11_ cbx_4__6_/bottom_grid_pin_12_
+ cbx_4__6_/bottom_grid_pin_13_ cbx_4__6_/bottom_grid_pin_14_ cbx_4__6_/bottom_grid_pin_15_
+ cbx_4__6_/bottom_grid_pin_1_ cbx_4__6_/bottom_grid_pin_2_ cbx_4__6_/REGOUT_FEEDTHROUGH
+ grid_clb_4__6_/top_width_0_height_0__pin_33_ sb_4__6_/left_bottom_grid_pin_34_ sb_3__6_/right_bottom_grid_pin_34_
+ sb_4__6_/left_bottom_grid_pin_35_ sb_3__6_/right_bottom_grid_pin_35_ sb_4__6_/left_bottom_grid_pin_36_
+ sb_3__6_/right_bottom_grid_pin_36_ sb_4__6_/left_bottom_grid_pin_37_ sb_3__6_/right_bottom_grid_pin_37_
+ sb_4__6_/left_bottom_grid_pin_38_ sb_3__6_/right_bottom_grid_pin_38_ sb_4__6_/left_bottom_grid_pin_39_
+ sb_3__6_/right_bottom_grid_pin_39_ cbx_4__6_/bottom_grid_pin_3_ sb_4__6_/left_bottom_grid_pin_40_
+ sb_3__6_/right_bottom_grid_pin_40_ sb_4__6_/left_bottom_grid_pin_41_ sb_3__6_/right_bottom_grid_pin_41_
+ cbx_4__6_/bottom_grid_pin_4_ cbx_4__6_/bottom_grid_pin_5_ cbx_4__6_/bottom_grid_pin_6_
+ cbx_4__6_/bottom_grid_pin_7_ cbx_4__6_/bottom_grid_pin_8_ cbx_4__6_/bottom_grid_pin_9_
+ grid_clb
Xcbx_2__3_ cbx_2__3_/REGIN_FEEDTHROUGH cbx_2__3_/REGOUT_FEEDTHROUGH cbx_2__3_/SC_IN_BOT
+ cbx_2__3_/SC_IN_TOP cbx_2__3_/SC_OUT_BOT cbx_2__3_/SC_OUT_TOP VGND VPWR cbx_2__3_/bottom_grid_pin_0_
+ cbx_2__3_/bottom_grid_pin_10_ cbx_2__3_/bottom_grid_pin_11_ cbx_2__3_/bottom_grid_pin_12_
+ cbx_2__3_/bottom_grid_pin_13_ cbx_2__3_/bottom_grid_pin_14_ cbx_2__3_/bottom_grid_pin_15_
+ cbx_2__3_/bottom_grid_pin_1_ cbx_2__3_/bottom_grid_pin_2_ cbx_2__3_/bottom_grid_pin_3_
+ cbx_2__3_/bottom_grid_pin_4_ cbx_2__3_/bottom_grid_pin_5_ cbx_2__3_/bottom_grid_pin_6_
+ cbx_2__3_/bottom_grid_pin_7_ cbx_2__3_/bottom_grid_pin_8_ cbx_2__3_/bottom_grid_pin_9_
+ sb_2__3_/ccff_tail sb_1__3_/ccff_head cbx_2__3_/chanx_left_in[0] cbx_2__3_/chanx_left_in[10]
+ cbx_2__3_/chanx_left_in[11] cbx_2__3_/chanx_left_in[12] cbx_2__3_/chanx_left_in[13]
+ cbx_2__3_/chanx_left_in[14] cbx_2__3_/chanx_left_in[15] cbx_2__3_/chanx_left_in[16]
+ cbx_2__3_/chanx_left_in[17] cbx_2__3_/chanx_left_in[18] cbx_2__3_/chanx_left_in[19]
+ cbx_2__3_/chanx_left_in[1] cbx_2__3_/chanx_left_in[2] cbx_2__3_/chanx_left_in[3]
+ cbx_2__3_/chanx_left_in[4] cbx_2__3_/chanx_left_in[5] cbx_2__3_/chanx_left_in[6]
+ cbx_2__3_/chanx_left_in[7] cbx_2__3_/chanx_left_in[8] cbx_2__3_/chanx_left_in[9]
+ sb_1__3_/chanx_right_in[0] sb_1__3_/chanx_right_in[10] sb_1__3_/chanx_right_in[11]
+ sb_1__3_/chanx_right_in[12] sb_1__3_/chanx_right_in[13] sb_1__3_/chanx_right_in[14]
+ sb_1__3_/chanx_right_in[15] sb_1__3_/chanx_right_in[16] sb_1__3_/chanx_right_in[17]
+ sb_1__3_/chanx_right_in[18] sb_1__3_/chanx_right_in[19] sb_1__3_/chanx_right_in[1]
+ sb_1__3_/chanx_right_in[2] sb_1__3_/chanx_right_in[3] sb_1__3_/chanx_right_in[4]
+ sb_1__3_/chanx_right_in[5] sb_1__3_/chanx_right_in[6] sb_1__3_/chanx_right_in[7]
+ sb_1__3_/chanx_right_in[8] sb_1__3_/chanx_right_in[9] sb_2__3_/chanx_left_out[0]
+ sb_2__3_/chanx_left_out[10] sb_2__3_/chanx_left_out[11] sb_2__3_/chanx_left_out[12]
+ sb_2__3_/chanx_left_out[13] sb_2__3_/chanx_left_out[14] sb_2__3_/chanx_left_out[15]
+ sb_2__3_/chanx_left_out[16] sb_2__3_/chanx_left_out[17] sb_2__3_/chanx_left_out[18]
+ sb_2__3_/chanx_left_out[19] sb_2__3_/chanx_left_out[1] sb_2__3_/chanx_left_out[2]
+ sb_2__3_/chanx_left_out[3] sb_2__3_/chanx_left_out[4] sb_2__3_/chanx_left_out[5]
+ sb_2__3_/chanx_left_out[6] sb_2__3_/chanx_left_out[7] sb_2__3_/chanx_left_out[8]
+ sb_2__3_/chanx_left_out[9] sb_2__3_/chanx_left_in[0] sb_2__3_/chanx_left_in[10]
+ sb_2__3_/chanx_left_in[11] sb_2__3_/chanx_left_in[12] sb_2__3_/chanx_left_in[13]
+ sb_2__3_/chanx_left_in[14] sb_2__3_/chanx_left_in[15] sb_2__3_/chanx_left_in[16]
+ sb_2__3_/chanx_left_in[17] sb_2__3_/chanx_left_in[18] sb_2__3_/chanx_left_in[19]
+ sb_2__3_/chanx_left_in[1] sb_2__3_/chanx_left_in[2] sb_2__3_/chanx_left_in[3] sb_2__3_/chanx_left_in[4]
+ sb_2__3_/chanx_left_in[5] sb_2__3_/chanx_left_in[6] sb_2__3_/chanx_left_in[7] sb_2__3_/chanx_left_in[8]
+ sb_2__3_/chanx_left_in[9] cbx_2__3_/clk_1_N_out cbx_2__3_/clk_1_S_out sb_1__3_/clk_1_E_out
+ cbx_2__3_/clk_2_E_out cbx_2__3_/clk_2_W_in cbx_2__3_/clk_2_W_out cbx_2__3_/clk_3_E_out
+ cbx_2__3_/clk_3_W_in cbx_2__3_/clk_3_W_out cbx_2__3_/prog_clk_0_N_in cbx_2__3_/prog_clk_0_W_out
+ cbx_2__3_/prog_clk_1_N_out cbx_2__3_/prog_clk_1_S_out sb_1__3_/prog_clk_1_E_out
+ cbx_2__3_/prog_clk_2_E_out cbx_2__3_/prog_clk_2_W_in cbx_2__3_/prog_clk_2_W_out
+ cbx_2__3_/prog_clk_3_E_out cbx_2__3_/prog_clk_3_W_in cbx_2__3_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_6__0_ sb_6__0_/SC_IN_TOP sb_6__0_/SC_OUT_TOP sb_6__0_/Test_en_N_out sb_6__0_/Test_en_S_in
+ VGND VPWR sb_6__0_/ccff_head sb_6__0_/ccff_tail sb_6__0_/chanx_left_in[0] sb_6__0_/chanx_left_in[10]
+ sb_6__0_/chanx_left_in[11] sb_6__0_/chanx_left_in[12] sb_6__0_/chanx_left_in[13]
+ sb_6__0_/chanx_left_in[14] sb_6__0_/chanx_left_in[15] sb_6__0_/chanx_left_in[16]
+ sb_6__0_/chanx_left_in[17] sb_6__0_/chanx_left_in[18] sb_6__0_/chanx_left_in[19]
+ sb_6__0_/chanx_left_in[1] sb_6__0_/chanx_left_in[2] sb_6__0_/chanx_left_in[3] sb_6__0_/chanx_left_in[4]
+ sb_6__0_/chanx_left_in[5] sb_6__0_/chanx_left_in[6] sb_6__0_/chanx_left_in[7] sb_6__0_/chanx_left_in[8]
+ sb_6__0_/chanx_left_in[9] sb_6__0_/chanx_left_out[0] sb_6__0_/chanx_left_out[10]
+ sb_6__0_/chanx_left_out[11] sb_6__0_/chanx_left_out[12] sb_6__0_/chanx_left_out[13]
+ sb_6__0_/chanx_left_out[14] sb_6__0_/chanx_left_out[15] sb_6__0_/chanx_left_out[16]
+ sb_6__0_/chanx_left_out[17] sb_6__0_/chanx_left_out[18] sb_6__0_/chanx_left_out[19]
+ sb_6__0_/chanx_left_out[1] sb_6__0_/chanx_left_out[2] sb_6__0_/chanx_left_out[3]
+ sb_6__0_/chanx_left_out[4] sb_6__0_/chanx_left_out[5] sb_6__0_/chanx_left_out[6]
+ sb_6__0_/chanx_left_out[7] sb_6__0_/chanx_left_out[8] sb_6__0_/chanx_left_out[9]
+ sb_6__0_/chanx_right_in[0] sb_6__0_/chanx_right_in[10] sb_6__0_/chanx_right_in[11]
+ sb_6__0_/chanx_right_in[12] sb_6__0_/chanx_right_in[13] sb_6__0_/chanx_right_in[14]
+ sb_6__0_/chanx_right_in[15] sb_6__0_/chanx_right_in[16] sb_6__0_/chanx_right_in[17]
+ sb_6__0_/chanx_right_in[18] sb_6__0_/chanx_right_in[19] sb_6__0_/chanx_right_in[1]
+ sb_6__0_/chanx_right_in[2] sb_6__0_/chanx_right_in[3] sb_6__0_/chanx_right_in[4]
+ sb_6__0_/chanx_right_in[5] sb_6__0_/chanx_right_in[6] sb_6__0_/chanx_right_in[7]
+ sb_6__0_/chanx_right_in[8] sb_6__0_/chanx_right_in[9] cbx_7__0_/chanx_left_in[0]
+ cbx_7__0_/chanx_left_in[10] cbx_7__0_/chanx_left_in[11] cbx_7__0_/chanx_left_in[12]
+ cbx_7__0_/chanx_left_in[13] cbx_7__0_/chanx_left_in[14] cbx_7__0_/chanx_left_in[15]
+ cbx_7__0_/chanx_left_in[16] cbx_7__0_/chanx_left_in[17] cbx_7__0_/chanx_left_in[18]
+ cbx_7__0_/chanx_left_in[19] cbx_7__0_/chanx_left_in[1] cbx_7__0_/chanx_left_in[2]
+ cbx_7__0_/chanx_left_in[3] cbx_7__0_/chanx_left_in[4] cbx_7__0_/chanx_left_in[5]
+ cbx_7__0_/chanx_left_in[6] cbx_7__0_/chanx_left_in[7] cbx_7__0_/chanx_left_in[8]
+ cbx_7__0_/chanx_left_in[9] sb_6__0_/chany_top_in[0] sb_6__0_/chany_top_in[10] sb_6__0_/chany_top_in[11]
+ sb_6__0_/chany_top_in[12] sb_6__0_/chany_top_in[13] sb_6__0_/chany_top_in[14] sb_6__0_/chany_top_in[15]
+ sb_6__0_/chany_top_in[16] sb_6__0_/chany_top_in[17] sb_6__0_/chany_top_in[18] sb_6__0_/chany_top_in[19]
+ sb_6__0_/chany_top_in[1] sb_6__0_/chany_top_in[2] sb_6__0_/chany_top_in[3] sb_6__0_/chany_top_in[4]
+ sb_6__0_/chany_top_in[5] sb_6__0_/chany_top_in[6] sb_6__0_/chany_top_in[7] sb_6__0_/chany_top_in[8]
+ sb_6__0_/chany_top_in[9] sb_6__0_/chany_top_out[0] sb_6__0_/chany_top_out[10] sb_6__0_/chany_top_out[11]
+ sb_6__0_/chany_top_out[12] sb_6__0_/chany_top_out[13] sb_6__0_/chany_top_out[14]
+ sb_6__0_/chany_top_out[15] sb_6__0_/chany_top_out[16] sb_6__0_/chany_top_out[17]
+ sb_6__0_/chany_top_out[18] sb_6__0_/chany_top_out[19] sb_6__0_/chany_top_out[1]
+ sb_6__0_/chany_top_out[2] sb_6__0_/chany_top_out[3] sb_6__0_/chany_top_out[4] sb_6__0_/chany_top_out[5]
+ sb_6__0_/chany_top_out[6] sb_6__0_/chany_top_out[7] sb_6__0_/chany_top_out[8] sb_6__0_/chany_top_out[9]
+ sb_6__0_/clk_3_N_out sb_6__0_/clk_3_S_in sb_6__0_/left_bottom_grid_pin_11_ sb_6__0_/left_bottom_grid_pin_13_
+ sb_6__0_/left_bottom_grid_pin_15_ sb_6__0_/left_bottom_grid_pin_17_ sb_6__0_/left_bottom_grid_pin_1_
+ sb_6__0_/left_bottom_grid_pin_3_ sb_6__0_/left_bottom_grid_pin_5_ sb_6__0_/left_bottom_grid_pin_7_
+ sb_6__0_/left_bottom_grid_pin_9_ sb_6__0_/prog_clk_0_N_in sb_6__0_/prog_clk_3_N_out
+ sb_6__0_/prog_clk_3_S_in sb_6__0_/right_bottom_grid_pin_11_ sb_6__0_/right_bottom_grid_pin_13_
+ sb_6__0_/right_bottom_grid_pin_15_ sb_6__0_/right_bottom_grid_pin_17_ sb_6__0_/right_bottom_grid_pin_1_
+ sb_6__0_/right_bottom_grid_pin_3_ sb_6__0_/right_bottom_grid_pin_5_ sb_6__0_/right_bottom_grid_pin_7_
+ sb_6__0_/right_bottom_grid_pin_9_ sb_6__0_/top_left_grid_pin_42_ sb_6__0_/top_left_grid_pin_43_
+ sb_6__0_/top_left_grid_pin_44_ sb_6__0_/top_left_grid_pin_45_ sb_6__0_/top_left_grid_pin_46_
+ sb_6__0_/top_left_grid_pin_47_ sb_6__0_/top_left_grid_pin_48_ sb_6__0_/top_left_grid_pin_49_
+ sb_1__0_
Xgrid_clb_1__3_ cbx_1__3_/SC_OUT_BOT cbx_1__2_/SC_IN_TOP grid_clb_1__3_/SC_OUT_TOP
+ cby_1__3_/Test_en_W_out grid_clb_1__3_/Test_en_E_out cby_1__3_/Test_en_W_out grid_clb_1__3_/Test_en_W_out
+ VGND VPWR cbx_1__2_/REGIN_FEEDTHROUGH grid_clb_1__3_/bottom_width_0_height_0__pin_51_
+ cby_0__3_/ccff_tail cby_1__3_/ccff_head cbx_1__3_/clk_1_S_out cbx_1__3_/clk_1_S_out
+ cby_1__3_/prog_clk_0_W_in cbx_1__3_/prog_clk_1_S_out grid_clb_1__3_/prog_clk_0_N_out
+ cbx_1__3_/prog_clk_1_S_out cbx_1__2_/prog_clk_0_N_in cby_0__3_/prog_clk_0_E_in cby_1__3_/left_grid_pin_16_
+ cby_1__3_/left_grid_pin_17_ cby_1__3_/left_grid_pin_18_ cby_1__3_/left_grid_pin_19_
+ cby_1__3_/left_grid_pin_20_ cby_1__3_/left_grid_pin_21_ cby_1__3_/left_grid_pin_22_
+ cby_1__3_/left_grid_pin_23_ cby_1__3_/left_grid_pin_24_ cby_1__3_/left_grid_pin_25_
+ cby_1__3_/left_grid_pin_26_ cby_1__3_/left_grid_pin_27_ cby_1__3_/left_grid_pin_28_
+ cby_1__3_/left_grid_pin_29_ cby_1__3_/left_grid_pin_30_ cby_1__3_/left_grid_pin_31_
+ sb_1__2_/top_left_grid_pin_42_ sb_1__3_/bottom_left_grid_pin_42_ sb_1__2_/top_left_grid_pin_43_
+ sb_1__3_/bottom_left_grid_pin_43_ sb_1__2_/top_left_grid_pin_44_ sb_1__3_/bottom_left_grid_pin_44_
+ sb_1__2_/top_left_grid_pin_45_ sb_1__3_/bottom_left_grid_pin_45_ sb_1__2_/top_left_grid_pin_46_
+ sb_1__3_/bottom_left_grid_pin_46_ sb_1__2_/top_left_grid_pin_47_ sb_1__3_/bottom_left_grid_pin_47_
+ sb_1__2_/top_left_grid_pin_48_ sb_1__3_/bottom_left_grid_pin_48_ sb_1__2_/top_left_grid_pin_49_
+ sb_1__3_/bottom_left_grid_pin_49_ cbx_1__3_/bottom_grid_pin_0_ cbx_1__3_/bottom_grid_pin_10_
+ cbx_1__3_/bottom_grid_pin_11_ cbx_1__3_/bottom_grid_pin_12_ cbx_1__3_/bottom_grid_pin_13_
+ cbx_1__3_/bottom_grid_pin_14_ cbx_1__3_/bottom_grid_pin_15_ cbx_1__3_/bottom_grid_pin_1_
+ cbx_1__3_/bottom_grid_pin_2_ cbx_1__3_/REGOUT_FEEDTHROUGH grid_clb_1__3_/top_width_0_height_0__pin_33_
+ sb_1__3_/left_bottom_grid_pin_34_ sb_0__3_/right_bottom_grid_pin_34_ sb_1__3_/left_bottom_grid_pin_35_
+ sb_0__3_/right_bottom_grid_pin_35_ sb_1__3_/left_bottom_grid_pin_36_ sb_0__3_/right_bottom_grid_pin_36_
+ sb_1__3_/left_bottom_grid_pin_37_ sb_0__3_/right_bottom_grid_pin_37_ sb_1__3_/left_bottom_grid_pin_38_
+ sb_0__3_/right_bottom_grid_pin_38_ sb_1__3_/left_bottom_grid_pin_39_ sb_0__3_/right_bottom_grid_pin_39_
+ cbx_1__3_/bottom_grid_pin_3_ sb_1__3_/left_bottom_grid_pin_40_ sb_0__3_/right_bottom_grid_pin_40_
+ sb_1__3_/left_bottom_grid_pin_41_ sb_0__3_/right_bottom_grid_pin_41_ cbx_1__3_/bottom_grid_pin_4_
+ cbx_1__3_/bottom_grid_pin_5_ cbx_1__3_/bottom_grid_pin_6_ cbx_1__3_/bottom_grid_pin_7_
+ cbx_1__3_/bottom_grid_pin_8_ cbx_1__3_/bottom_grid_pin_9_ grid_clb
Xcby_8__7_ IO_ISOL_N VGND VPWR cby_8__7_/ccff_head sb_8__6_/ccff_head sb_8__6_/chany_top_out[0]
+ sb_8__6_/chany_top_out[10] sb_8__6_/chany_top_out[11] sb_8__6_/chany_top_out[12]
+ sb_8__6_/chany_top_out[13] sb_8__6_/chany_top_out[14] sb_8__6_/chany_top_out[15]
+ sb_8__6_/chany_top_out[16] sb_8__6_/chany_top_out[17] sb_8__6_/chany_top_out[18]
+ sb_8__6_/chany_top_out[19] sb_8__6_/chany_top_out[1] sb_8__6_/chany_top_out[2] sb_8__6_/chany_top_out[3]
+ sb_8__6_/chany_top_out[4] sb_8__6_/chany_top_out[5] sb_8__6_/chany_top_out[6] sb_8__6_/chany_top_out[7]
+ sb_8__6_/chany_top_out[8] sb_8__6_/chany_top_out[9] sb_8__6_/chany_top_in[0] sb_8__6_/chany_top_in[10]
+ sb_8__6_/chany_top_in[11] sb_8__6_/chany_top_in[12] sb_8__6_/chany_top_in[13] sb_8__6_/chany_top_in[14]
+ sb_8__6_/chany_top_in[15] sb_8__6_/chany_top_in[16] sb_8__6_/chany_top_in[17] sb_8__6_/chany_top_in[18]
+ sb_8__6_/chany_top_in[19] sb_8__6_/chany_top_in[1] sb_8__6_/chany_top_in[2] sb_8__6_/chany_top_in[3]
+ sb_8__6_/chany_top_in[4] sb_8__6_/chany_top_in[5] sb_8__6_/chany_top_in[6] sb_8__6_/chany_top_in[7]
+ sb_8__6_/chany_top_in[8] sb_8__6_/chany_top_in[9] cby_8__7_/chany_top_in[0] cby_8__7_/chany_top_in[10]
+ cby_8__7_/chany_top_in[11] cby_8__7_/chany_top_in[12] cby_8__7_/chany_top_in[13]
+ cby_8__7_/chany_top_in[14] cby_8__7_/chany_top_in[15] cby_8__7_/chany_top_in[16]
+ cby_8__7_/chany_top_in[17] cby_8__7_/chany_top_in[18] cby_8__7_/chany_top_in[19]
+ cby_8__7_/chany_top_in[1] cby_8__7_/chany_top_in[2] cby_8__7_/chany_top_in[3] cby_8__7_/chany_top_in[4]
+ cby_8__7_/chany_top_in[5] cby_8__7_/chany_top_in[6] cby_8__7_/chany_top_in[7] cby_8__7_/chany_top_in[8]
+ cby_8__7_/chany_top_in[9] cby_8__7_/chany_top_out[0] cby_8__7_/chany_top_out[10]
+ cby_8__7_/chany_top_out[11] cby_8__7_/chany_top_out[12] cby_8__7_/chany_top_out[13]
+ cby_8__7_/chany_top_out[14] cby_8__7_/chany_top_out[15] cby_8__7_/chany_top_out[16]
+ cby_8__7_/chany_top_out[17] cby_8__7_/chany_top_out[18] cby_8__7_/chany_top_out[19]
+ cby_8__7_/chany_top_out[1] cby_8__7_/chany_top_out[2] cby_8__7_/chany_top_out[3]
+ cby_8__7_/chany_top_out[4] cby_8__7_/chany_top_out[5] cby_8__7_/chany_top_out[6]
+ cby_8__7_/chany_top_out[7] cby_8__7_/chany_top_out[8] cby_8__7_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
+ cby_8__7_/left_grid_pin_16_ cby_8__7_/left_grid_pin_17_ cby_8__7_/left_grid_pin_18_
+ cby_8__7_/left_grid_pin_19_ cby_8__7_/left_grid_pin_20_ cby_8__7_/left_grid_pin_21_
+ cby_8__7_/left_grid_pin_22_ cby_8__7_/left_grid_pin_23_ cby_8__7_/left_grid_pin_24_
+ cby_8__7_/left_grid_pin_25_ cby_8__7_/left_grid_pin_26_ cby_8__7_/left_grid_pin_27_
+ cby_8__7_/left_grid_pin_28_ cby_8__7_/left_grid_pin_29_ cby_8__7_/left_grid_pin_30_
+ cby_8__7_/left_grid_pin_31_ cby_8__7_/right_grid_pin_0_ sb_8__6_/top_right_grid_pin_1_
+ sb_8__7_/bottom_right_grid_pin_1_ cby_8__7_/prog_clk_0_N_out sb_8__6_/prog_clk_0_N_in
+ cby_8__7_/prog_clk_0_W_in cby_8__7_/right_grid_pin_0_ cby_2__1_
Xcbx_8__8_ IO_ISOL_N cbx_8__8_/SC_IN_BOT cbx_8__8_/SC_IN_TOP cbx_8__8_/SC_OUT_BOT
+ sb_8__8_/SC_IN_BOT VGND VPWR cbx_8__8_/bottom_grid_pin_0_ cbx_8__8_/bottom_grid_pin_10_
+ cbx_8__8_/bottom_grid_pin_11_ cbx_8__8_/bottom_grid_pin_12_ cbx_8__8_/bottom_grid_pin_13_
+ cbx_8__8_/bottom_grid_pin_14_ cbx_8__8_/bottom_grid_pin_15_ cbx_8__8_/bottom_grid_pin_1_
+ cbx_8__8_/bottom_grid_pin_2_ cbx_8__8_/bottom_grid_pin_3_ cbx_8__8_/bottom_grid_pin_4_
+ cbx_8__8_/bottom_grid_pin_5_ cbx_8__8_/bottom_grid_pin_6_ cbx_8__8_/bottom_grid_pin_7_
+ cbx_8__8_/bottom_grid_pin_8_ cbx_8__8_/bottom_grid_pin_9_ cbx_8__8_/top_grid_pin_0_
+ sb_8__8_/left_top_grid_pin_1_ sb_7__8_/right_top_grid_pin_1_ sb_8__8_/ccff_tail
+ sb_7__8_/ccff_head cbx_8__8_/chanx_left_in[0] cbx_8__8_/chanx_left_in[10] cbx_8__8_/chanx_left_in[11]
+ cbx_8__8_/chanx_left_in[12] cbx_8__8_/chanx_left_in[13] cbx_8__8_/chanx_left_in[14]
+ cbx_8__8_/chanx_left_in[15] cbx_8__8_/chanx_left_in[16] cbx_8__8_/chanx_left_in[17]
+ cbx_8__8_/chanx_left_in[18] cbx_8__8_/chanx_left_in[19] cbx_8__8_/chanx_left_in[1]
+ cbx_8__8_/chanx_left_in[2] cbx_8__8_/chanx_left_in[3] cbx_8__8_/chanx_left_in[4]
+ cbx_8__8_/chanx_left_in[5] cbx_8__8_/chanx_left_in[6] cbx_8__8_/chanx_left_in[7]
+ cbx_8__8_/chanx_left_in[8] cbx_8__8_/chanx_left_in[9] sb_7__8_/chanx_right_in[0]
+ sb_7__8_/chanx_right_in[10] sb_7__8_/chanx_right_in[11] sb_7__8_/chanx_right_in[12]
+ sb_7__8_/chanx_right_in[13] sb_7__8_/chanx_right_in[14] sb_7__8_/chanx_right_in[15]
+ sb_7__8_/chanx_right_in[16] sb_7__8_/chanx_right_in[17] sb_7__8_/chanx_right_in[18]
+ sb_7__8_/chanx_right_in[19] sb_7__8_/chanx_right_in[1] sb_7__8_/chanx_right_in[2]
+ sb_7__8_/chanx_right_in[3] sb_7__8_/chanx_right_in[4] sb_7__8_/chanx_right_in[5]
+ sb_7__8_/chanx_right_in[6] sb_7__8_/chanx_right_in[7] sb_7__8_/chanx_right_in[8]
+ sb_7__8_/chanx_right_in[9] sb_8__8_/chanx_left_out[0] sb_8__8_/chanx_left_out[10]
+ sb_8__8_/chanx_left_out[11] sb_8__8_/chanx_left_out[12] sb_8__8_/chanx_left_out[13]
+ sb_8__8_/chanx_left_out[14] sb_8__8_/chanx_left_out[15] sb_8__8_/chanx_left_out[16]
+ sb_8__8_/chanx_left_out[17] sb_8__8_/chanx_left_out[18] sb_8__8_/chanx_left_out[19]
+ sb_8__8_/chanx_left_out[1] sb_8__8_/chanx_left_out[2] sb_8__8_/chanx_left_out[3]
+ sb_8__8_/chanx_left_out[4] sb_8__8_/chanx_left_out[5] sb_8__8_/chanx_left_out[6]
+ sb_8__8_/chanx_left_out[7] sb_8__8_/chanx_left_out[8] sb_8__8_/chanx_left_out[9]
+ sb_8__8_/chanx_left_in[0] sb_8__8_/chanx_left_in[10] sb_8__8_/chanx_left_in[11]
+ sb_8__8_/chanx_left_in[12] sb_8__8_/chanx_left_in[13] sb_8__8_/chanx_left_in[14]
+ sb_8__8_/chanx_left_in[15] sb_8__8_/chanx_left_in[16] sb_8__8_/chanx_left_in[17]
+ sb_8__8_/chanx_left_in[18] sb_8__8_/chanx_left_in[19] sb_8__8_/chanx_left_in[1]
+ sb_8__8_/chanx_left_in[2] sb_8__8_/chanx_left_in[3] sb_8__8_/chanx_left_in[4] sb_8__8_/chanx_left_in[5]
+ sb_8__8_/chanx_left_in[6] sb_8__8_/chanx_left_in[7] sb_8__8_/chanx_left_in[8] sb_8__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
+ cbx_8__8_/prog_clk_0_S_in cbx_8__8_/prog_clk_0_W_out cbx_8__8_/top_grid_pin_0_ cbx_1__2_
Xcby_5__4_ cby_5__4_/Test_en_W_in cby_5__4_/Test_en_E_out cby_5__4_/Test_en_N_out
+ cby_5__4_/Test_en_W_in cby_5__4_/Test_en_W_in cby_5__4_/Test_en_W_out VGND VPWR
+ cby_5__4_/ccff_head cby_5__4_/ccff_tail sb_5__3_/chany_top_out[0] sb_5__3_/chany_top_out[10]
+ sb_5__3_/chany_top_out[11] sb_5__3_/chany_top_out[12] sb_5__3_/chany_top_out[13]
+ sb_5__3_/chany_top_out[14] sb_5__3_/chany_top_out[15] sb_5__3_/chany_top_out[16]
+ sb_5__3_/chany_top_out[17] sb_5__3_/chany_top_out[18] sb_5__3_/chany_top_out[19]
+ sb_5__3_/chany_top_out[1] sb_5__3_/chany_top_out[2] sb_5__3_/chany_top_out[3] sb_5__3_/chany_top_out[4]
+ sb_5__3_/chany_top_out[5] sb_5__3_/chany_top_out[6] sb_5__3_/chany_top_out[7] sb_5__3_/chany_top_out[8]
+ sb_5__3_/chany_top_out[9] sb_5__3_/chany_top_in[0] sb_5__3_/chany_top_in[10] sb_5__3_/chany_top_in[11]
+ sb_5__3_/chany_top_in[12] sb_5__3_/chany_top_in[13] sb_5__3_/chany_top_in[14] sb_5__3_/chany_top_in[15]
+ sb_5__3_/chany_top_in[16] sb_5__3_/chany_top_in[17] sb_5__3_/chany_top_in[18] sb_5__3_/chany_top_in[19]
+ sb_5__3_/chany_top_in[1] sb_5__3_/chany_top_in[2] sb_5__3_/chany_top_in[3] sb_5__3_/chany_top_in[4]
+ sb_5__3_/chany_top_in[5] sb_5__3_/chany_top_in[6] sb_5__3_/chany_top_in[7] sb_5__3_/chany_top_in[8]
+ sb_5__3_/chany_top_in[9] cby_5__4_/chany_top_in[0] cby_5__4_/chany_top_in[10] cby_5__4_/chany_top_in[11]
+ cby_5__4_/chany_top_in[12] cby_5__4_/chany_top_in[13] cby_5__4_/chany_top_in[14]
+ cby_5__4_/chany_top_in[15] cby_5__4_/chany_top_in[16] cby_5__4_/chany_top_in[17]
+ cby_5__4_/chany_top_in[18] cby_5__4_/chany_top_in[19] cby_5__4_/chany_top_in[1]
+ cby_5__4_/chany_top_in[2] cby_5__4_/chany_top_in[3] cby_5__4_/chany_top_in[4] cby_5__4_/chany_top_in[5]
+ cby_5__4_/chany_top_in[6] cby_5__4_/chany_top_in[7] cby_5__4_/chany_top_in[8] cby_5__4_/chany_top_in[9]
+ cby_5__4_/chany_top_out[0] cby_5__4_/chany_top_out[10] cby_5__4_/chany_top_out[11]
+ cby_5__4_/chany_top_out[12] cby_5__4_/chany_top_out[13] cby_5__4_/chany_top_out[14]
+ cby_5__4_/chany_top_out[15] cby_5__4_/chany_top_out[16] cby_5__4_/chany_top_out[17]
+ cby_5__4_/chany_top_out[18] cby_5__4_/chany_top_out[19] cby_5__4_/chany_top_out[1]
+ cby_5__4_/chany_top_out[2] cby_5__4_/chany_top_out[3] cby_5__4_/chany_top_out[4]
+ cby_5__4_/chany_top_out[5] cby_5__4_/chany_top_out[6] cby_5__4_/chany_top_out[7]
+ cby_5__4_/chany_top_out[8] cby_5__4_/chany_top_out[9] cby_5__4_/clk_2_N_out cby_5__4_/clk_2_S_in
+ cby_5__4_/clk_2_S_out cby_5__4_/clk_3_N_out cby_5__4_/clk_3_S_in cby_5__4_/clk_3_S_out
+ cby_5__4_/left_grid_pin_16_ cby_5__4_/left_grid_pin_17_ cby_5__4_/left_grid_pin_18_
+ cby_5__4_/left_grid_pin_19_ cby_5__4_/left_grid_pin_20_ cby_5__4_/left_grid_pin_21_
+ cby_5__4_/left_grid_pin_22_ cby_5__4_/left_grid_pin_23_ cby_5__4_/left_grid_pin_24_
+ cby_5__4_/left_grid_pin_25_ cby_5__4_/left_grid_pin_26_ cby_5__4_/left_grid_pin_27_
+ cby_5__4_/left_grid_pin_28_ cby_5__4_/left_grid_pin_29_ cby_5__4_/left_grid_pin_30_
+ cby_5__4_/left_grid_pin_31_ cby_5__4_/prog_clk_0_N_out sb_5__3_/prog_clk_0_N_in
+ cby_5__4_/prog_clk_0_W_in cby_5__4_/prog_clk_2_N_out cby_5__4_/prog_clk_2_S_in cby_5__4_/prog_clk_2_S_out
+ cby_5__4_/prog_clk_3_N_out cby_5__4_/prog_clk_3_S_in cby_5__4_/prog_clk_3_S_out
+ cby_1__1_
Xcby_2__1_ cby_2__1_/Test_en_W_in cby_2__1_/Test_en_E_out cby_2__1_/Test_en_N_out
+ cby_2__1_/Test_en_W_in cby_2__1_/Test_en_W_in cby_2__1_/Test_en_W_out VGND VPWR
+ cby_2__1_/ccff_head cby_2__1_/ccff_tail sb_2__0_/chany_top_out[0] sb_2__0_/chany_top_out[10]
+ sb_2__0_/chany_top_out[11] sb_2__0_/chany_top_out[12] sb_2__0_/chany_top_out[13]
+ sb_2__0_/chany_top_out[14] sb_2__0_/chany_top_out[15] sb_2__0_/chany_top_out[16]
+ sb_2__0_/chany_top_out[17] sb_2__0_/chany_top_out[18] sb_2__0_/chany_top_out[19]
+ sb_2__0_/chany_top_out[1] sb_2__0_/chany_top_out[2] sb_2__0_/chany_top_out[3] sb_2__0_/chany_top_out[4]
+ sb_2__0_/chany_top_out[5] sb_2__0_/chany_top_out[6] sb_2__0_/chany_top_out[7] sb_2__0_/chany_top_out[8]
+ sb_2__0_/chany_top_out[9] sb_2__0_/chany_top_in[0] sb_2__0_/chany_top_in[10] sb_2__0_/chany_top_in[11]
+ sb_2__0_/chany_top_in[12] sb_2__0_/chany_top_in[13] sb_2__0_/chany_top_in[14] sb_2__0_/chany_top_in[15]
+ sb_2__0_/chany_top_in[16] sb_2__0_/chany_top_in[17] sb_2__0_/chany_top_in[18] sb_2__0_/chany_top_in[19]
+ sb_2__0_/chany_top_in[1] sb_2__0_/chany_top_in[2] sb_2__0_/chany_top_in[3] sb_2__0_/chany_top_in[4]
+ sb_2__0_/chany_top_in[5] sb_2__0_/chany_top_in[6] sb_2__0_/chany_top_in[7] sb_2__0_/chany_top_in[8]
+ sb_2__0_/chany_top_in[9] cby_2__1_/chany_top_in[0] cby_2__1_/chany_top_in[10] cby_2__1_/chany_top_in[11]
+ cby_2__1_/chany_top_in[12] cby_2__1_/chany_top_in[13] cby_2__1_/chany_top_in[14]
+ cby_2__1_/chany_top_in[15] cby_2__1_/chany_top_in[16] cby_2__1_/chany_top_in[17]
+ cby_2__1_/chany_top_in[18] cby_2__1_/chany_top_in[19] cby_2__1_/chany_top_in[1]
+ cby_2__1_/chany_top_in[2] cby_2__1_/chany_top_in[3] cby_2__1_/chany_top_in[4] cby_2__1_/chany_top_in[5]
+ cby_2__1_/chany_top_in[6] cby_2__1_/chany_top_in[7] cby_2__1_/chany_top_in[8] cby_2__1_/chany_top_in[9]
+ cby_2__1_/chany_top_out[0] cby_2__1_/chany_top_out[10] cby_2__1_/chany_top_out[11]
+ cby_2__1_/chany_top_out[12] cby_2__1_/chany_top_out[13] cby_2__1_/chany_top_out[14]
+ cby_2__1_/chany_top_out[15] cby_2__1_/chany_top_out[16] cby_2__1_/chany_top_out[17]
+ cby_2__1_/chany_top_out[18] cby_2__1_/chany_top_out[19] cby_2__1_/chany_top_out[1]
+ cby_2__1_/chany_top_out[2] cby_2__1_/chany_top_out[3] cby_2__1_/chany_top_out[4]
+ cby_2__1_/chany_top_out[5] cby_2__1_/chany_top_out[6] cby_2__1_/chany_top_out[7]
+ cby_2__1_/chany_top_out[8] cby_2__1_/chany_top_out[9] cby_2__1_/clk_2_N_out cby_2__1_/clk_2_S_in
+ cby_2__1_/clk_2_S_out cby_2__1_/clk_3_N_out cby_2__1_/clk_3_S_in cby_2__1_/clk_3_S_out
+ cby_2__1_/left_grid_pin_16_ cby_2__1_/left_grid_pin_17_ cby_2__1_/left_grid_pin_18_
+ cby_2__1_/left_grid_pin_19_ cby_2__1_/left_grid_pin_20_ cby_2__1_/left_grid_pin_21_
+ cby_2__1_/left_grid_pin_22_ cby_2__1_/left_grid_pin_23_ cby_2__1_/left_grid_pin_24_
+ cby_2__1_/left_grid_pin_25_ cby_2__1_/left_grid_pin_26_ cby_2__1_/left_grid_pin_27_
+ cby_2__1_/left_grid_pin_28_ cby_2__1_/left_grid_pin_29_ cby_2__1_/left_grid_pin_30_
+ cby_2__1_/left_grid_pin_31_ cby_2__1_/prog_clk_0_N_out sb_2__0_/prog_clk_0_N_in
+ cby_2__1_/prog_clk_0_W_in cby_2__1_/prog_clk_2_N_out cby_2__1_/prog_clk_2_S_in cby_2__1_/prog_clk_2_S_out
+ cby_2__1_/prog_clk_3_N_out cby_2__1_/prog_clk_3_S_in cby_2__1_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_7__8_ cbx_7__8_/SC_OUT_BOT cbx_7__7_/SC_IN_TOP grid_clb_7__8_/SC_OUT_TOP
+ cby_6__8_/Test_en_E_out cby_7__8_/Test_en_W_in cby_6__8_/Test_en_E_out grid_clb_7__8_/Test_en_W_out
+ VGND VPWR cbx_7__7_/REGIN_FEEDTHROUGH grid_clb_7__8_/bottom_width_0_height_0__pin_51_
+ cby_6__8_/ccff_tail cby_7__8_/ccff_head cbx_7__7_/clk_1_N_out cbx_7__7_/clk_1_N_out
+ cby_7__8_/prog_clk_0_W_in cbx_7__7_/prog_clk_1_N_out cbx_7__8_/prog_clk_0_S_in cbx_7__7_/prog_clk_1_N_out
+ cbx_7__7_/prog_clk_0_N_in grid_clb_7__8_/prog_clk_0_W_out cby_7__8_/left_grid_pin_16_
+ cby_7__8_/left_grid_pin_17_ cby_7__8_/left_grid_pin_18_ cby_7__8_/left_grid_pin_19_
+ cby_7__8_/left_grid_pin_20_ cby_7__8_/left_grid_pin_21_ cby_7__8_/left_grid_pin_22_
+ cby_7__8_/left_grid_pin_23_ cby_7__8_/left_grid_pin_24_ cby_7__8_/left_grid_pin_25_
+ cby_7__8_/left_grid_pin_26_ cby_7__8_/left_grid_pin_27_ cby_7__8_/left_grid_pin_28_
+ cby_7__8_/left_grid_pin_29_ cby_7__8_/left_grid_pin_30_ cby_7__8_/left_grid_pin_31_
+ sb_7__7_/top_left_grid_pin_42_ sb_7__8_/bottom_left_grid_pin_42_ sb_7__7_/top_left_grid_pin_43_
+ sb_7__8_/bottom_left_grid_pin_43_ sb_7__7_/top_left_grid_pin_44_ sb_7__8_/bottom_left_grid_pin_44_
+ sb_7__7_/top_left_grid_pin_45_ sb_7__8_/bottom_left_grid_pin_45_ sb_7__7_/top_left_grid_pin_46_
+ sb_7__8_/bottom_left_grid_pin_46_ sb_7__7_/top_left_grid_pin_47_ sb_7__8_/bottom_left_grid_pin_47_
+ sb_7__7_/top_left_grid_pin_48_ sb_7__8_/bottom_left_grid_pin_48_ sb_7__7_/top_left_grid_pin_49_
+ sb_7__8_/bottom_left_grid_pin_49_ cbx_7__8_/bottom_grid_pin_0_ cbx_7__8_/bottom_grid_pin_10_
+ cbx_7__8_/bottom_grid_pin_11_ cbx_7__8_/bottom_grid_pin_12_ cbx_7__8_/bottom_grid_pin_13_
+ cbx_7__8_/bottom_grid_pin_14_ cbx_7__8_/bottom_grid_pin_15_ cbx_7__8_/bottom_grid_pin_1_
+ cbx_7__8_/bottom_grid_pin_2_ tie_array/x[6] grid_clb_7__8_/top_width_0_height_0__pin_33_
+ sb_7__8_/left_bottom_grid_pin_34_ sb_6__8_/right_bottom_grid_pin_34_ sb_7__8_/left_bottom_grid_pin_35_
+ sb_6__8_/right_bottom_grid_pin_35_ sb_7__8_/left_bottom_grid_pin_36_ sb_6__8_/right_bottom_grid_pin_36_
+ sb_7__8_/left_bottom_grid_pin_37_ sb_6__8_/right_bottom_grid_pin_37_ sb_7__8_/left_bottom_grid_pin_38_
+ sb_6__8_/right_bottom_grid_pin_38_ sb_7__8_/left_bottom_grid_pin_39_ sb_6__8_/right_bottom_grid_pin_39_
+ cbx_7__8_/bottom_grid_pin_3_ sb_7__8_/left_bottom_grid_pin_40_ sb_6__8_/right_bottom_grid_pin_40_
+ sb_7__8_/left_bottom_grid_pin_41_ sb_6__8_/right_bottom_grid_pin_41_ cbx_7__8_/bottom_grid_pin_4_
+ cbx_7__8_/bottom_grid_pin_5_ cbx_7__8_/bottom_grid_pin_6_ cbx_7__8_/bottom_grid_pin_7_
+ cbx_7__8_/bottom_grid_pin_8_ cbx_7__8_/bottom_grid_pin_9_ grid_clb
Xcbx_5__5_ cbx_5__5_/REGIN_FEEDTHROUGH cbx_5__5_/REGOUT_FEEDTHROUGH cbx_5__5_/SC_IN_BOT
+ cbx_5__5_/SC_IN_TOP cbx_5__5_/SC_OUT_BOT cbx_5__5_/SC_OUT_TOP VGND VPWR cbx_5__5_/bottom_grid_pin_0_
+ cbx_5__5_/bottom_grid_pin_10_ cbx_5__5_/bottom_grid_pin_11_ cbx_5__5_/bottom_grid_pin_12_
+ cbx_5__5_/bottom_grid_pin_13_ cbx_5__5_/bottom_grid_pin_14_ cbx_5__5_/bottom_grid_pin_15_
+ cbx_5__5_/bottom_grid_pin_1_ cbx_5__5_/bottom_grid_pin_2_ cbx_5__5_/bottom_grid_pin_3_
+ cbx_5__5_/bottom_grid_pin_4_ cbx_5__5_/bottom_grid_pin_5_ cbx_5__5_/bottom_grid_pin_6_
+ cbx_5__5_/bottom_grid_pin_7_ cbx_5__5_/bottom_grid_pin_8_ cbx_5__5_/bottom_grid_pin_9_
+ sb_5__5_/ccff_tail sb_4__5_/ccff_head cbx_5__5_/chanx_left_in[0] cbx_5__5_/chanx_left_in[10]
+ cbx_5__5_/chanx_left_in[11] cbx_5__5_/chanx_left_in[12] cbx_5__5_/chanx_left_in[13]
+ cbx_5__5_/chanx_left_in[14] cbx_5__5_/chanx_left_in[15] cbx_5__5_/chanx_left_in[16]
+ cbx_5__5_/chanx_left_in[17] cbx_5__5_/chanx_left_in[18] cbx_5__5_/chanx_left_in[19]
+ cbx_5__5_/chanx_left_in[1] cbx_5__5_/chanx_left_in[2] cbx_5__5_/chanx_left_in[3]
+ cbx_5__5_/chanx_left_in[4] cbx_5__5_/chanx_left_in[5] cbx_5__5_/chanx_left_in[6]
+ cbx_5__5_/chanx_left_in[7] cbx_5__5_/chanx_left_in[8] cbx_5__5_/chanx_left_in[9]
+ sb_4__5_/chanx_right_in[0] sb_4__5_/chanx_right_in[10] sb_4__5_/chanx_right_in[11]
+ sb_4__5_/chanx_right_in[12] sb_4__5_/chanx_right_in[13] sb_4__5_/chanx_right_in[14]
+ sb_4__5_/chanx_right_in[15] sb_4__5_/chanx_right_in[16] sb_4__5_/chanx_right_in[17]
+ sb_4__5_/chanx_right_in[18] sb_4__5_/chanx_right_in[19] sb_4__5_/chanx_right_in[1]
+ sb_4__5_/chanx_right_in[2] sb_4__5_/chanx_right_in[3] sb_4__5_/chanx_right_in[4]
+ sb_4__5_/chanx_right_in[5] sb_4__5_/chanx_right_in[6] sb_4__5_/chanx_right_in[7]
+ sb_4__5_/chanx_right_in[8] sb_4__5_/chanx_right_in[9] sb_5__5_/chanx_left_out[0]
+ sb_5__5_/chanx_left_out[10] sb_5__5_/chanx_left_out[11] sb_5__5_/chanx_left_out[12]
+ sb_5__5_/chanx_left_out[13] sb_5__5_/chanx_left_out[14] sb_5__5_/chanx_left_out[15]
+ sb_5__5_/chanx_left_out[16] sb_5__5_/chanx_left_out[17] sb_5__5_/chanx_left_out[18]
+ sb_5__5_/chanx_left_out[19] sb_5__5_/chanx_left_out[1] sb_5__5_/chanx_left_out[2]
+ sb_5__5_/chanx_left_out[3] sb_5__5_/chanx_left_out[4] sb_5__5_/chanx_left_out[5]
+ sb_5__5_/chanx_left_out[6] sb_5__5_/chanx_left_out[7] sb_5__5_/chanx_left_out[8]
+ sb_5__5_/chanx_left_out[9] sb_5__5_/chanx_left_in[0] sb_5__5_/chanx_left_in[10]
+ sb_5__5_/chanx_left_in[11] sb_5__5_/chanx_left_in[12] sb_5__5_/chanx_left_in[13]
+ sb_5__5_/chanx_left_in[14] sb_5__5_/chanx_left_in[15] sb_5__5_/chanx_left_in[16]
+ sb_5__5_/chanx_left_in[17] sb_5__5_/chanx_left_in[18] sb_5__5_/chanx_left_in[19]
+ sb_5__5_/chanx_left_in[1] sb_5__5_/chanx_left_in[2] sb_5__5_/chanx_left_in[3] sb_5__5_/chanx_left_in[4]
+ sb_5__5_/chanx_left_in[5] sb_5__5_/chanx_left_in[6] sb_5__5_/chanx_left_in[7] sb_5__5_/chanx_left_in[8]
+ sb_5__5_/chanx_left_in[9] cbx_5__5_/clk_1_N_out cbx_5__5_/clk_1_S_out sb_5__5_/clk_1_W_out
+ cbx_5__5_/clk_2_E_out cbx_5__5_/clk_2_W_in cbx_5__5_/clk_2_W_out cbx_5__5_/clk_3_E_out
+ cbx_5__5_/clk_3_W_in cbx_5__5_/clk_3_W_out cbx_5__5_/prog_clk_0_N_in cbx_5__5_/prog_clk_0_W_out
+ cbx_5__5_/prog_clk_1_N_out cbx_5__5_/prog_clk_1_S_out sb_5__5_/prog_clk_1_W_out
+ cbx_5__5_/prog_clk_2_E_out cbx_5__5_/prog_clk_2_W_in cbx_5__5_/prog_clk_2_W_out
+ cbx_5__5_/prog_clk_3_E_out cbx_5__5_/prog_clk_3_W_in cbx_5__5_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_4__5_ cbx_4__4_/SC_OUT_TOP grid_clb_4__5_/SC_OUT_BOT cbx_4__5_/SC_IN_BOT
+ cby_4__5_/Test_en_W_out grid_clb_4__5_/Test_en_E_out cby_4__5_/Test_en_W_out cby_3__5_/Test_en_W_in
+ VGND VPWR cbx_4__4_/REGIN_FEEDTHROUGH grid_clb_4__5_/bottom_width_0_height_0__pin_51_
+ cby_3__5_/ccff_tail cby_4__5_/ccff_head cbx_4__5_/clk_1_S_out cbx_4__5_/clk_1_S_out
+ cby_4__5_/prog_clk_0_W_in cbx_4__5_/prog_clk_1_S_out grid_clb_4__5_/prog_clk_0_N_out
+ cbx_4__5_/prog_clk_1_S_out cbx_4__4_/prog_clk_0_N_in grid_clb_4__5_/prog_clk_0_W_out
+ cby_4__5_/left_grid_pin_16_ cby_4__5_/left_grid_pin_17_ cby_4__5_/left_grid_pin_18_
+ cby_4__5_/left_grid_pin_19_ cby_4__5_/left_grid_pin_20_ cby_4__5_/left_grid_pin_21_
+ cby_4__5_/left_grid_pin_22_ cby_4__5_/left_grid_pin_23_ cby_4__5_/left_grid_pin_24_
+ cby_4__5_/left_grid_pin_25_ cby_4__5_/left_grid_pin_26_ cby_4__5_/left_grid_pin_27_
+ cby_4__5_/left_grid_pin_28_ cby_4__5_/left_grid_pin_29_ cby_4__5_/left_grid_pin_30_
+ cby_4__5_/left_grid_pin_31_ sb_4__4_/top_left_grid_pin_42_ sb_4__5_/bottom_left_grid_pin_42_
+ sb_4__4_/top_left_grid_pin_43_ sb_4__5_/bottom_left_grid_pin_43_ sb_4__4_/top_left_grid_pin_44_
+ sb_4__5_/bottom_left_grid_pin_44_ sb_4__4_/top_left_grid_pin_45_ sb_4__5_/bottom_left_grid_pin_45_
+ sb_4__4_/top_left_grid_pin_46_ sb_4__5_/bottom_left_grid_pin_46_ sb_4__4_/top_left_grid_pin_47_
+ sb_4__5_/bottom_left_grid_pin_47_ sb_4__4_/top_left_grid_pin_48_ sb_4__5_/bottom_left_grid_pin_48_
+ sb_4__4_/top_left_grid_pin_49_ sb_4__5_/bottom_left_grid_pin_49_ cbx_4__5_/bottom_grid_pin_0_
+ cbx_4__5_/bottom_grid_pin_10_ cbx_4__5_/bottom_grid_pin_11_ cbx_4__5_/bottom_grid_pin_12_
+ cbx_4__5_/bottom_grid_pin_13_ cbx_4__5_/bottom_grid_pin_14_ cbx_4__5_/bottom_grid_pin_15_
+ cbx_4__5_/bottom_grid_pin_1_ cbx_4__5_/bottom_grid_pin_2_ cbx_4__5_/REGOUT_FEEDTHROUGH
+ grid_clb_4__5_/top_width_0_height_0__pin_33_ sb_4__5_/left_bottom_grid_pin_34_ sb_3__5_/right_bottom_grid_pin_34_
+ sb_4__5_/left_bottom_grid_pin_35_ sb_3__5_/right_bottom_grid_pin_35_ sb_4__5_/left_bottom_grid_pin_36_
+ sb_3__5_/right_bottom_grid_pin_36_ sb_4__5_/left_bottom_grid_pin_37_ sb_3__5_/right_bottom_grid_pin_37_
+ sb_4__5_/left_bottom_grid_pin_38_ sb_3__5_/right_bottom_grid_pin_38_ sb_4__5_/left_bottom_grid_pin_39_
+ sb_3__5_/right_bottom_grid_pin_39_ cbx_4__5_/bottom_grid_pin_3_ sb_4__5_/left_bottom_grid_pin_40_
+ sb_3__5_/right_bottom_grid_pin_40_ sb_4__5_/left_bottom_grid_pin_41_ sb_3__5_/right_bottom_grid_pin_41_
+ cbx_4__5_/bottom_grid_pin_4_ cbx_4__5_/bottom_grid_pin_5_ cbx_4__5_/bottom_grid_pin_6_
+ cbx_4__5_/bottom_grid_pin_7_ cbx_4__5_/bottom_grid_pin_8_ cbx_4__5_/bottom_grid_pin_9_
+ grid_clb
Xcbx_2__2_ cbx_2__2_/REGIN_FEEDTHROUGH cbx_2__2_/REGOUT_FEEDTHROUGH cbx_2__2_/SC_IN_BOT
+ cbx_2__2_/SC_IN_TOP cbx_2__2_/SC_OUT_BOT cbx_2__2_/SC_OUT_TOP VGND VPWR cbx_2__2_/bottom_grid_pin_0_
+ cbx_2__2_/bottom_grid_pin_10_ cbx_2__2_/bottom_grid_pin_11_ cbx_2__2_/bottom_grid_pin_12_
+ cbx_2__2_/bottom_grid_pin_13_ cbx_2__2_/bottom_grid_pin_14_ cbx_2__2_/bottom_grid_pin_15_
+ cbx_2__2_/bottom_grid_pin_1_ cbx_2__2_/bottom_grid_pin_2_ cbx_2__2_/bottom_grid_pin_3_
+ cbx_2__2_/bottom_grid_pin_4_ cbx_2__2_/bottom_grid_pin_5_ cbx_2__2_/bottom_grid_pin_6_
+ cbx_2__2_/bottom_grid_pin_7_ cbx_2__2_/bottom_grid_pin_8_ cbx_2__2_/bottom_grid_pin_9_
+ sb_2__2_/ccff_tail sb_1__2_/ccff_head cbx_2__2_/chanx_left_in[0] cbx_2__2_/chanx_left_in[10]
+ cbx_2__2_/chanx_left_in[11] cbx_2__2_/chanx_left_in[12] cbx_2__2_/chanx_left_in[13]
+ cbx_2__2_/chanx_left_in[14] cbx_2__2_/chanx_left_in[15] cbx_2__2_/chanx_left_in[16]
+ cbx_2__2_/chanx_left_in[17] cbx_2__2_/chanx_left_in[18] cbx_2__2_/chanx_left_in[19]
+ cbx_2__2_/chanx_left_in[1] cbx_2__2_/chanx_left_in[2] cbx_2__2_/chanx_left_in[3]
+ cbx_2__2_/chanx_left_in[4] cbx_2__2_/chanx_left_in[5] cbx_2__2_/chanx_left_in[6]
+ cbx_2__2_/chanx_left_in[7] cbx_2__2_/chanx_left_in[8] cbx_2__2_/chanx_left_in[9]
+ sb_1__2_/chanx_right_in[0] sb_1__2_/chanx_right_in[10] sb_1__2_/chanx_right_in[11]
+ sb_1__2_/chanx_right_in[12] sb_1__2_/chanx_right_in[13] sb_1__2_/chanx_right_in[14]
+ sb_1__2_/chanx_right_in[15] sb_1__2_/chanx_right_in[16] sb_1__2_/chanx_right_in[17]
+ sb_1__2_/chanx_right_in[18] sb_1__2_/chanx_right_in[19] sb_1__2_/chanx_right_in[1]
+ sb_1__2_/chanx_right_in[2] sb_1__2_/chanx_right_in[3] sb_1__2_/chanx_right_in[4]
+ sb_1__2_/chanx_right_in[5] sb_1__2_/chanx_right_in[6] sb_1__2_/chanx_right_in[7]
+ sb_1__2_/chanx_right_in[8] sb_1__2_/chanx_right_in[9] sb_2__2_/chanx_left_out[0]
+ sb_2__2_/chanx_left_out[10] sb_2__2_/chanx_left_out[11] sb_2__2_/chanx_left_out[12]
+ sb_2__2_/chanx_left_out[13] sb_2__2_/chanx_left_out[14] sb_2__2_/chanx_left_out[15]
+ sb_2__2_/chanx_left_out[16] sb_2__2_/chanx_left_out[17] sb_2__2_/chanx_left_out[18]
+ sb_2__2_/chanx_left_out[19] sb_2__2_/chanx_left_out[1] sb_2__2_/chanx_left_out[2]
+ sb_2__2_/chanx_left_out[3] sb_2__2_/chanx_left_out[4] sb_2__2_/chanx_left_out[5]
+ sb_2__2_/chanx_left_out[6] sb_2__2_/chanx_left_out[7] sb_2__2_/chanx_left_out[8]
+ sb_2__2_/chanx_left_out[9] sb_2__2_/chanx_left_in[0] sb_2__2_/chanx_left_in[10]
+ sb_2__2_/chanx_left_in[11] sb_2__2_/chanx_left_in[12] sb_2__2_/chanx_left_in[13]
+ sb_2__2_/chanx_left_in[14] sb_2__2_/chanx_left_in[15] sb_2__2_/chanx_left_in[16]
+ sb_2__2_/chanx_left_in[17] sb_2__2_/chanx_left_in[18] sb_2__2_/chanx_left_in[19]
+ sb_2__2_/chanx_left_in[1] sb_2__2_/chanx_left_in[2] sb_2__2_/chanx_left_in[3] sb_2__2_/chanx_left_in[4]
+ sb_2__2_/chanx_left_in[5] sb_2__2_/chanx_left_in[6] sb_2__2_/chanx_left_in[7] sb_2__2_/chanx_left_in[8]
+ sb_2__2_/chanx_left_in[9] cbx_2__2_/clk_1_N_out cbx_2__2_/clk_1_S_out cbx_2__2_/clk_1_W_in
+ cbx_2__2_/clk_2_E_out sb_2__2_/clk_2_W_out sb_1__2_/clk_2_N_in cbx_2__2_/clk_3_E_out
+ cbx_2__2_/clk_3_W_in cbx_2__2_/clk_3_W_out cbx_2__2_/prog_clk_0_N_in cbx_2__2_/prog_clk_0_W_out
+ cbx_2__2_/prog_clk_1_N_out cbx_2__2_/prog_clk_1_S_out cbx_2__2_/prog_clk_1_W_in
+ cbx_2__2_/prog_clk_2_E_out sb_2__2_/prog_clk_2_W_out sb_1__2_/prog_clk_2_N_in cbx_2__2_/prog_clk_3_E_out
+ cbx_2__2_/prog_clk_3_W_in cbx_2__2_/prog_clk_3_W_out cbx_1__1_
Xsb_2__7_ sb_2__7_/Test_en_N_out sb_2__7_/Test_en_S_in VGND VPWR sb_2__7_/bottom_left_grid_pin_42_
+ sb_2__7_/bottom_left_grid_pin_43_ sb_2__7_/bottom_left_grid_pin_44_ sb_2__7_/bottom_left_grid_pin_45_
+ sb_2__7_/bottom_left_grid_pin_46_ sb_2__7_/bottom_left_grid_pin_47_ sb_2__7_/bottom_left_grid_pin_48_
+ sb_2__7_/bottom_left_grid_pin_49_ sb_2__7_/ccff_head sb_2__7_/ccff_tail sb_2__7_/chanx_left_in[0]
+ sb_2__7_/chanx_left_in[10] sb_2__7_/chanx_left_in[11] sb_2__7_/chanx_left_in[12]
+ sb_2__7_/chanx_left_in[13] sb_2__7_/chanx_left_in[14] sb_2__7_/chanx_left_in[15]
+ sb_2__7_/chanx_left_in[16] sb_2__7_/chanx_left_in[17] sb_2__7_/chanx_left_in[18]
+ sb_2__7_/chanx_left_in[19] sb_2__7_/chanx_left_in[1] sb_2__7_/chanx_left_in[2] sb_2__7_/chanx_left_in[3]
+ sb_2__7_/chanx_left_in[4] sb_2__7_/chanx_left_in[5] sb_2__7_/chanx_left_in[6] sb_2__7_/chanx_left_in[7]
+ sb_2__7_/chanx_left_in[8] sb_2__7_/chanx_left_in[9] sb_2__7_/chanx_left_out[0] sb_2__7_/chanx_left_out[10]
+ sb_2__7_/chanx_left_out[11] sb_2__7_/chanx_left_out[12] sb_2__7_/chanx_left_out[13]
+ sb_2__7_/chanx_left_out[14] sb_2__7_/chanx_left_out[15] sb_2__7_/chanx_left_out[16]
+ sb_2__7_/chanx_left_out[17] sb_2__7_/chanx_left_out[18] sb_2__7_/chanx_left_out[19]
+ sb_2__7_/chanx_left_out[1] sb_2__7_/chanx_left_out[2] sb_2__7_/chanx_left_out[3]
+ sb_2__7_/chanx_left_out[4] sb_2__7_/chanx_left_out[5] sb_2__7_/chanx_left_out[6]
+ sb_2__7_/chanx_left_out[7] sb_2__7_/chanx_left_out[8] sb_2__7_/chanx_left_out[9]
+ sb_2__7_/chanx_right_in[0] sb_2__7_/chanx_right_in[10] sb_2__7_/chanx_right_in[11]
+ sb_2__7_/chanx_right_in[12] sb_2__7_/chanx_right_in[13] sb_2__7_/chanx_right_in[14]
+ sb_2__7_/chanx_right_in[15] sb_2__7_/chanx_right_in[16] sb_2__7_/chanx_right_in[17]
+ sb_2__7_/chanx_right_in[18] sb_2__7_/chanx_right_in[19] sb_2__7_/chanx_right_in[1]
+ sb_2__7_/chanx_right_in[2] sb_2__7_/chanx_right_in[3] sb_2__7_/chanx_right_in[4]
+ sb_2__7_/chanx_right_in[5] sb_2__7_/chanx_right_in[6] sb_2__7_/chanx_right_in[7]
+ sb_2__7_/chanx_right_in[8] sb_2__7_/chanx_right_in[9] cbx_3__7_/chanx_left_in[0]
+ cbx_3__7_/chanx_left_in[10] cbx_3__7_/chanx_left_in[11] cbx_3__7_/chanx_left_in[12]
+ cbx_3__7_/chanx_left_in[13] cbx_3__7_/chanx_left_in[14] cbx_3__7_/chanx_left_in[15]
+ cbx_3__7_/chanx_left_in[16] cbx_3__7_/chanx_left_in[17] cbx_3__7_/chanx_left_in[18]
+ cbx_3__7_/chanx_left_in[19] cbx_3__7_/chanx_left_in[1] cbx_3__7_/chanx_left_in[2]
+ cbx_3__7_/chanx_left_in[3] cbx_3__7_/chanx_left_in[4] cbx_3__7_/chanx_left_in[5]
+ cbx_3__7_/chanx_left_in[6] cbx_3__7_/chanx_left_in[7] cbx_3__7_/chanx_left_in[8]
+ cbx_3__7_/chanx_left_in[9] cby_2__7_/chany_top_out[0] cby_2__7_/chany_top_out[10]
+ cby_2__7_/chany_top_out[11] cby_2__7_/chany_top_out[12] cby_2__7_/chany_top_out[13]
+ cby_2__7_/chany_top_out[14] cby_2__7_/chany_top_out[15] cby_2__7_/chany_top_out[16]
+ cby_2__7_/chany_top_out[17] cby_2__7_/chany_top_out[18] cby_2__7_/chany_top_out[19]
+ cby_2__7_/chany_top_out[1] cby_2__7_/chany_top_out[2] cby_2__7_/chany_top_out[3]
+ cby_2__7_/chany_top_out[4] cby_2__7_/chany_top_out[5] cby_2__7_/chany_top_out[6]
+ cby_2__7_/chany_top_out[7] cby_2__7_/chany_top_out[8] cby_2__7_/chany_top_out[9]
+ cby_2__7_/chany_top_in[0] cby_2__7_/chany_top_in[10] cby_2__7_/chany_top_in[11]
+ cby_2__7_/chany_top_in[12] cby_2__7_/chany_top_in[13] cby_2__7_/chany_top_in[14]
+ cby_2__7_/chany_top_in[15] cby_2__7_/chany_top_in[16] cby_2__7_/chany_top_in[17]
+ cby_2__7_/chany_top_in[18] cby_2__7_/chany_top_in[19] cby_2__7_/chany_top_in[1]
+ cby_2__7_/chany_top_in[2] cby_2__7_/chany_top_in[3] cby_2__7_/chany_top_in[4] cby_2__7_/chany_top_in[5]
+ cby_2__7_/chany_top_in[6] cby_2__7_/chany_top_in[7] cby_2__7_/chany_top_in[8] cby_2__7_/chany_top_in[9]
+ sb_2__7_/chany_top_in[0] sb_2__7_/chany_top_in[10] sb_2__7_/chany_top_in[11] sb_2__7_/chany_top_in[12]
+ sb_2__7_/chany_top_in[13] sb_2__7_/chany_top_in[14] sb_2__7_/chany_top_in[15] sb_2__7_/chany_top_in[16]
+ sb_2__7_/chany_top_in[17] sb_2__7_/chany_top_in[18] sb_2__7_/chany_top_in[19] sb_2__7_/chany_top_in[1]
+ sb_2__7_/chany_top_in[2] sb_2__7_/chany_top_in[3] sb_2__7_/chany_top_in[4] sb_2__7_/chany_top_in[5]
+ sb_2__7_/chany_top_in[6] sb_2__7_/chany_top_in[7] sb_2__7_/chany_top_in[8] sb_2__7_/chany_top_in[9]
+ sb_2__7_/chany_top_out[0] sb_2__7_/chany_top_out[10] sb_2__7_/chany_top_out[11]
+ sb_2__7_/chany_top_out[12] sb_2__7_/chany_top_out[13] sb_2__7_/chany_top_out[14]
+ sb_2__7_/chany_top_out[15] sb_2__7_/chany_top_out[16] sb_2__7_/chany_top_out[17]
+ sb_2__7_/chany_top_out[18] sb_2__7_/chany_top_out[19] sb_2__7_/chany_top_out[1]
+ sb_2__7_/chany_top_out[2] sb_2__7_/chany_top_out[3] sb_2__7_/chany_top_out[4] sb_2__7_/chany_top_out[5]
+ sb_2__7_/chany_top_out[6] sb_2__7_/chany_top_out[7] sb_2__7_/chany_top_out[8] sb_2__7_/chany_top_out[9]
+ sb_2__7_/clk_1_E_out sb_2__7_/clk_1_N_in sb_2__7_/clk_1_W_out sb_2__7_/clk_2_E_out
+ sb_2__7_/clk_2_N_in sb_2__7_/clk_2_N_out sb_2__7_/clk_2_S_out sb_2__7_/clk_2_W_out
+ sb_2__7_/clk_3_E_out sb_2__7_/clk_3_N_in sb_2__7_/clk_3_N_out sb_2__7_/clk_3_S_out
+ sb_2__7_/clk_3_W_out sb_2__7_/left_bottom_grid_pin_34_ sb_2__7_/left_bottom_grid_pin_35_
+ sb_2__7_/left_bottom_grid_pin_36_ sb_2__7_/left_bottom_grid_pin_37_ sb_2__7_/left_bottom_grid_pin_38_
+ sb_2__7_/left_bottom_grid_pin_39_ sb_2__7_/left_bottom_grid_pin_40_ sb_2__7_/left_bottom_grid_pin_41_
+ sb_2__7_/prog_clk_0_N_in sb_2__7_/prog_clk_1_E_out sb_2__7_/prog_clk_1_N_in sb_2__7_/prog_clk_1_W_out
+ sb_2__7_/prog_clk_2_E_out sb_2__7_/prog_clk_2_N_in sb_2__7_/prog_clk_2_N_out sb_2__7_/prog_clk_2_S_out
+ sb_2__7_/prog_clk_2_W_out sb_2__7_/prog_clk_3_E_out sb_2__7_/prog_clk_3_N_in sb_2__7_/prog_clk_3_N_out
+ sb_2__7_/prog_clk_3_S_out sb_2__7_/prog_clk_3_W_out sb_2__7_/right_bottom_grid_pin_34_
+ sb_2__7_/right_bottom_grid_pin_35_ sb_2__7_/right_bottom_grid_pin_36_ sb_2__7_/right_bottom_grid_pin_37_
+ sb_2__7_/right_bottom_grid_pin_38_ sb_2__7_/right_bottom_grid_pin_39_ sb_2__7_/right_bottom_grid_pin_40_
+ sb_2__7_/right_bottom_grid_pin_41_ sb_2__7_/top_left_grid_pin_42_ sb_2__7_/top_left_grid_pin_43_
+ sb_2__7_/top_left_grid_pin_44_ sb_2__7_/top_left_grid_pin_45_ sb_2__7_/top_left_grid_pin_46_
+ sb_2__7_/top_left_grid_pin_47_ sb_2__7_/top_left_grid_pin_48_ sb_2__7_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_1__2_ cbx_1__2_/SC_OUT_BOT cbx_1__1_/SC_IN_TOP grid_clb_1__2_/SC_OUT_TOP
+ cby_1__2_/Test_en_W_out grid_clb_1__2_/Test_en_E_out cby_1__2_/Test_en_W_out grid_clb_1__2_/Test_en_W_out
+ VGND VPWR cbx_1__1_/REGIN_FEEDTHROUGH grid_clb_1__2_/bottom_width_0_height_0__pin_51_
+ cby_0__2_/ccff_tail cby_1__2_/ccff_head cbx_1__1_/clk_1_N_out cbx_1__1_/clk_1_N_out
+ cby_1__2_/prog_clk_0_W_in cbx_1__1_/prog_clk_1_N_out grid_clb_1__2_/prog_clk_0_N_out
+ cbx_1__1_/prog_clk_1_N_out cbx_1__1_/prog_clk_0_N_in cby_0__2_/prog_clk_0_E_in cby_1__2_/left_grid_pin_16_
+ cby_1__2_/left_grid_pin_17_ cby_1__2_/left_grid_pin_18_ cby_1__2_/left_grid_pin_19_
+ cby_1__2_/left_grid_pin_20_ cby_1__2_/left_grid_pin_21_ cby_1__2_/left_grid_pin_22_
+ cby_1__2_/left_grid_pin_23_ cby_1__2_/left_grid_pin_24_ cby_1__2_/left_grid_pin_25_
+ cby_1__2_/left_grid_pin_26_ cby_1__2_/left_grid_pin_27_ cby_1__2_/left_grid_pin_28_
+ cby_1__2_/left_grid_pin_29_ cby_1__2_/left_grid_pin_30_ cby_1__2_/left_grid_pin_31_
+ sb_1__1_/top_left_grid_pin_42_ sb_1__2_/bottom_left_grid_pin_42_ sb_1__1_/top_left_grid_pin_43_
+ sb_1__2_/bottom_left_grid_pin_43_ sb_1__1_/top_left_grid_pin_44_ sb_1__2_/bottom_left_grid_pin_44_
+ sb_1__1_/top_left_grid_pin_45_ sb_1__2_/bottom_left_grid_pin_45_ sb_1__1_/top_left_grid_pin_46_
+ sb_1__2_/bottom_left_grid_pin_46_ sb_1__1_/top_left_grid_pin_47_ sb_1__2_/bottom_left_grid_pin_47_
+ sb_1__1_/top_left_grid_pin_48_ sb_1__2_/bottom_left_grid_pin_48_ sb_1__1_/top_left_grid_pin_49_
+ sb_1__2_/bottom_left_grid_pin_49_ cbx_1__2_/bottom_grid_pin_0_ cbx_1__2_/bottom_grid_pin_10_
+ cbx_1__2_/bottom_grid_pin_11_ cbx_1__2_/bottom_grid_pin_12_ cbx_1__2_/bottom_grid_pin_13_
+ cbx_1__2_/bottom_grid_pin_14_ cbx_1__2_/bottom_grid_pin_15_ cbx_1__2_/bottom_grid_pin_1_
+ cbx_1__2_/bottom_grid_pin_2_ cbx_1__2_/REGOUT_FEEDTHROUGH grid_clb_1__2_/top_width_0_height_0__pin_33_
+ sb_1__2_/left_bottom_grid_pin_34_ sb_0__2_/right_bottom_grid_pin_34_ sb_1__2_/left_bottom_grid_pin_35_
+ sb_0__2_/right_bottom_grid_pin_35_ sb_1__2_/left_bottom_grid_pin_36_ sb_0__2_/right_bottom_grid_pin_36_
+ sb_1__2_/left_bottom_grid_pin_37_ sb_0__2_/right_bottom_grid_pin_37_ sb_1__2_/left_bottom_grid_pin_38_
+ sb_0__2_/right_bottom_grid_pin_38_ sb_1__2_/left_bottom_grid_pin_39_ sb_0__2_/right_bottom_grid_pin_39_
+ cbx_1__2_/bottom_grid_pin_3_ sb_1__2_/left_bottom_grid_pin_40_ sb_0__2_/right_bottom_grid_pin_40_
+ sb_1__2_/left_bottom_grid_pin_41_ sb_0__2_/right_bottom_grid_pin_41_ cbx_1__2_/bottom_grid_pin_4_
+ cbx_1__2_/bottom_grid_pin_5_ cbx_1__2_/bottom_grid_pin_6_ cbx_1__2_/bottom_grid_pin_7_
+ cbx_1__2_/bottom_grid_pin_8_ cbx_1__2_/bottom_grid_pin_9_ grid_clb
Xcby_8__6_ IO_ISOL_N VGND VPWR cby_8__6_/ccff_head sb_8__5_/ccff_head sb_8__5_/chany_top_out[0]
+ sb_8__5_/chany_top_out[10] sb_8__5_/chany_top_out[11] sb_8__5_/chany_top_out[12]
+ sb_8__5_/chany_top_out[13] sb_8__5_/chany_top_out[14] sb_8__5_/chany_top_out[15]
+ sb_8__5_/chany_top_out[16] sb_8__5_/chany_top_out[17] sb_8__5_/chany_top_out[18]
+ sb_8__5_/chany_top_out[19] sb_8__5_/chany_top_out[1] sb_8__5_/chany_top_out[2] sb_8__5_/chany_top_out[3]
+ sb_8__5_/chany_top_out[4] sb_8__5_/chany_top_out[5] sb_8__5_/chany_top_out[6] sb_8__5_/chany_top_out[7]
+ sb_8__5_/chany_top_out[8] sb_8__5_/chany_top_out[9] sb_8__5_/chany_top_in[0] sb_8__5_/chany_top_in[10]
+ sb_8__5_/chany_top_in[11] sb_8__5_/chany_top_in[12] sb_8__5_/chany_top_in[13] sb_8__5_/chany_top_in[14]
+ sb_8__5_/chany_top_in[15] sb_8__5_/chany_top_in[16] sb_8__5_/chany_top_in[17] sb_8__5_/chany_top_in[18]
+ sb_8__5_/chany_top_in[19] sb_8__5_/chany_top_in[1] sb_8__5_/chany_top_in[2] sb_8__5_/chany_top_in[3]
+ sb_8__5_/chany_top_in[4] sb_8__5_/chany_top_in[5] sb_8__5_/chany_top_in[6] sb_8__5_/chany_top_in[7]
+ sb_8__5_/chany_top_in[8] sb_8__5_/chany_top_in[9] cby_8__6_/chany_top_in[0] cby_8__6_/chany_top_in[10]
+ cby_8__6_/chany_top_in[11] cby_8__6_/chany_top_in[12] cby_8__6_/chany_top_in[13]
+ cby_8__6_/chany_top_in[14] cby_8__6_/chany_top_in[15] cby_8__6_/chany_top_in[16]
+ cby_8__6_/chany_top_in[17] cby_8__6_/chany_top_in[18] cby_8__6_/chany_top_in[19]
+ cby_8__6_/chany_top_in[1] cby_8__6_/chany_top_in[2] cby_8__6_/chany_top_in[3] cby_8__6_/chany_top_in[4]
+ cby_8__6_/chany_top_in[5] cby_8__6_/chany_top_in[6] cby_8__6_/chany_top_in[7] cby_8__6_/chany_top_in[8]
+ cby_8__6_/chany_top_in[9] cby_8__6_/chany_top_out[0] cby_8__6_/chany_top_out[10]
+ cby_8__6_/chany_top_out[11] cby_8__6_/chany_top_out[12] cby_8__6_/chany_top_out[13]
+ cby_8__6_/chany_top_out[14] cby_8__6_/chany_top_out[15] cby_8__6_/chany_top_out[16]
+ cby_8__6_/chany_top_out[17] cby_8__6_/chany_top_out[18] cby_8__6_/chany_top_out[19]
+ cby_8__6_/chany_top_out[1] cby_8__6_/chany_top_out[2] cby_8__6_/chany_top_out[3]
+ cby_8__6_/chany_top_out[4] cby_8__6_/chany_top_out[5] cby_8__6_/chany_top_out[6]
+ cby_8__6_/chany_top_out[7] cby_8__6_/chany_top_out[8] cby_8__6_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
+ cby_8__6_/left_grid_pin_16_ cby_8__6_/left_grid_pin_17_ cby_8__6_/left_grid_pin_18_
+ cby_8__6_/left_grid_pin_19_ cby_8__6_/left_grid_pin_20_ cby_8__6_/left_grid_pin_21_
+ cby_8__6_/left_grid_pin_22_ cby_8__6_/left_grid_pin_23_ cby_8__6_/left_grid_pin_24_
+ cby_8__6_/left_grid_pin_25_ cby_8__6_/left_grid_pin_26_ cby_8__6_/left_grid_pin_27_
+ cby_8__6_/left_grid_pin_28_ cby_8__6_/left_grid_pin_29_ cby_8__6_/left_grid_pin_30_
+ cby_8__6_/left_grid_pin_31_ cby_8__6_/right_grid_pin_0_ sb_8__5_/top_right_grid_pin_1_
+ sb_8__6_/bottom_right_grid_pin_1_ cby_8__6_/prog_clk_0_N_out sb_8__5_/prog_clk_0_N_in
+ cby_8__6_/prog_clk_0_W_in cby_8__6_/right_grid_pin_0_ cby_2__1_
Xcby_5__3_ cby_5__3_/Test_en_W_in cby_5__3_/Test_en_E_out cby_5__3_/Test_en_N_out
+ cby_5__3_/Test_en_W_in cby_5__3_/Test_en_W_in cby_5__3_/Test_en_W_out VGND VPWR
+ cby_5__3_/ccff_head cby_5__3_/ccff_tail sb_5__2_/chany_top_out[0] sb_5__2_/chany_top_out[10]
+ sb_5__2_/chany_top_out[11] sb_5__2_/chany_top_out[12] sb_5__2_/chany_top_out[13]
+ sb_5__2_/chany_top_out[14] sb_5__2_/chany_top_out[15] sb_5__2_/chany_top_out[16]
+ sb_5__2_/chany_top_out[17] sb_5__2_/chany_top_out[18] sb_5__2_/chany_top_out[19]
+ sb_5__2_/chany_top_out[1] sb_5__2_/chany_top_out[2] sb_5__2_/chany_top_out[3] sb_5__2_/chany_top_out[4]
+ sb_5__2_/chany_top_out[5] sb_5__2_/chany_top_out[6] sb_5__2_/chany_top_out[7] sb_5__2_/chany_top_out[8]
+ sb_5__2_/chany_top_out[9] sb_5__2_/chany_top_in[0] sb_5__2_/chany_top_in[10] sb_5__2_/chany_top_in[11]
+ sb_5__2_/chany_top_in[12] sb_5__2_/chany_top_in[13] sb_5__2_/chany_top_in[14] sb_5__2_/chany_top_in[15]
+ sb_5__2_/chany_top_in[16] sb_5__2_/chany_top_in[17] sb_5__2_/chany_top_in[18] sb_5__2_/chany_top_in[19]
+ sb_5__2_/chany_top_in[1] sb_5__2_/chany_top_in[2] sb_5__2_/chany_top_in[3] sb_5__2_/chany_top_in[4]
+ sb_5__2_/chany_top_in[5] sb_5__2_/chany_top_in[6] sb_5__2_/chany_top_in[7] sb_5__2_/chany_top_in[8]
+ sb_5__2_/chany_top_in[9] cby_5__3_/chany_top_in[0] cby_5__3_/chany_top_in[10] cby_5__3_/chany_top_in[11]
+ cby_5__3_/chany_top_in[12] cby_5__3_/chany_top_in[13] cby_5__3_/chany_top_in[14]
+ cby_5__3_/chany_top_in[15] cby_5__3_/chany_top_in[16] cby_5__3_/chany_top_in[17]
+ cby_5__3_/chany_top_in[18] cby_5__3_/chany_top_in[19] cby_5__3_/chany_top_in[1]
+ cby_5__3_/chany_top_in[2] cby_5__3_/chany_top_in[3] cby_5__3_/chany_top_in[4] cby_5__3_/chany_top_in[5]
+ cby_5__3_/chany_top_in[6] cby_5__3_/chany_top_in[7] cby_5__3_/chany_top_in[8] cby_5__3_/chany_top_in[9]
+ cby_5__3_/chany_top_out[0] cby_5__3_/chany_top_out[10] cby_5__3_/chany_top_out[11]
+ cby_5__3_/chany_top_out[12] cby_5__3_/chany_top_out[13] cby_5__3_/chany_top_out[14]
+ cby_5__3_/chany_top_out[15] cby_5__3_/chany_top_out[16] cby_5__3_/chany_top_out[17]
+ cby_5__3_/chany_top_out[18] cby_5__3_/chany_top_out[19] cby_5__3_/chany_top_out[1]
+ cby_5__3_/chany_top_out[2] cby_5__3_/chany_top_out[3] cby_5__3_/chany_top_out[4]
+ cby_5__3_/chany_top_out[5] cby_5__3_/chany_top_out[6] cby_5__3_/chany_top_out[7]
+ cby_5__3_/chany_top_out[8] cby_5__3_/chany_top_out[9] sb_5__3_/clk_1_N_in sb_5__2_/clk_2_N_out
+ cby_5__3_/clk_2_S_out cby_5__3_/clk_3_N_out cby_5__3_/clk_3_S_in cby_5__3_/clk_3_S_out
+ cby_5__3_/left_grid_pin_16_ cby_5__3_/left_grid_pin_17_ cby_5__3_/left_grid_pin_18_
+ cby_5__3_/left_grid_pin_19_ cby_5__3_/left_grid_pin_20_ cby_5__3_/left_grid_pin_21_
+ cby_5__3_/left_grid_pin_22_ cby_5__3_/left_grid_pin_23_ cby_5__3_/left_grid_pin_24_
+ cby_5__3_/left_grid_pin_25_ cby_5__3_/left_grid_pin_26_ cby_5__3_/left_grid_pin_27_
+ cby_5__3_/left_grid_pin_28_ cby_5__3_/left_grid_pin_29_ cby_5__3_/left_grid_pin_30_
+ cby_5__3_/left_grid_pin_31_ cby_5__3_/prog_clk_0_N_out sb_5__2_/prog_clk_0_N_in
+ cby_5__3_/prog_clk_0_W_in sb_5__3_/prog_clk_1_N_in sb_5__2_/prog_clk_2_N_out cby_5__3_/prog_clk_2_S_out
+ cby_5__3_/prog_clk_3_N_out cby_5__3_/prog_clk_3_S_in cby_5__3_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_8__7_ cbx_8__7_/REGIN_FEEDTHROUGH cbx_8__7_/REGOUT_FEEDTHROUGH cbx_8__7_/SC_IN_BOT
+ cbx_8__7_/SC_IN_TOP cbx_8__7_/SC_OUT_BOT cbx_8__7_/SC_OUT_TOP VGND VPWR cbx_8__7_/bottom_grid_pin_0_
+ cbx_8__7_/bottom_grid_pin_10_ cbx_8__7_/bottom_grid_pin_11_ cbx_8__7_/bottom_grid_pin_12_
+ cbx_8__7_/bottom_grid_pin_13_ cbx_8__7_/bottom_grid_pin_14_ cbx_8__7_/bottom_grid_pin_15_
+ cbx_8__7_/bottom_grid_pin_1_ cbx_8__7_/bottom_grid_pin_2_ cbx_8__7_/bottom_grid_pin_3_
+ cbx_8__7_/bottom_grid_pin_4_ cbx_8__7_/bottom_grid_pin_5_ cbx_8__7_/bottom_grid_pin_6_
+ cbx_8__7_/bottom_grid_pin_7_ cbx_8__7_/bottom_grid_pin_8_ cbx_8__7_/bottom_grid_pin_9_
+ sb_8__7_/ccff_tail sb_7__7_/ccff_head cbx_8__7_/chanx_left_in[0] cbx_8__7_/chanx_left_in[10]
+ cbx_8__7_/chanx_left_in[11] cbx_8__7_/chanx_left_in[12] cbx_8__7_/chanx_left_in[13]
+ cbx_8__7_/chanx_left_in[14] cbx_8__7_/chanx_left_in[15] cbx_8__7_/chanx_left_in[16]
+ cbx_8__7_/chanx_left_in[17] cbx_8__7_/chanx_left_in[18] cbx_8__7_/chanx_left_in[19]
+ cbx_8__7_/chanx_left_in[1] cbx_8__7_/chanx_left_in[2] cbx_8__7_/chanx_left_in[3]
+ cbx_8__7_/chanx_left_in[4] cbx_8__7_/chanx_left_in[5] cbx_8__7_/chanx_left_in[6]
+ cbx_8__7_/chanx_left_in[7] cbx_8__7_/chanx_left_in[8] cbx_8__7_/chanx_left_in[9]
+ sb_7__7_/chanx_right_in[0] sb_7__7_/chanx_right_in[10] sb_7__7_/chanx_right_in[11]
+ sb_7__7_/chanx_right_in[12] sb_7__7_/chanx_right_in[13] sb_7__7_/chanx_right_in[14]
+ sb_7__7_/chanx_right_in[15] sb_7__7_/chanx_right_in[16] sb_7__7_/chanx_right_in[17]
+ sb_7__7_/chanx_right_in[18] sb_7__7_/chanx_right_in[19] sb_7__7_/chanx_right_in[1]
+ sb_7__7_/chanx_right_in[2] sb_7__7_/chanx_right_in[3] sb_7__7_/chanx_right_in[4]
+ sb_7__7_/chanx_right_in[5] sb_7__7_/chanx_right_in[6] sb_7__7_/chanx_right_in[7]
+ sb_7__7_/chanx_right_in[8] sb_7__7_/chanx_right_in[9] sb_8__7_/chanx_left_out[0]
+ sb_8__7_/chanx_left_out[10] sb_8__7_/chanx_left_out[11] sb_8__7_/chanx_left_out[12]
+ sb_8__7_/chanx_left_out[13] sb_8__7_/chanx_left_out[14] sb_8__7_/chanx_left_out[15]
+ sb_8__7_/chanx_left_out[16] sb_8__7_/chanx_left_out[17] sb_8__7_/chanx_left_out[18]
+ sb_8__7_/chanx_left_out[19] sb_8__7_/chanx_left_out[1] sb_8__7_/chanx_left_out[2]
+ sb_8__7_/chanx_left_out[3] sb_8__7_/chanx_left_out[4] sb_8__7_/chanx_left_out[5]
+ sb_8__7_/chanx_left_out[6] sb_8__7_/chanx_left_out[7] sb_8__7_/chanx_left_out[8]
+ sb_8__7_/chanx_left_out[9] sb_8__7_/chanx_left_in[0] sb_8__7_/chanx_left_in[10]
+ sb_8__7_/chanx_left_in[11] sb_8__7_/chanx_left_in[12] sb_8__7_/chanx_left_in[13]
+ sb_8__7_/chanx_left_in[14] sb_8__7_/chanx_left_in[15] sb_8__7_/chanx_left_in[16]
+ sb_8__7_/chanx_left_in[17] sb_8__7_/chanx_left_in[18] sb_8__7_/chanx_left_in[19]
+ sb_8__7_/chanx_left_in[1] sb_8__7_/chanx_left_in[2] sb_8__7_/chanx_left_in[3] sb_8__7_/chanx_left_in[4]
+ sb_8__7_/chanx_left_in[5] sb_8__7_/chanx_left_in[6] sb_8__7_/chanx_left_in[7] sb_8__7_/chanx_left_in[8]
+ sb_8__7_/chanx_left_in[9] cbx_8__7_/clk_1_N_out cbx_8__7_/clk_1_S_out sb_7__7_/clk_1_E_out
+ cbx_8__7_/clk_2_E_out cbx_8__7_/clk_2_W_in cbx_8__7_/clk_2_W_out cbx_8__7_/clk_3_E_out
+ cbx_8__7_/clk_3_W_in cbx_8__7_/clk_3_W_out cbx_8__7_/prog_clk_0_N_in cbx_8__7_/prog_clk_0_W_out
+ cbx_8__7_/prog_clk_1_N_out cbx_8__7_/prog_clk_1_S_out sb_7__7_/prog_clk_1_E_out
+ cbx_8__7_/prog_clk_2_E_out cbx_8__7_/prog_clk_2_W_in cbx_8__7_/prog_clk_2_W_out
+ cbx_8__7_/prog_clk_3_E_out cbx_8__7_/prog_clk_3_W_in cbx_8__7_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_7__7_ cbx_7__7_/SC_OUT_BOT cbx_7__6_/SC_IN_TOP grid_clb_7__7_/SC_OUT_TOP
+ cby_6__7_/Test_en_E_out cby_7__7_/Test_en_W_in cby_6__7_/Test_en_E_out grid_clb_7__7_/Test_en_W_out
+ VGND VPWR cbx_7__6_/REGIN_FEEDTHROUGH grid_clb_7__7_/bottom_width_0_height_0__pin_51_
+ cby_6__7_/ccff_tail cby_7__7_/ccff_head cbx_7__7_/clk_1_S_out cbx_7__7_/clk_1_S_out
+ cby_7__7_/prog_clk_0_W_in cbx_7__7_/prog_clk_1_S_out grid_clb_7__7_/prog_clk_0_N_out
+ cbx_7__7_/prog_clk_1_S_out cbx_7__6_/prog_clk_0_N_in grid_clb_7__7_/prog_clk_0_W_out
+ cby_7__7_/left_grid_pin_16_ cby_7__7_/left_grid_pin_17_ cby_7__7_/left_grid_pin_18_
+ cby_7__7_/left_grid_pin_19_ cby_7__7_/left_grid_pin_20_ cby_7__7_/left_grid_pin_21_
+ cby_7__7_/left_grid_pin_22_ cby_7__7_/left_grid_pin_23_ cby_7__7_/left_grid_pin_24_
+ cby_7__7_/left_grid_pin_25_ cby_7__7_/left_grid_pin_26_ cby_7__7_/left_grid_pin_27_
+ cby_7__7_/left_grid_pin_28_ cby_7__7_/left_grid_pin_29_ cby_7__7_/left_grid_pin_30_
+ cby_7__7_/left_grid_pin_31_ sb_7__6_/top_left_grid_pin_42_ sb_7__7_/bottom_left_grid_pin_42_
+ sb_7__6_/top_left_grid_pin_43_ sb_7__7_/bottom_left_grid_pin_43_ sb_7__6_/top_left_grid_pin_44_
+ sb_7__7_/bottom_left_grid_pin_44_ sb_7__6_/top_left_grid_pin_45_ sb_7__7_/bottom_left_grid_pin_45_
+ sb_7__6_/top_left_grid_pin_46_ sb_7__7_/bottom_left_grid_pin_46_ sb_7__6_/top_left_grid_pin_47_
+ sb_7__7_/bottom_left_grid_pin_47_ sb_7__6_/top_left_grid_pin_48_ sb_7__7_/bottom_left_grid_pin_48_
+ sb_7__6_/top_left_grid_pin_49_ sb_7__7_/bottom_left_grid_pin_49_ cbx_7__7_/bottom_grid_pin_0_
+ cbx_7__7_/bottom_grid_pin_10_ cbx_7__7_/bottom_grid_pin_11_ cbx_7__7_/bottom_grid_pin_12_
+ cbx_7__7_/bottom_grid_pin_13_ cbx_7__7_/bottom_grid_pin_14_ cbx_7__7_/bottom_grid_pin_15_
+ cbx_7__7_/bottom_grid_pin_1_ cbx_7__7_/bottom_grid_pin_2_ cbx_7__7_/REGOUT_FEEDTHROUGH
+ grid_clb_7__7_/top_width_0_height_0__pin_33_ sb_7__7_/left_bottom_grid_pin_34_ sb_6__7_/right_bottom_grid_pin_34_
+ sb_7__7_/left_bottom_grid_pin_35_ sb_6__7_/right_bottom_grid_pin_35_ sb_7__7_/left_bottom_grid_pin_36_
+ sb_6__7_/right_bottom_grid_pin_36_ sb_7__7_/left_bottom_grid_pin_37_ sb_6__7_/right_bottom_grid_pin_37_
+ sb_7__7_/left_bottom_grid_pin_38_ sb_6__7_/right_bottom_grid_pin_38_ sb_7__7_/left_bottom_grid_pin_39_
+ sb_6__7_/right_bottom_grid_pin_39_ cbx_7__7_/bottom_grid_pin_3_ sb_7__7_/left_bottom_grid_pin_40_
+ sb_6__7_/right_bottom_grid_pin_40_ sb_7__7_/left_bottom_grid_pin_41_ sb_6__7_/right_bottom_grid_pin_41_
+ cbx_7__7_/bottom_grid_pin_4_ cbx_7__7_/bottom_grid_pin_5_ cbx_7__7_/bottom_grid_pin_6_
+ cbx_7__7_/bottom_grid_pin_7_ cbx_7__7_/bottom_grid_pin_8_ cbx_7__7_/bottom_grid_pin_9_
+ grid_clb
Xcbx_5__4_ cbx_5__4_/REGIN_FEEDTHROUGH cbx_5__4_/REGOUT_FEEDTHROUGH cbx_5__4_/SC_IN_BOT
+ cbx_5__4_/SC_IN_TOP cbx_5__4_/SC_OUT_BOT cbx_5__4_/SC_OUT_TOP VGND VPWR cbx_5__4_/bottom_grid_pin_0_
+ cbx_5__4_/bottom_grid_pin_10_ cbx_5__4_/bottom_grid_pin_11_ cbx_5__4_/bottom_grid_pin_12_
+ cbx_5__4_/bottom_grid_pin_13_ cbx_5__4_/bottom_grid_pin_14_ cbx_5__4_/bottom_grid_pin_15_
+ cbx_5__4_/bottom_grid_pin_1_ cbx_5__4_/bottom_grid_pin_2_ cbx_5__4_/bottom_grid_pin_3_
+ cbx_5__4_/bottom_grid_pin_4_ cbx_5__4_/bottom_grid_pin_5_ cbx_5__4_/bottom_grid_pin_6_
+ cbx_5__4_/bottom_grid_pin_7_ cbx_5__4_/bottom_grid_pin_8_ cbx_5__4_/bottom_grid_pin_9_
+ sb_5__4_/ccff_tail sb_4__4_/ccff_head cbx_5__4_/chanx_left_in[0] cbx_5__4_/chanx_left_in[10]
+ cbx_5__4_/chanx_left_in[11] cbx_5__4_/chanx_left_in[12] cbx_5__4_/chanx_left_in[13]
+ cbx_5__4_/chanx_left_in[14] cbx_5__4_/chanx_left_in[15] cbx_5__4_/chanx_left_in[16]
+ cbx_5__4_/chanx_left_in[17] cbx_5__4_/chanx_left_in[18] cbx_5__4_/chanx_left_in[19]
+ cbx_5__4_/chanx_left_in[1] cbx_5__4_/chanx_left_in[2] cbx_5__4_/chanx_left_in[3]
+ cbx_5__4_/chanx_left_in[4] cbx_5__4_/chanx_left_in[5] cbx_5__4_/chanx_left_in[6]
+ cbx_5__4_/chanx_left_in[7] cbx_5__4_/chanx_left_in[8] cbx_5__4_/chanx_left_in[9]
+ sb_4__4_/chanx_right_in[0] sb_4__4_/chanx_right_in[10] sb_4__4_/chanx_right_in[11]
+ sb_4__4_/chanx_right_in[12] sb_4__4_/chanx_right_in[13] sb_4__4_/chanx_right_in[14]
+ sb_4__4_/chanx_right_in[15] sb_4__4_/chanx_right_in[16] sb_4__4_/chanx_right_in[17]
+ sb_4__4_/chanx_right_in[18] sb_4__4_/chanx_right_in[19] sb_4__4_/chanx_right_in[1]
+ sb_4__4_/chanx_right_in[2] sb_4__4_/chanx_right_in[3] sb_4__4_/chanx_right_in[4]
+ sb_4__4_/chanx_right_in[5] sb_4__4_/chanx_right_in[6] sb_4__4_/chanx_right_in[7]
+ sb_4__4_/chanx_right_in[8] sb_4__4_/chanx_right_in[9] sb_5__4_/chanx_left_out[0]
+ sb_5__4_/chanx_left_out[10] sb_5__4_/chanx_left_out[11] sb_5__4_/chanx_left_out[12]
+ sb_5__4_/chanx_left_out[13] sb_5__4_/chanx_left_out[14] sb_5__4_/chanx_left_out[15]
+ sb_5__4_/chanx_left_out[16] sb_5__4_/chanx_left_out[17] sb_5__4_/chanx_left_out[18]
+ sb_5__4_/chanx_left_out[19] sb_5__4_/chanx_left_out[1] sb_5__4_/chanx_left_out[2]
+ sb_5__4_/chanx_left_out[3] sb_5__4_/chanx_left_out[4] sb_5__4_/chanx_left_out[5]
+ sb_5__4_/chanx_left_out[6] sb_5__4_/chanx_left_out[7] sb_5__4_/chanx_left_out[8]
+ sb_5__4_/chanx_left_out[9] sb_5__4_/chanx_left_in[0] sb_5__4_/chanx_left_in[10]
+ sb_5__4_/chanx_left_in[11] sb_5__4_/chanx_left_in[12] sb_5__4_/chanx_left_in[13]
+ sb_5__4_/chanx_left_in[14] sb_5__4_/chanx_left_in[15] sb_5__4_/chanx_left_in[16]
+ sb_5__4_/chanx_left_in[17] sb_5__4_/chanx_left_in[18] sb_5__4_/chanx_left_in[19]
+ sb_5__4_/chanx_left_in[1] sb_5__4_/chanx_left_in[2] sb_5__4_/chanx_left_in[3] sb_5__4_/chanx_left_in[4]
+ sb_5__4_/chanx_left_in[5] sb_5__4_/chanx_left_in[6] sb_5__4_/chanx_left_in[7] sb_5__4_/chanx_left_in[8]
+ sb_5__4_/chanx_left_in[9] cbx_5__4_/clk_1_N_out cbx_5__4_/clk_1_S_out cbx_5__4_/clk_1_W_in
+ cbx_5__4_/clk_2_E_out cbx_5__4_/clk_2_W_in cbx_5__4_/clk_2_W_out sb_5__4_/clk_3_N_in
+ sb_4__4_/clk_3_E_out cbx_5__4_/clk_3_W_out cbx_5__4_/prog_clk_0_N_in cbx_5__4_/prog_clk_0_W_out
+ cbx_5__4_/prog_clk_1_N_out cbx_5__4_/prog_clk_1_S_out cbx_5__4_/prog_clk_1_W_in
+ cbx_5__4_/prog_clk_2_E_out cbx_5__4_/prog_clk_2_W_in cbx_5__4_/prog_clk_2_W_out
+ sb_5__4_/prog_clk_3_N_in sb_4__4_/prog_clk_3_E_out cbx_5__4_/prog_clk_3_W_out cbx_1__1_
Xsb_2__6_ sb_2__6_/Test_en_N_out sb_2__6_/Test_en_S_in VGND VPWR sb_2__6_/bottom_left_grid_pin_42_
+ sb_2__6_/bottom_left_grid_pin_43_ sb_2__6_/bottom_left_grid_pin_44_ sb_2__6_/bottom_left_grid_pin_45_
+ sb_2__6_/bottom_left_grid_pin_46_ sb_2__6_/bottom_left_grid_pin_47_ sb_2__6_/bottom_left_grid_pin_48_
+ sb_2__6_/bottom_left_grid_pin_49_ sb_2__6_/ccff_head sb_2__6_/ccff_tail sb_2__6_/chanx_left_in[0]
+ sb_2__6_/chanx_left_in[10] sb_2__6_/chanx_left_in[11] sb_2__6_/chanx_left_in[12]
+ sb_2__6_/chanx_left_in[13] sb_2__6_/chanx_left_in[14] sb_2__6_/chanx_left_in[15]
+ sb_2__6_/chanx_left_in[16] sb_2__6_/chanx_left_in[17] sb_2__6_/chanx_left_in[18]
+ sb_2__6_/chanx_left_in[19] sb_2__6_/chanx_left_in[1] sb_2__6_/chanx_left_in[2] sb_2__6_/chanx_left_in[3]
+ sb_2__6_/chanx_left_in[4] sb_2__6_/chanx_left_in[5] sb_2__6_/chanx_left_in[6] sb_2__6_/chanx_left_in[7]
+ sb_2__6_/chanx_left_in[8] sb_2__6_/chanx_left_in[9] sb_2__6_/chanx_left_out[0] sb_2__6_/chanx_left_out[10]
+ sb_2__6_/chanx_left_out[11] sb_2__6_/chanx_left_out[12] sb_2__6_/chanx_left_out[13]
+ sb_2__6_/chanx_left_out[14] sb_2__6_/chanx_left_out[15] sb_2__6_/chanx_left_out[16]
+ sb_2__6_/chanx_left_out[17] sb_2__6_/chanx_left_out[18] sb_2__6_/chanx_left_out[19]
+ sb_2__6_/chanx_left_out[1] sb_2__6_/chanx_left_out[2] sb_2__6_/chanx_left_out[3]
+ sb_2__6_/chanx_left_out[4] sb_2__6_/chanx_left_out[5] sb_2__6_/chanx_left_out[6]
+ sb_2__6_/chanx_left_out[7] sb_2__6_/chanx_left_out[8] sb_2__6_/chanx_left_out[9]
+ sb_2__6_/chanx_right_in[0] sb_2__6_/chanx_right_in[10] sb_2__6_/chanx_right_in[11]
+ sb_2__6_/chanx_right_in[12] sb_2__6_/chanx_right_in[13] sb_2__6_/chanx_right_in[14]
+ sb_2__6_/chanx_right_in[15] sb_2__6_/chanx_right_in[16] sb_2__6_/chanx_right_in[17]
+ sb_2__6_/chanx_right_in[18] sb_2__6_/chanx_right_in[19] sb_2__6_/chanx_right_in[1]
+ sb_2__6_/chanx_right_in[2] sb_2__6_/chanx_right_in[3] sb_2__6_/chanx_right_in[4]
+ sb_2__6_/chanx_right_in[5] sb_2__6_/chanx_right_in[6] sb_2__6_/chanx_right_in[7]
+ sb_2__6_/chanx_right_in[8] sb_2__6_/chanx_right_in[9] cbx_3__6_/chanx_left_in[0]
+ cbx_3__6_/chanx_left_in[10] cbx_3__6_/chanx_left_in[11] cbx_3__6_/chanx_left_in[12]
+ cbx_3__6_/chanx_left_in[13] cbx_3__6_/chanx_left_in[14] cbx_3__6_/chanx_left_in[15]
+ cbx_3__6_/chanx_left_in[16] cbx_3__6_/chanx_left_in[17] cbx_3__6_/chanx_left_in[18]
+ cbx_3__6_/chanx_left_in[19] cbx_3__6_/chanx_left_in[1] cbx_3__6_/chanx_left_in[2]
+ cbx_3__6_/chanx_left_in[3] cbx_3__6_/chanx_left_in[4] cbx_3__6_/chanx_left_in[5]
+ cbx_3__6_/chanx_left_in[6] cbx_3__6_/chanx_left_in[7] cbx_3__6_/chanx_left_in[8]
+ cbx_3__6_/chanx_left_in[9] cby_2__6_/chany_top_out[0] cby_2__6_/chany_top_out[10]
+ cby_2__6_/chany_top_out[11] cby_2__6_/chany_top_out[12] cby_2__6_/chany_top_out[13]
+ cby_2__6_/chany_top_out[14] cby_2__6_/chany_top_out[15] cby_2__6_/chany_top_out[16]
+ cby_2__6_/chany_top_out[17] cby_2__6_/chany_top_out[18] cby_2__6_/chany_top_out[19]
+ cby_2__6_/chany_top_out[1] cby_2__6_/chany_top_out[2] cby_2__6_/chany_top_out[3]
+ cby_2__6_/chany_top_out[4] cby_2__6_/chany_top_out[5] cby_2__6_/chany_top_out[6]
+ cby_2__6_/chany_top_out[7] cby_2__6_/chany_top_out[8] cby_2__6_/chany_top_out[9]
+ cby_2__6_/chany_top_in[0] cby_2__6_/chany_top_in[10] cby_2__6_/chany_top_in[11]
+ cby_2__6_/chany_top_in[12] cby_2__6_/chany_top_in[13] cby_2__6_/chany_top_in[14]
+ cby_2__6_/chany_top_in[15] cby_2__6_/chany_top_in[16] cby_2__6_/chany_top_in[17]
+ cby_2__6_/chany_top_in[18] cby_2__6_/chany_top_in[19] cby_2__6_/chany_top_in[1]
+ cby_2__6_/chany_top_in[2] cby_2__6_/chany_top_in[3] cby_2__6_/chany_top_in[4] cby_2__6_/chany_top_in[5]
+ cby_2__6_/chany_top_in[6] cby_2__6_/chany_top_in[7] cby_2__6_/chany_top_in[8] cby_2__6_/chany_top_in[9]
+ sb_2__6_/chany_top_in[0] sb_2__6_/chany_top_in[10] sb_2__6_/chany_top_in[11] sb_2__6_/chany_top_in[12]
+ sb_2__6_/chany_top_in[13] sb_2__6_/chany_top_in[14] sb_2__6_/chany_top_in[15] sb_2__6_/chany_top_in[16]
+ sb_2__6_/chany_top_in[17] sb_2__6_/chany_top_in[18] sb_2__6_/chany_top_in[19] sb_2__6_/chany_top_in[1]
+ sb_2__6_/chany_top_in[2] sb_2__6_/chany_top_in[3] sb_2__6_/chany_top_in[4] sb_2__6_/chany_top_in[5]
+ sb_2__6_/chany_top_in[6] sb_2__6_/chany_top_in[7] sb_2__6_/chany_top_in[8] sb_2__6_/chany_top_in[9]
+ sb_2__6_/chany_top_out[0] sb_2__6_/chany_top_out[10] sb_2__6_/chany_top_out[11]
+ sb_2__6_/chany_top_out[12] sb_2__6_/chany_top_out[13] sb_2__6_/chany_top_out[14]
+ sb_2__6_/chany_top_out[15] sb_2__6_/chany_top_out[16] sb_2__6_/chany_top_out[17]
+ sb_2__6_/chany_top_out[18] sb_2__6_/chany_top_out[19] sb_2__6_/chany_top_out[1]
+ sb_2__6_/chany_top_out[2] sb_2__6_/chany_top_out[3] sb_2__6_/chany_top_out[4] sb_2__6_/chany_top_out[5]
+ sb_2__6_/chany_top_out[6] sb_2__6_/chany_top_out[7] sb_2__6_/chany_top_out[8] sb_2__6_/chany_top_out[9]
+ sb_2__6_/clk_1_E_out sb_2__6_/clk_1_N_in sb_2__6_/clk_1_W_out sb_2__6_/clk_2_E_out
+ sb_2__6_/clk_2_N_in sb_2__6_/clk_2_N_out sb_2__6_/clk_2_S_out sb_2__6_/clk_2_W_out
+ sb_2__6_/clk_3_E_out sb_2__6_/clk_3_N_in sb_2__6_/clk_3_N_out sb_2__6_/clk_3_S_out
+ sb_2__6_/clk_3_W_out sb_2__6_/left_bottom_grid_pin_34_ sb_2__6_/left_bottom_grid_pin_35_
+ sb_2__6_/left_bottom_grid_pin_36_ sb_2__6_/left_bottom_grid_pin_37_ sb_2__6_/left_bottom_grid_pin_38_
+ sb_2__6_/left_bottom_grid_pin_39_ sb_2__6_/left_bottom_grid_pin_40_ sb_2__6_/left_bottom_grid_pin_41_
+ sb_2__6_/prog_clk_0_N_in sb_2__6_/prog_clk_1_E_out sb_2__6_/prog_clk_1_N_in sb_2__6_/prog_clk_1_W_out
+ sb_2__6_/prog_clk_2_E_out sb_2__6_/prog_clk_2_N_in sb_2__6_/prog_clk_2_N_out sb_2__6_/prog_clk_2_S_out
+ sb_2__6_/prog_clk_2_W_out sb_2__6_/prog_clk_3_E_out sb_2__6_/prog_clk_3_N_in sb_2__6_/prog_clk_3_N_out
+ sb_2__6_/prog_clk_3_S_out sb_2__6_/prog_clk_3_W_out sb_2__6_/right_bottom_grid_pin_34_
+ sb_2__6_/right_bottom_grid_pin_35_ sb_2__6_/right_bottom_grid_pin_36_ sb_2__6_/right_bottom_grid_pin_37_
+ sb_2__6_/right_bottom_grid_pin_38_ sb_2__6_/right_bottom_grid_pin_39_ sb_2__6_/right_bottom_grid_pin_40_
+ sb_2__6_/right_bottom_grid_pin_41_ sb_2__6_/top_left_grid_pin_42_ sb_2__6_/top_left_grid_pin_43_
+ sb_2__6_/top_left_grid_pin_44_ sb_2__6_/top_left_grid_pin_45_ sb_2__6_/top_left_grid_pin_46_
+ sb_2__6_/top_left_grid_pin_47_ sb_2__6_/top_left_grid_pin_48_ sb_2__6_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_4__4_ cbx_4__3_/SC_OUT_TOP grid_clb_4__4_/SC_OUT_BOT cbx_4__4_/SC_IN_BOT
+ cby_4__4_/Test_en_W_out grid_clb_4__4_/Test_en_E_out cby_4__4_/Test_en_W_out cby_3__4_/Test_en_W_in
+ VGND VPWR cbx_4__3_/REGIN_FEEDTHROUGH grid_clb_4__4_/bottom_width_0_height_0__pin_51_
+ cby_3__4_/ccff_tail cby_4__4_/ccff_head cbx_4__3_/clk_1_N_out cbx_4__3_/clk_1_N_out
+ cby_4__4_/prog_clk_0_W_in cbx_4__3_/prog_clk_1_N_out grid_clb_4__4_/prog_clk_0_N_out
+ cbx_4__3_/prog_clk_1_N_out cbx_4__3_/prog_clk_0_N_in grid_clb_4__4_/prog_clk_0_W_out
+ cby_4__4_/left_grid_pin_16_ cby_4__4_/left_grid_pin_17_ cby_4__4_/left_grid_pin_18_
+ cby_4__4_/left_grid_pin_19_ cby_4__4_/left_grid_pin_20_ cby_4__4_/left_grid_pin_21_
+ cby_4__4_/left_grid_pin_22_ cby_4__4_/left_grid_pin_23_ cby_4__4_/left_grid_pin_24_
+ cby_4__4_/left_grid_pin_25_ cby_4__4_/left_grid_pin_26_ cby_4__4_/left_grid_pin_27_
+ cby_4__4_/left_grid_pin_28_ cby_4__4_/left_grid_pin_29_ cby_4__4_/left_grid_pin_30_
+ cby_4__4_/left_grid_pin_31_ sb_4__3_/top_left_grid_pin_42_ sb_4__4_/bottom_left_grid_pin_42_
+ sb_4__3_/top_left_grid_pin_43_ sb_4__4_/bottom_left_grid_pin_43_ sb_4__3_/top_left_grid_pin_44_
+ sb_4__4_/bottom_left_grid_pin_44_ sb_4__3_/top_left_grid_pin_45_ sb_4__4_/bottom_left_grid_pin_45_
+ sb_4__3_/top_left_grid_pin_46_ sb_4__4_/bottom_left_grid_pin_46_ sb_4__3_/top_left_grid_pin_47_
+ sb_4__4_/bottom_left_grid_pin_47_ sb_4__3_/top_left_grid_pin_48_ sb_4__4_/bottom_left_grid_pin_48_
+ sb_4__3_/top_left_grid_pin_49_ sb_4__4_/bottom_left_grid_pin_49_ cbx_4__4_/bottom_grid_pin_0_
+ cbx_4__4_/bottom_grid_pin_10_ cbx_4__4_/bottom_grid_pin_11_ cbx_4__4_/bottom_grid_pin_12_
+ cbx_4__4_/bottom_grid_pin_13_ cbx_4__4_/bottom_grid_pin_14_ cbx_4__4_/bottom_grid_pin_15_
+ cbx_4__4_/bottom_grid_pin_1_ cbx_4__4_/bottom_grid_pin_2_ cbx_4__4_/REGOUT_FEEDTHROUGH
+ grid_clb_4__4_/top_width_0_height_0__pin_33_ sb_4__4_/left_bottom_grid_pin_34_ sb_3__4_/right_bottom_grid_pin_34_
+ sb_4__4_/left_bottom_grid_pin_35_ sb_3__4_/right_bottom_grid_pin_35_ sb_4__4_/left_bottom_grid_pin_36_
+ sb_3__4_/right_bottom_grid_pin_36_ sb_4__4_/left_bottom_grid_pin_37_ sb_3__4_/right_bottom_grid_pin_37_
+ sb_4__4_/left_bottom_grid_pin_38_ sb_3__4_/right_bottom_grid_pin_38_ sb_4__4_/left_bottom_grid_pin_39_
+ sb_3__4_/right_bottom_grid_pin_39_ cbx_4__4_/bottom_grid_pin_3_ sb_4__4_/left_bottom_grid_pin_40_
+ sb_3__4_/right_bottom_grid_pin_40_ sb_4__4_/left_bottom_grid_pin_41_ sb_3__4_/right_bottom_grid_pin_41_
+ cbx_4__4_/bottom_grid_pin_4_ cbx_4__4_/bottom_grid_pin_5_ cbx_4__4_/bottom_grid_pin_6_
+ cbx_4__4_/bottom_grid_pin_7_ cbx_4__4_/bottom_grid_pin_8_ cbx_4__4_/bottom_grid_pin_9_
+ grid_clb
Xgrid_clb_1__1_ cbx_1__1_/SC_OUT_BOT cbx_1__0_/SC_IN_TOP grid_clb_1__1_/SC_OUT_TOP
+ cby_1__1_/Test_en_W_out grid_clb_1__1_/Test_en_E_out cby_1__1_/Test_en_W_out grid_clb_1__1_/Test_en_W_out
+ VGND VPWR grid_clb_1__1_/bottom_width_0_height_0__pin_50_ grid_clb_1__1_/bottom_width_0_height_0__pin_51_
+ cby_0__1_/ccff_tail cby_1__1_/ccff_head cbx_1__1_/clk_1_S_out cbx_1__1_/clk_1_S_out
+ cby_1__1_/prog_clk_0_W_in cbx_1__1_/prog_clk_1_S_out grid_clb_1__1_/prog_clk_0_N_out
+ cbx_1__1_/prog_clk_1_S_out cbx_1__0_/prog_clk_0_N_in cby_0__1_/prog_clk_0_E_in cby_1__1_/left_grid_pin_16_
+ cby_1__1_/left_grid_pin_17_ cby_1__1_/left_grid_pin_18_ cby_1__1_/left_grid_pin_19_
+ cby_1__1_/left_grid_pin_20_ cby_1__1_/left_grid_pin_21_ cby_1__1_/left_grid_pin_22_
+ cby_1__1_/left_grid_pin_23_ cby_1__1_/left_grid_pin_24_ cby_1__1_/left_grid_pin_25_
+ cby_1__1_/left_grid_pin_26_ cby_1__1_/left_grid_pin_27_ cby_1__1_/left_grid_pin_28_
+ cby_1__1_/left_grid_pin_29_ cby_1__1_/left_grid_pin_30_ cby_1__1_/left_grid_pin_31_
+ sb_1__0_/top_left_grid_pin_42_ sb_1__1_/bottom_left_grid_pin_42_ sb_1__0_/top_left_grid_pin_43_
+ sb_1__1_/bottom_left_grid_pin_43_ sb_1__0_/top_left_grid_pin_44_ sb_1__1_/bottom_left_grid_pin_44_
+ sb_1__0_/top_left_grid_pin_45_ sb_1__1_/bottom_left_grid_pin_45_ sb_1__0_/top_left_grid_pin_46_
+ sb_1__1_/bottom_left_grid_pin_46_ sb_1__0_/top_left_grid_pin_47_ sb_1__1_/bottom_left_grid_pin_47_
+ sb_1__0_/top_left_grid_pin_48_ sb_1__1_/bottom_left_grid_pin_48_ sb_1__0_/top_left_grid_pin_49_
+ sb_1__1_/bottom_left_grid_pin_49_ cbx_1__1_/bottom_grid_pin_0_ cbx_1__1_/bottom_grid_pin_10_
+ cbx_1__1_/bottom_grid_pin_11_ cbx_1__1_/bottom_grid_pin_12_ cbx_1__1_/bottom_grid_pin_13_
+ cbx_1__1_/bottom_grid_pin_14_ cbx_1__1_/bottom_grid_pin_15_ cbx_1__1_/bottom_grid_pin_1_
+ cbx_1__1_/bottom_grid_pin_2_ cbx_1__1_/REGOUT_FEEDTHROUGH grid_clb_1__1_/top_width_0_height_0__pin_33_
+ sb_1__1_/left_bottom_grid_pin_34_ sb_0__1_/right_bottom_grid_pin_34_ sb_1__1_/left_bottom_grid_pin_35_
+ sb_0__1_/right_bottom_grid_pin_35_ sb_1__1_/left_bottom_grid_pin_36_ sb_0__1_/right_bottom_grid_pin_36_
+ sb_1__1_/left_bottom_grid_pin_37_ sb_0__1_/right_bottom_grid_pin_37_ sb_1__1_/left_bottom_grid_pin_38_
+ sb_0__1_/right_bottom_grid_pin_38_ sb_1__1_/left_bottom_grid_pin_39_ sb_0__1_/right_bottom_grid_pin_39_
+ cbx_1__1_/bottom_grid_pin_3_ sb_1__1_/left_bottom_grid_pin_40_ sb_0__1_/right_bottom_grid_pin_40_
+ sb_1__1_/left_bottom_grid_pin_41_ sb_0__1_/right_bottom_grid_pin_41_ cbx_1__1_/bottom_grid_pin_4_
+ cbx_1__1_/bottom_grid_pin_5_ cbx_1__1_/bottom_grid_pin_6_ cbx_1__1_/bottom_grid_pin_7_
+ cbx_1__1_/bottom_grid_pin_8_ cbx_1__1_/bottom_grid_pin_9_ grid_clb
Xcbx_2__1_ cbx_2__1_/REGIN_FEEDTHROUGH cbx_2__1_/REGOUT_FEEDTHROUGH cbx_2__1_/SC_IN_BOT
+ cbx_2__1_/SC_IN_TOP cbx_2__1_/SC_OUT_BOT cbx_2__1_/SC_OUT_TOP VGND VPWR cbx_2__1_/bottom_grid_pin_0_
+ cbx_2__1_/bottom_grid_pin_10_ cbx_2__1_/bottom_grid_pin_11_ cbx_2__1_/bottom_grid_pin_12_
+ cbx_2__1_/bottom_grid_pin_13_ cbx_2__1_/bottom_grid_pin_14_ cbx_2__1_/bottom_grid_pin_15_
+ cbx_2__1_/bottom_grid_pin_1_ cbx_2__1_/bottom_grid_pin_2_ cbx_2__1_/bottom_grid_pin_3_
+ cbx_2__1_/bottom_grid_pin_4_ cbx_2__1_/bottom_grid_pin_5_ cbx_2__1_/bottom_grid_pin_6_
+ cbx_2__1_/bottom_grid_pin_7_ cbx_2__1_/bottom_grid_pin_8_ cbx_2__1_/bottom_grid_pin_9_
+ sb_2__1_/ccff_tail sb_1__1_/ccff_head cbx_2__1_/chanx_left_in[0] cbx_2__1_/chanx_left_in[10]
+ cbx_2__1_/chanx_left_in[11] cbx_2__1_/chanx_left_in[12] cbx_2__1_/chanx_left_in[13]
+ cbx_2__1_/chanx_left_in[14] cbx_2__1_/chanx_left_in[15] cbx_2__1_/chanx_left_in[16]
+ cbx_2__1_/chanx_left_in[17] cbx_2__1_/chanx_left_in[18] cbx_2__1_/chanx_left_in[19]
+ cbx_2__1_/chanx_left_in[1] cbx_2__1_/chanx_left_in[2] cbx_2__1_/chanx_left_in[3]
+ cbx_2__1_/chanx_left_in[4] cbx_2__1_/chanx_left_in[5] cbx_2__1_/chanx_left_in[6]
+ cbx_2__1_/chanx_left_in[7] cbx_2__1_/chanx_left_in[8] cbx_2__1_/chanx_left_in[9]
+ sb_1__1_/chanx_right_in[0] sb_1__1_/chanx_right_in[10] sb_1__1_/chanx_right_in[11]
+ sb_1__1_/chanx_right_in[12] sb_1__1_/chanx_right_in[13] sb_1__1_/chanx_right_in[14]
+ sb_1__1_/chanx_right_in[15] sb_1__1_/chanx_right_in[16] sb_1__1_/chanx_right_in[17]
+ sb_1__1_/chanx_right_in[18] sb_1__1_/chanx_right_in[19] sb_1__1_/chanx_right_in[1]
+ sb_1__1_/chanx_right_in[2] sb_1__1_/chanx_right_in[3] sb_1__1_/chanx_right_in[4]
+ sb_1__1_/chanx_right_in[5] sb_1__1_/chanx_right_in[6] sb_1__1_/chanx_right_in[7]
+ sb_1__1_/chanx_right_in[8] sb_1__1_/chanx_right_in[9] sb_2__1_/chanx_left_out[0]
+ sb_2__1_/chanx_left_out[10] sb_2__1_/chanx_left_out[11] sb_2__1_/chanx_left_out[12]
+ sb_2__1_/chanx_left_out[13] sb_2__1_/chanx_left_out[14] sb_2__1_/chanx_left_out[15]
+ sb_2__1_/chanx_left_out[16] sb_2__1_/chanx_left_out[17] sb_2__1_/chanx_left_out[18]
+ sb_2__1_/chanx_left_out[19] sb_2__1_/chanx_left_out[1] sb_2__1_/chanx_left_out[2]
+ sb_2__1_/chanx_left_out[3] sb_2__1_/chanx_left_out[4] sb_2__1_/chanx_left_out[5]
+ sb_2__1_/chanx_left_out[6] sb_2__1_/chanx_left_out[7] sb_2__1_/chanx_left_out[8]
+ sb_2__1_/chanx_left_out[9] sb_2__1_/chanx_left_in[0] sb_2__1_/chanx_left_in[10]
+ sb_2__1_/chanx_left_in[11] sb_2__1_/chanx_left_in[12] sb_2__1_/chanx_left_in[13]
+ sb_2__1_/chanx_left_in[14] sb_2__1_/chanx_left_in[15] sb_2__1_/chanx_left_in[16]
+ sb_2__1_/chanx_left_in[17] sb_2__1_/chanx_left_in[18] sb_2__1_/chanx_left_in[19]
+ sb_2__1_/chanx_left_in[1] sb_2__1_/chanx_left_in[2] sb_2__1_/chanx_left_in[3] sb_2__1_/chanx_left_in[4]
+ sb_2__1_/chanx_left_in[5] sb_2__1_/chanx_left_in[6] sb_2__1_/chanx_left_in[7] sb_2__1_/chanx_left_in[8]
+ sb_2__1_/chanx_left_in[9] cbx_2__1_/clk_1_N_out cbx_2__1_/clk_1_S_out sb_1__1_/clk_1_E_out
+ cbx_2__1_/clk_2_E_out cbx_2__1_/clk_2_W_in cbx_2__1_/clk_2_W_out cbx_2__1_/clk_3_E_out
+ cbx_2__1_/clk_3_W_in cbx_2__1_/clk_3_W_out cbx_2__1_/prog_clk_0_N_in cbx_2__1_/prog_clk_0_W_out
+ cbx_2__1_/prog_clk_1_N_out cbx_2__1_/prog_clk_1_S_out sb_1__1_/prog_clk_1_E_out
+ cbx_2__1_/prog_clk_2_E_out cbx_2__1_/prog_clk_2_W_in cbx_2__1_/prog_clk_2_W_out
+ cbx_2__1_/prog_clk_3_E_out cbx_2__1_/prog_clk_3_W_in cbx_2__1_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_8__5_ IO_ISOL_N VGND VPWR cby_8__5_/ccff_head sb_8__4_/ccff_head sb_8__4_/chany_top_out[0]
+ sb_8__4_/chany_top_out[10] sb_8__4_/chany_top_out[11] sb_8__4_/chany_top_out[12]
+ sb_8__4_/chany_top_out[13] sb_8__4_/chany_top_out[14] sb_8__4_/chany_top_out[15]
+ sb_8__4_/chany_top_out[16] sb_8__4_/chany_top_out[17] sb_8__4_/chany_top_out[18]
+ sb_8__4_/chany_top_out[19] sb_8__4_/chany_top_out[1] sb_8__4_/chany_top_out[2] sb_8__4_/chany_top_out[3]
+ sb_8__4_/chany_top_out[4] sb_8__4_/chany_top_out[5] sb_8__4_/chany_top_out[6] sb_8__4_/chany_top_out[7]
+ sb_8__4_/chany_top_out[8] sb_8__4_/chany_top_out[9] sb_8__4_/chany_top_in[0] sb_8__4_/chany_top_in[10]
+ sb_8__4_/chany_top_in[11] sb_8__4_/chany_top_in[12] sb_8__4_/chany_top_in[13] sb_8__4_/chany_top_in[14]
+ sb_8__4_/chany_top_in[15] sb_8__4_/chany_top_in[16] sb_8__4_/chany_top_in[17] sb_8__4_/chany_top_in[18]
+ sb_8__4_/chany_top_in[19] sb_8__4_/chany_top_in[1] sb_8__4_/chany_top_in[2] sb_8__4_/chany_top_in[3]
+ sb_8__4_/chany_top_in[4] sb_8__4_/chany_top_in[5] sb_8__4_/chany_top_in[6] sb_8__4_/chany_top_in[7]
+ sb_8__4_/chany_top_in[8] sb_8__4_/chany_top_in[9] cby_8__5_/chany_top_in[0] cby_8__5_/chany_top_in[10]
+ cby_8__5_/chany_top_in[11] cby_8__5_/chany_top_in[12] cby_8__5_/chany_top_in[13]
+ cby_8__5_/chany_top_in[14] cby_8__5_/chany_top_in[15] cby_8__5_/chany_top_in[16]
+ cby_8__5_/chany_top_in[17] cby_8__5_/chany_top_in[18] cby_8__5_/chany_top_in[19]
+ cby_8__5_/chany_top_in[1] cby_8__5_/chany_top_in[2] cby_8__5_/chany_top_in[3] cby_8__5_/chany_top_in[4]
+ cby_8__5_/chany_top_in[5] cby_8__5_/chany_top_in[6] cby_8__5_/chany_top_in[7] cby_8__5_/chany_top_in[8]
+ cby_8__5_/chany_top_in[9] cby_8__5_/chany_top_out[0] cby_8__5_/chany_top_out[10]
+ cby_8__5_/chany_top_out[11] cby_8__5_/chany_top_out[12] cby_8__5_/chany_top_out[13]
+ cby_8__5_/chany_top_out[14] cby_8__5_/chany_top_out[15] cby_8__5_/chany_top_out[16]
+ cby_8__5_/chany_top_out[17] cby_8__5_/chany_top_out[18] cby_8__5_/chany_top_out[19]
+ cby_8__5_/chany_top_out[1] cby_8__5_/chany_top_out[2] cby_8__5_/chany_top_out[3]
+ cby_8__5_/chany_top_out[4] cby_8__5_/chany_top_out[5] cby_8__5_/chany_top_out[6]
+ cby_8__5_/chany_top_out[7] cby_8__5_/chany_top_out[8] cby_8__5_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
+ cby_8__5_/left_grid_pin_16_ cby_8__5_/left_grid_pin_17_ cby_8__5_/left_grid_pin_18_
+ cby_8__5_/left_grid_pin_19_ cby_8__5_/left_grid_pin_20_ cby_8__5_/left_grid_pin_21_
+ cby_8__5_/left_grid_pin_22_ cby_8__5_/left_grid_pin_23_ cby_8__5_/left_grid_pin_24_
+ cby_8__5_/left_grid_pin_25_ cby_8__5_/left_grid_pin_26_ cby_8__5_/left_grid_pin_27_
+ cby_8__5_/left_grid_pin_28_ cby_8__5_/left_grid_pin_29_ cby_8__5_/left_grid_pin_30_
+ cby_8__5_/left_grid_pin_31_ cby_8__5_/right_grid_pin_0_ sb_8__4_/top_right_grid_pin_1_
+ sb_8__5_/bottom_right_grid_pin_1_ cby_8__5_/prog_clk_0_N_out sb_8__4_/prog_clk_0_N_in
+ cby_8__5_/prog_clk_0_W_in cby_8__5_/right_grid_pin_0_ cby_2__1_
Xcbx_8__6_ cbx_8__6_/REGIN_FEEDTHROUGH cbx_8__6_/REGOUT_FEEDTHROUGH cbx_8__6_/SC_IN_BOT
+ cbx_8__6_/SC_IN_TOP cbx_8__6_/SC_OUT_BOT cbx_8__6_/SC_OUT_TOP VGND VPWR cbx_8__6_/bottom_grid_pin_0_
+ cbx_8__6_/bottom_grid_pin_10_ cbx_8__6_/bottom_grid_pin_11_ cbx_8__6_/bottom_grid_pin_12_
+ cbx_8__6_/bottom_grid_pin_13_ cbx_8__6_/bottom_grid_pin_14_ cbx_8__6_/bottom_grid_pin_15_
+ cbx_8__6_/bottom_grid_pin_1_ cbx_8__6_/bottom_grid_pin_2_ cbx_8__6_/bottom_grid_pin_3_
+ cbx_8__6_/bottom_grid_pin_4_ cbx_8__6_/bottom_grid_pin_5_ cbx_8__6_/bottom_grid_pin_6_
+ cbx_8__6_/bottom_grid_pin_7_ cbx_8__6_/bottom_grid_pin_8_ cbx_8__6_/bottom_grid_pin_9_
+ sb_8__6_/ccff_tail sb_7__6_/ccff_head cbx_8__6_/chanx_left_in[0] cbx_8__6_/chanx_left_in[10]
+ cbx_8__6_/chanx_left_in[11] cbx_8__6_/chanx_left_in[12] cbx_8__6_/chanx_left_in[13]
+ cbx_8__6_/chanx_left_in[14] cbx_8__6_/chanx_left_in[15] cbx_8__6_/chanx_left_in[16]
+ cbx_8__6_/chanx_left_in[17] cbx_8__6_/chanx_left_in[18] cbx_8__6_/chanx_left_in[19]
+ cbx_8__6_/chanx_left_in[1] cbx_8__6_/chanx_left_in[2] cbx_8__6_/chanx_left_in[3]
+ cbx_8__6_/chanx_left_in[4] cbx_8__6_/chanx_left_in[5] cbx_8__6_/chanx_left_in[6]
+ cbx_8__6_/chanx_left_in[7] cbx_8__6_/chanx_left_in[8] cbx_8__6_/chanx_left_in[9]
+ sb_7__6_/chanx_right_in[0] sb_7__6_/chanx_right_in[10] sb_7__6_/chanx_right_in[11]
+ sb_7__6_/chanx_right_in[12] sb_7__6_/chanx_right_in[13] sb_7__6_/chanx_right_in[14]
+ sb_7__6_/chanx_right_in[15] sb_7__6_/chanx_right_in[16] sb_7__6_/chanx_right_in[17]
+ sb_7__6_/chanx_right_in[18] sb_7__6_/chanx_right_in[19] sb_7__6_/chanx_right_in[1]
+ sb_7__6_/chanx_right_in[2] sb_7__6_/chanx_right_in[3] sb_7__6_/chanx_right_in[4]
+ sb_7__6_/chanx_right_in[5] sb_7__6_/chanx_right_in[6] sb_7__6_/chanx_right_in[7]
+ sb_7__6_/chanx_right_in[8] sb_7__6_/chanx_right_in[9] sb_8__6_/chanx_left_out[0]
+ sb_8__6_/chanx_left_out[10] sb_8__6_/chanx_left_out[11] sb_8__6_/chanx_left_out[12]
+ sb_8__6_/chanx_left_out[13] sb_8__6_/chanx_left_out[14] sb_8__6_/chanx_left_out[15]
+ sb_8__6_/chanx_left_out[16] sb_8__6_/chanx_left_out[17] sb_8__6_/chanx_left_out[18]
+ sb_8__6_/chanx_left_out[19] sb_8__6_/chanx_left_out[1] sb_8__6_/chanx_left_out[2]
+ sb_8__6_/chanx_left_out[3] sb_8__6_/chanx_left_out[4] sb_8__6_/chanx_left_out[5]
+ sb_8__6_/chanx_left_out[6] sb_8__6_/chanx_left_out[7] sb_8__6_/chanx_left_out[8]
+ sb_8__6_/chanx_left_out[9] sb_8__6_/chanx_left_in[0] sb_8__6_/chanx_left_in[10]
+ sb_8__6_/chanx_left_in[11] sb_8__6_/chanx_left_in[12] sb_8__6_/chanx_left_in[13]
+ sb_8__6_/chanx_left_in[14] sb_8__6_/chanx_left_in[15] sb_8__6_/chanx_left_in[16]
+ sb_8__6_/chanx_left_in[17] sb_8__6_/chanx_left_in[18] sb_8__6_/chanx_left_in[19]
+ sb_8__6_/chanx_left_in[1] sb_8__6_/chanx_left_in[2] sb_8__6_/chanx_left_in[3] sb_8__6_/chanx_left_in[4]
+ sb_8__6_/chanx_left_in[5] sb_8__6_/chanx_left_in[6] sb_8__6_/chanx_left_in[7] sb_8__6_/chanx_left_in[8]
+ sb_8__6_/chanx_left_in[9] cbx_8__6_/clk_1_N_out cbx_8__6_/clk_1_S_out cbx_8__6_/clk_1_W_in
+ cbx_8__6_/clk_2_E_out cbx_8__6_/clk_2_W_in cbx_8__6_/clk_2_W_out cbx_8__6_/clk_3_E_out
+ cbx_8__6_/clk_3_W_in cbx_8__6_/clk_3_W_out cbx_8__6_/prog_clk_0_N_in cbx_8__6_/prog_clk_0_W_out
+ cbx_8__6_/prog_clk_1_N_out cbx_8__6_/prog_clk_1_S_out cbx_8__6_/prog_clk_1_W_in
+ cbx_8__6_/prog_clk_2_E_out cbx_8__6_/prog_clk_2_W_in cbx_8__6_/prog_clk_2_W_out
+ cbx_8__6_/prog_clk_3_E_out cbx_8__6_/prog_clk_3_W_in cbx_8__6_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_5__2_ cby_5__2_/Test_en_W_in cby_5__2_/Test_en_E_out cby_5__2_/Test_en_N_out
+ cby_5__2_/Test_en_W_in cby_5__2_/Test_en_W_in cby_5__2_/Test_en_W_out VGND VPWR
+ cby_5__2_/ccff_head cby_5__2_/ccff_tail sb_5__1_/chany_top_out[0] sb_5__1_/chany_top_out[10]
+ sb_5__1_/chany_top_out[11] sb_5__1_/chany_top_out[12] sb_5__1_/chany_top_out[13]
+ sb_5__1_/chany_top_out[14] sb_5__1_/chany_top_out[15] sb_5__1_/chany_top_out[16]
+ sb_5__1_/chany_top_out[17] sb_5__1_/chany_top_out[18] sb_5__1_/chany_top_out[19]
+ sb_5__1_/chany_top_out[1] sb_5__1_/chany_top_out[2] sb_5__1_/chany_top_out[3] sb_5__1_/chany_top_out[4]
+ sb_5__1_/chany_top_out[5] sb_5__1_/chany_top_out[6] sb_5__1_/chany_top_out[7] sb_5__1_/chany_top_out[8]
+ sb_5__1_/chany_top_out[9] sb_5__1_/chany_top_in[0] sb_5__1_/chany_top_in[10] sb_5__1_/chany_top_in[11]
+ sb_5__1_/chany_top_in[12] sb_5__1_/chany_top_in[13] sb_5__1_/chany_top_in[14] sb_5__1_/chany_top_in[15]
+ sb_5__1_/chany_top_in[16] sb_5__1_/chany_top_in[17] sb_5__1_/chany_top_in[18] sb_5__1_/chany_top_in[19]
+ sb_5__1_/chany_top_in[1] sb_5__1_/chany_top_in[2] sb_5__1_/chany_top_in[3] sb_5__1_/chany_top_in[4]
+ sb_5__1_/chany_top_in[5] sb_5__1_/chany_top_in[6] sb_5__1_/chany_top_in[7] sb_5__1_/chany_top_in[8]
+ sb_5__1_/chany_top_in[9] cby_5__2_/chany_top_in[0] cby_5__2_/chany_top_in[10] cby_5__2_/chany_top_in[11]
+ cby_5__2_/chany_top_in[12] cby_5__2_/chany_top_in[13] cby_5__2_/chany_top_in[14]
+ cby_5__2_/chany_top_in[15] cby_5__2_/chany_top_in[16] cby_5__2_/chany_top_in[17]
+ cby_5__2_/chany_top_in[18] cby_5__2_/chany_top_in[19] cby_5__2_/chany_top_in[1]
+ cby_5__2_/chany_top_in[2] cby_5__2_/chany_top_in[3] cby_5__2_/chany_top_in[4] cby_5__2_/chany_top_in[5]
+ cby_5__2_/chany_top_in[6] cby_5__2_/chany_top_in[7] cby_5__2_/chany_top_in[8] cby_5__2_/chany_top_in[9]
+ cby_5__2_/chany_top_out[0] cby_5__2_/chany_top_out[10] cby_5__2_/chany_top_out[11]
+ cby_5__2_/chany_top_out[12] cby_5__2_/chany_top_out[13] cby_5__2_/chany_top_out[14]
+ cby_5__2_/chany_top_out[15] cby_5__2_/chany_top_out[16] cby_5__2_/chany_top_out[17]
+ cby_5__2_/chany_top_out[18] cby_5__2_/chany_top_out[19] cby_5__2_/chany_top_out[1]
+ cby_5__2_/chany_top_out[2] cby_5__2_/chany_top_out[3] cby_5__2_/chany_top_out[4]
+ cby_5__2_/chany_top_out[5] cby_5__2_/chany_top_out[6] cby_5__2_/chany_top_out[7]
+ cby_5__2_/chany_top_out[8] cby_5__2_/chany_top_out[9] cby_5__2_/clk_2_N_out sb_5__2_/clk_2_S_out
+ sb_5__1_/clk_1_N_in cby_5__2_/clk_3_N_out cby_5__2_/clk_3_S_in cby_5__2_/clk_3_S_out
+ cby_5__2_/left_grid_pin_16_ cby_5__2_/left_grid_pin_17_ cby_5__2_/left_grid_pin_18_
+ cby_5__2_/left_grid_pin_19_ cby_5__2_/left_grid_pin_20_ cby_5__2_/left_grid_pin_21_
+ cby_5__2_/left_grid_pin_22_ cby_5__2_/left_grid_pin_23_ cby_5__2_/left_grid_pin_24_
+ cby_5__2_/left_grid_pin_25_ cby_5__2_/left_grid_pin_26_ cby_5__2_/left_grid_pin_27_
+ cby_5__2_/left_grid_pin_28_ cby_5__2_/left_grid_pin_29_ cby_5__2_/left_grid_pin_30_
+ cby_5__2_/left_grid_pin_31_ cby_5__2_/prog_clk_0_N_out sb_5__1_/prog_clk_0_N_in
+ cby_5__2_/prog_clk_0_W_in cby_5__2_/prog_clk_2_N_out sb_5__2_/prog_clk_2_S_out sb_5__1_/prog_clk_1_N_in
+ cby_5__2_/prog_clk_3_N_out cby_5__2_/prog_clk_3_S_in cby_5__2_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_7__6_ cbx_7__6_/SC_OUT_BOT cbx_7__5_/SC_IN_TOP grid_clb_7__6_/SC_OUT_TOP
+ cby_6__6_/Test_en_E_out cby_7__6_/Test_en_W_in cby_6__6_/Test_en_E_out grid_clb_7__6_/Test_en_W_out
+ VGND VPWR cbx_7__5_/REGIN_FEEDTHROUGH grid_clb_7__6_/bottom_width_0_height_0__pin_51_
+ cby_6__6_/ccff_tail cby_7__6_/ccff_head cbx_7__5_/clk_1_N_out cbx_7__5_/clk_1_N_out
+ cby_7__6_/prog_clk_0_W_in cbx_7__5_/prog_clk_1_N_out grid_clb_7__6_/prog_clk_0_N_out
+ cbx_7__5_/prog_clk_1_N_out cbx_7__5_/prog_clk_0_N_in grid_clb_7__6_/prog_clk_0_W_out
+ cby_7__6_/left_grid_pin_16_ cby_7__6_/left_grid_pin_17_ cby_7__6_/left_grid_pin_18_
+ cby_7__6_/left_grid_pin_19_ cby_7__6_/left_grid_pin_20_ cby_7__6_/left_grid_pin_21_
+ cby_7__6_/left_grid_pin_22_ cby_7__6_/left_grid_pin_23_ cby_7__6_/left_grid_pin_24_
+ cby_7__6_/left_grid_pin_25_ cby_7__6_/left_grid_pin_26_ cby_7__6_/left_grid_pin_27_
+ cby_7__6_/left_grid_pin_28_ cby_7__6_/left_grid_pin_29_ cby_7__6_/left_grid_pin_30_
+ cby_7__6_/left_grid_pin_31_ sb_7__5_/top_left_grid_pin_42_ sb_7__6_/bottom_left_grid_pin_42_
+ sb_7__5_/top_left_grid_pin_43_ sb_7__6_/bottom_left_grid_pin_43_ sb_7__5_/top_left_grid_pin_44_
+ sb_7__6_/bottom_left_grid_pin_44_ sb_7__5_/top_left_grid_pin_45_ sb_7__6_/bottom_left_grid_pin_45_
+ sb_7__5_/top_left_grid_pin_46_ sb_7__6_/bottom_left_grid_pin_46_ sb_7__5_/top_left_grid_pin_47_
+ sb_7__6_/bottom_left_grid_pin_47_ sb_7__5_/top_left_grid_pin_48_ sb_7__6_/bottom_left_grid_pin_48_
+ sb_7__5_/top_left_grid_pin_49_ sb_7__6_/bottom_left_grid_pin_49_ cbx_7__6_/bottom_grid_pin_0_
+ cbx_7__6_/bottom_grid_pin_10_ cbx_7__6_/bottom_grid_pin_11_ cbx_7__6_/bottom_grid_pin_12_
+ cbx_7__6_/bottom_grid_pin_13_ cbx_7__6_/bottom_grid_pin_14_ cbx_7__6_/bottom_grid_pin_15_
+ cbx_7__6_/bottom_grid_pin_1_ cbx_7__6_/bottom_grid_pin_2_ cbx_7__6_/REGOUT_FEEDTHROUGH
+ grid_clb_7__6_/top_width_0_height_0__pin_33_ sb_7__6_/left_bottom_grid_pin_34_ sb_6__6_/right_bottom_grid_pin_34_
+ sb_7__6_/left_bottom_grid_pin_35_ sb_6__6_/right_bottom_grid_pin_35_ sb_7__6_/left_bottom_grid_pin_36_
+ sb_6__6_/right_bottom_grid_pin_36_ sb_7__6_/left_bottom_grid_pin_37_ sb_6__6_/right_bottom_grid_pin_37_
+ sb_7__6_/left_bottom_grid_pin_38_ sb_6__6_/right_bottom_grid_pin_38_ sb_7__6_/left_bottom_grid_pin_39_
+ sb_6__6_/right_bottom_grid_pin_39_ cbx_7__6_/bottom_grid_pin_3_ sb_7__6_/left_bottom_grid_pin_40_
+ sb_6__6_/right_bottom_grid_pin_40_ sb_7__6_/left_bottom_grid_pin_41_ sb_6__6_/right_bottom_grid_pin_41_
+ cbx_7__6_/bottom_grid_pin_4_ cbx_7__6_/bottom_grid_pin_5_ cbx_7__6_/bottom_grid_pin_6_
+ cbx_7__6_/bottom_grid_pin_7_ cbx_7__6_/bottom_grid_pin_8_ cbx_7__6_/bottom_grid_pin_9_
+ grid_clb
Xcbx_5__3_ cbx_5__3_/REGIN_FEEDTHROUGH cbx_5__3_/REGOUT_FEEDTHROUGH cbx_5__3_/SC_IN_BOT
+ cbx_5__3_/SC_IN_TOP cbx_5__3_/SC_OUT_BOT cbx_5__3_/SC_OUT_TOP VGND VPWR cbx_5__3_/bottom_grid_pin_0_
+ cbx_5__3_/bottom_grid_pin_10_ cbx_5__3_/bottom_grid_pin_11_ cbx_5__3_/bottom_grid_pin_12_
+ cbx_5__3_/bottom_grid_pin_13_ cbx_5__3_/bottom_grid_pin_14_ cbx_5__3_/bottom_grid_pin_15_
+ cbx_5__3_/bottom_grid_pin_1_ cbx_5__3_/bottom_grid_pin_2_ cbx_5__3_/bottom_grid_pin_3_
+ cbx_5__3_/bottom_grid_pin_4_ cbx_5__3_/bottom_grid_pin_5_ cbx_5__3_/bottom_grid_pin_6_
+ cbx_5__3_/bottom_grid_pin_7_ cbx_5__3_/bottom_grid_pin_8_ cbx_5__3_/bottom_grid_pin_9_
+ sb_5__3_/ccff_tail sb_4__3_/ccff_head cbx_5__3_/chanx_left_in[0] cbx_5__3_/chanx_left_in[10]
+ cbx_5__3_/chanx_left_in[11] cbx_5__3_/chanx_left_in[12] cbx_5__3_/chanx_left_in[13]
+ cbx_5__3_/chanx_left_in[14] cbx_5__3_/chanx_left_in[15] cbx_5__3_/chanx_left_in[16]
+ cbx_5__3_/chanx_left_in[17] cbx_5__3_/chanx_left_in[18] cbx_5__3_/chanx_left_in[19]
+ cbx_5__3_/chanx_left_in[1] cbx_5__3_/chanx_left_in[2] cbx_5__3_/chanx_left_in[3]
+ cbx_5__3_/chanx_left_in[4] cbx_5__3_/chanx_left_in[5] cbx_5__3_/chanx_left_in[6]
+ cbx_5__3_/chanx_left_in[7] cbx_5__3_/chanx_left_in[8] cbx_5__3_/chanx_left_in[9]
+ sb_4__3_/chanx_right_in[0] sb_4__3_/chanx_right_in[10] sb_4__3_/chanx_right_in[11]
+ sb_4__3_/chanx_right_in[12] sb_4__3_/chanx_right_in[13] sb_4__3_/chanx_right_in[14]
+ sb_4__3_/chanx_right_in[15] sb_4__3_/chanx_right_in[16] sb_4__3_/chanx_right_in[17]
+ sb_4__3_/chanx_right_in[18] sb_4__3_/chanx_right_in[19] sb_4__3_/chanx_right_in[1]
+ sb_4__3_/chanx_right_in[2] sb_4__3_/chanx_right_in[3] sb_4__3_/chanx_right_in[4]
+ sb_4__3_/chanx_right_in[5] sb_4__3_/chanx_right_in[6] sb_4__3_/chanx_right_in[7]
+ sb_4__3_/chanx_right_in[8] sb_4__3_/chanx_right_in[9] sb_5__3_/chanx_left_out[0]
+ sb_5__3_/chanx_left_out[10] sb_5__3_/chanx_left_out[11] sb_5__3_/chanx_left_out[12]
+ sb_5__3_/chanx_left_out[13] sb_5__3_/chanx_left_out[14] sb_5__3_/chanx_left_out[15]
+ sb_5__3_/chanx_left_out[16] sb_5__3_/chanx_left_out[17] sb_5__3_/chanx_left_out[18]
+ sb_5__3_/chanx_left_out[19] sb_5__3_/chanx_left_out[1] sb_5__3_/chanx_left_out[2]
+ sb_5__3_/chanx_left_out[3] sb_5__3_/chanx_left_out[4] sb_5__3_/chanx_left_out[5]
+ sb_5__3_/chanx_left_out[6] sb_5__3_/chanx_left_out[7] sb_5__3_/chanx_left_out[8]
+ sb_5__3_/chanx_left_out[9] sb_5__3_/chanx_left_in[0] sb_5__3_/chanx_left_in[10]
+ sb_5__3_/chanx_left_in[11] sb_5__3_/chanx_left_in[12] sb_5__3_/chanx_left_in[13]
+ sb_5__3_/chanx_left_in[14] sb_5__3_/chanx_left_in[15] sb_5__3_/chanx_left_in[16]
+ sb_5__3_/chanx_left_in[17] sb_5__3_/chanx_left_in[18] sb_5__3_/chanx_left_in[19]
+ sb_5__3_/chanx_left_in[1] sb_5__3_/chanx_left_in[2] sb_5__3_/chanx_left_in[3] sb_5__3_/chanx_left_in[4]
+ sb_5__3_/chanx_left_in[5] sb_5__3_/chanx_left_in[6] sb_5__3_/chanx_left_in[7] sb_5__3_/chanx_left_in[8]
+ sb_5__3_/chanx_left_in[9] cbx_5__3_/clk_1_N_out cbx_5__3_/clk_1_S_out sb_5__3_/clk_1_W_out
+ cbx_5__3_/clk_2_E_out cbx_5__3_/clk_2_W_in cbx_5__3_/clk_2_W_out cbx_5__3_/clk_3_E_out
+ cbx_5__3_/clk_3_W_in cbx_5__3_/clk_3_W_out cbx_5__3_/prog_clk_0_N_in cbx_5__3_/prog_clk_0_W_out
+ cbx_5__3_/prog_clk_1_N_out cbx_5__3_/prog_clk_1_S_out sb_5__3_/prog_clk_1_W_out
+ cbx_5__3_/prog_clk_2_E_out cbx_5__3_/prog_clk_2_W_in cbx_5__3_/prog_clk_2_W_out
+ cbx_5__3_/prog_clk_3_E_out cbx_5__3_/prog_clk_3_W_in cbx_5__3_/prog_clk_3_W_out
+ cbx_1__1_
Xcbx_2__0_ IO_ISOL_N sb_1__0_/SC_OUT_TOP cbx_2__0_/SC_IN_TOP cbx_2__0_/SC_OUT_BOT
+ cbx_2__0_/SC_OUT_TOP VGND VPWR cbx_2__0_/bottom_grid_pin_0_ cbx_2__0_/bottom_grid_pin_10_
+ cbx_2__0_/bottom_grid_pin_12_ cbx_2__0_/bottom_grid_pin_14_ cbx_2__0_/bottom_grid_pin_16_
+ cbx_2__0_/bottom_grid_pin_2_ cbx_2__0_/bottom_grid_pin_4_ cbx_2__0_/bottom_grid_pin_6_
+ cbx_2__0_/bottom_grid_pin_8_ sb_2__0_/ccff_tail sb_1__0_/ccff_head cbx_2__0_/chanx_left_in[0]
+ cbx_2__0_/chanx_left_in[10] cbx_2__0_/chanx_left_in[11] cbx_2__0_/chanx_left_in[12]
+ cbx_2__0_/chanx_left_in[13] cbx_2__0_/chanx_left_in[14] cbx_2__0_/chanx_left_in[15]
+ cbx_2__0_/chanx_left_in[16] cbx_2__0_/chanx_left_in[17] cbx_2__0_/chanx_left_in[18]
+ cbx_2__0_/chanx_left_in[19] cbx_2__0_/chanx_left_in[1] cbx_2__0_/chanx_left_in[2]
+ cbx_2__0_/chanx_left_in[3] cbx_2__0_/chanx_left_in[4] cbx_2__0_/chanx_left_in[5]
+ cbx_2__0_/chanx_left_in[6] cbx_2__0_/chanx_left_in[7] cbx_2__0_/chanx_left_in[8]
+ cbx_2__0_/chanx_left_in[9] sb_1__0_/chanx_right_in[0] sb_1__0_/chanx_right_in[10]
+ sb_1__0_/chanx_right_in[11] sb_1__0_/chanx_right_in[12] sb_1__0_/chanx_right_in[13]
+ sb_1__0_/chanx_right_in[14] sb_1__0_/chanx_right_in[15] sb_1__0_/chanx_right_in[16]
+ sb_1__0_/chanx_right_in[17] sb_1__0_/chanx_right_in[18] sb_1__0_/chanx_right_in[19]
+ sb_1__0_/chanx_right_in[1] sb_1__0_/chanx_right_in[2] sb_1__0_/chanx_right_in[3]
+ sb_1__0_/chanx_right_in[4] sb_1__0_/chanx_right_in[5] sb_1__0_/chanx_right_in[6]
+ sb_1__0_/chanx_right_in[7] sb_1__0_/chanx_right_in[8] sb_1__0_/chanx_right_in[9]
+ sb_2__0_/chanx_left_out[0] sb_2__0_/chanx_left_out[10] sb_2__0_/chanx_left_out[11]
+ sb_2__0_/chanx_left_out[12] sb_2__0_/chanx_left_out[13] sb_2__0_/chanx_left_out[14]
+ sb_2__0_/chanx_left_out[15] sb_2__0_/chanx_left_out[16] sb_2__0_/chanx_left_out[17]
+ sb_2__0_/chanx_left_out[18] sb_2__0_/chanx_left_out[19] sb_2__0_/chanx_left_out[1]
+ sb_2__0_/chanx_left_out[2] sb_2__0_/chanx_left_out[3] sb_2__0_/chanx_left_out[4]
+ sb_2__0_/chanx_left_out[5] sb_2__0_/chanx_left_out[6] sb_2__0_/chanx_left_out[7]
+ sb_2__0_/chanx_left_out[8] sb_2__0_/chanx_left_out[9] sb_2__0_/chanx_left_in[0]
+ sb_2__0_/chanx_left_in[10] sb_2__0_/chanx_left_in[11] sb_2__0_/chanx_left_in[12]
+ sb_2__0_/chanx_left_in[13] sb_2__0_/chanx_left_in[14] sb_2__0_/chanx_left_in[15]
+ sb_2__0_/chanx_left_in[16] sb_2__0_/chanx_left_in[17] sb_2__0_/chanx_left_in[18]
+ sb_2__0_/chanx_left_in[19] sb_2__0_/chanx_left_in[1] sb_2__0_/chanx_left_in[2] sb_2__0_/chanx_left_in[3]
+ sb_2__0_/chanx_left_in[4] sb_2__0_/chanx_left_in[5] sb_2__0_/chanx_left_in[6] sb_2__0_/chanx_left_in[7]
+ sb_2__0_/chanx_left_in[8] sb_2__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78] cbx_2__0_/prog_clk_0_N_in
+ cbx_2__0_/prog_clk_0_W_out cbx_2__0_/bottom_grid_pin_0_ cbx_2__0_/bottom_grid_pin_10_
+ sb_2__0_/left_bottom_grid_pin_11_ sb_1__0_/right_bottom_grid_pin_11_ cbx_2__0_/bottom_grid_pin_12_
+ sb_2__0_/left_bottom_grid_pin_13_ sb_1__0_/right_bottom_grid_pin_13_ cbx_2__0_/bottom_grid_pin_14_
+ sb_2__0_/left_bottom_grid_pin_15_ sb_1__0_/right_bottom_grid_pin_15_ cbx_2__0_/bottom_grid_pin_16_
+ sb_2__0_/left_bottom_grid_pin_17_ sb_1__0_/right_bottom_grid_pin_17_ sb_2__0_/left_bottom_grid_pin_1_
+ sb_1__0_/right_bottom_grid_pin_1_ cbx_2__0_/bottom_grid_pin_2_ sb_2__0_/left_bottom_grid_pin_3_
+ sb_1__0_/right_bottom_grid_pin_3_ cbx_2__0_/bottom_grid_pin_4_ sb_2__0_/left_bottom_grid_pin_5_
+ sb_1__0_/right_bottom_grid_pin_5_ cbx_2__0_/bottom_grid_pin_6_ sb_2__0_/left_bottom_grid_pin_7_
+ sb_1__0_/right_bottom_grid_pin_7_ cbx_2__0_/bottom_grid_pin_8_ sb_2__0_/left_bottom_grid_pin_9_
+ sb_1__0_/right_bottom_grid_pin_9_ cbx_1__0_
Xgrid_clb_4__3_ cbx_4__2_/SC_OUT_TOP grid_clb_4__3_/SC_OUT_BOT cbx_4__3_/SC_IN_BOT
+ cby_4__3_/Test_en_W_out grid_clb_4__3_/Test_en_E_out cby_4__3_/Test_en_W_out cby_3__3_/Test_en_W_in
+ VGND VPWR cbx_4__2_/REGIN_FEEDTHROUGH grid_clb_4__3_/bottom_width_0_height_0__pin_51_
+ cby_3__3_/ccff_tail cby_4__3_/ccff_head cbx_4__3_/clk_1_S_out cbx_4__3_/clk_1_S_out
+ cby_4__3_/prog_clk_0_W_in cbx_4__3_/prog_clk_1_S_out grid_clb_4__3_/prog_clk_0_N_out
+ cbx_4__3_/prog_clk_1_S_out cbx_4__2_/prog_clk_0_N_in grid_clb_4__3_/prog_clk_0_W_out
+ cby_4__3_/left_grid_pin_16_ cby_4__3_/left_grid_pin_17_ cby_4__3_/left_grid_pin_18_
+ cby_4__3_/left_grid_pin_19_ cby_4__3_/left_grid_pin_20_ cby_4__3_/left_grid_pin_21_
+ cby_4__3_/left_grid_pin_22_ cby_4__3_/left_grid_pin_23_ cby_4__3_/left_grid_pin_24_
+ cby_4__3_/left_grid_pin_25_ cby_4__3_/left_grid_pin_26_ cby_4__3_/left_grid_pin_27_
+ cby_4__3_/left_grid_pin_28_ cby_4__3_/left_grid_pin_29_ cby_4__3_/left_grid_pin_30_
+ cby_4__3_/left_grid_pin_31_ sb_4__2_/top_left_grid_pin_42_ sb_4__3_/bottom_left_grid_pin_42_
+ sb_4__2_/top_left_grid_pin_43_ sb_4__3_/bottom_left_grid_pin_43_ sb_4__2_/top_left_grid_pin_44_
+ sb_4__3_/bottom_left_grid_pin_44_ sb_4__2_/top_left_grid_pin_45_ sb_4__3_/bottom_left_grid_pin_45_
+ sb_4__2_/top_left_grid_pin_46_ sb_4__3_/bottom_left_grid_pin_46_ sb_4__2_/top_left_grid_pin_47_
+ sb_4__3_/bottom_left_grid_pin_47_ sb_4__2_/top_left_grid_pin_48_ sb_4__3_/bottom_left_grid_pin_48_
+ sb_4__2_/top_left_grid_pin_49_ sb_4__3_/bottom_left_grid_pin_49_ cbx_4__3_/bottom_grid_pin_0_
+ cbx_4__3_/bottom_grid_pin_10_ cbx_4__3_/bottom_grid_pin_11_ cbx_4__3_/bottom_grid_pin_12_
+ cbx_4__3_/bottom_grid_pin_13_ cbx_4__3_/bottom_grid_pin_14_ cbx_4__3_/bottom_grid_pin_15_
+ cbx_4__3_/bottom_grid_pin_1_ cbx_4__3_/bottom_grid_pin_2_ cbx_4__3_/REGOUT_FEEDTHROUGH
+ grid_clb_4__3_/top_width_0_height_0__pin_33_ sb_4__3_/left_bottom_grid_pin_34_ sb_3__3_/right_bottom_grid_pin_34_
+ sb_4__3_/left_bottom_grid_pin_35_ sb_3__3_/right_bottom_grid_pin_35_ sb_4__3_/left_bottom_grid_pin_36_
+ sb_3__3_/right_bottom_grid_pin_36_ sb_4__3_/left_bottom_grid_pin_37_ sb_3__3_/right_bottom_grid_pin_37_
+ sb_4__3_/left_bottom_grid_pin_38_ sb_3__3_/right_bottom_grid_pin_38_ sb_4__3_/left_bottom_grid_pin_39_
+ sb_3__3_/right_bottom_grid_pin_39_ cbx_4__3_/bottom_grid_pin_3_ sb_4__3_/left_bottom_grid_pin_40_
+ sb_3__3_/right_bottom_grid_pin_40_ sb_4__3_/left_bottom_grid_pin_41_ sb_3__3_/right_bottom_grid_pin_41_
+ cbx_4__3_/bottom_grid_pin_4_ cbx_4__3_/bottom_grid_pin_5_ cbx_4__3_/bottom_grid_pin_6_
+ cbx_4__3_/bottom_grid_pin_7_ cbx_4__3_/bottom_grid_pin_8_ cbx_4__3_/bottom_grid_pin_9_
+ grid_clb
Xsb_5__8_ sb_5__8_/SC_IN_BOT sb_5__8_/SC_OUT_BOT VGND VPWR sb_5__8_/bottom_left_grid_pin_42_
+ sb_5__8_/bottom_left_grid_pin_43_ sb_5__8_/bottom_left_grid_pin_44_ sb_5__8_/bottom_left_grid_pin_45_
+ sb_5__8_/bottom_left_grid_pin_46_ sb_5__8_/bottom_left_grid_pin_47_ sb_5__8_/bottom_left_grid_pin_48_
+ sb_5__8_/bottom_left_grid_pin_49_ sb_5__8_/ccff_head sb_5__8_/ccff_tail sb_5__8_/chanx_left_in[0]
+ sb_5__8_/chanx_left_in[10] sb_5__8_/chanx_left_in[11] sb_5__8_/chanx_left_in[12]
+ sb_5__8_/chanx_left_in[13] sb_5__8_/chanx_left_in[14] sb_5__8_/chanx_left_in[15]
+ sb_5__8_/chanx_left_in[16] sb_5__8_/chanx_left_in[17] sb_5__8_/chanx_left_in[18]
+ sb_5__8_/chanx_left_in[19] sb_5__8_/chanx_left_in[1] sb_5__8_/chanx_left_in[2] sb_5__8_/chanx_left_in[3]
+ sb_5__8_/chanx_left_in[4] sb_5__8_/chanx_left_in[5] sb_5__8_/chanx_left_in[6] sb_5__8_/chanx_left_in[7]
+ sb_5__8_/chanx_left_in[8] sb_5__8_/chanx_left_in[9] sb_5__8_/chanx_left_out[0] sb_5__8_/chanx_left_out[10]
+ sb_5__8_/chanx_left_out[11] sb_5__8_/chanx_left_out[12] sb_5__8_/chanx_left_out[13]
+ sb_5__8_/chanx_left_out[14] sb_5__8_/chanx_left_out[15] sb_5__8_/chanx_left_out[16]
+ sb_5__8_/chanx_left_out[17] sb_5__8_/chanx_left_out[18] sb_5__8_/chanx_left_out[19]
+ sb_5__8_/chanx_left_out[1] sb_5__8_/chanx_left_out[2] sb_5__8_/chanx_left_out[3]
+ sb_5__8_/chanx_left_out[4] sb_5__8_/chanx_left_out[5] sb_5__8_/chanx_left_out[6]
+ sb_5__8_/chanx_left_out[7] sb_5__8_/chanx_left_out[8] sb_5__8_/chanx_left_out[9]
+ sb_5__8_/chanx_right_in[0] sb_5__8_/chanx_right_in[10] sb_5__8_/chanx_right_in[11]
+ sb_5__8_/chanx_right_in[12] sb_5__8_/chanx_right_in[13] sb_5__8_/chanx_right_in[14]
+ sb_5__8_/chanx_right_in[15] sb_5__8_/chanx_right_in[16] sb_5__8_/chanx_right_in[17]
+ sb_5__8_/chanx_right_in[18] sb_5__8_/chanx_right_in[19] sb_5__8_/chanx_right_in[1]
+ sb_5__8_/chanx_right_in[2] sb_5__8_/chanx_right_in[3] sb_5__8_/chanx_right_in[4]
+ sb_5__8_/chanx_right_in[5] sb_5__8_/chanx_right_in[6] sb_5__8_/chanx_right_in[7]
+ sb_5__8_/chanx_right_in[8] sb_5__8_/chanx_right_in[9] cbx_6__8_/chanx_left_in[0]
+ cbx_6__8_/chanx_left_in[10] cbx_6__8_/chanx_left_in[11] cbx_6__8_/chanx_left_in[12]
+ cbx_6__8_/chanx_left_in[13] cbx_6__8_/chanx_left_in[14] cbx_6__8_/chanx_left_in[15]
+ cbx_6__8_/chanx_left_in[16] cbx_6__8_/chanx_left_in[17] cbx_6__8_/chanx_left_in[18]
+ cbx_6__8_/chanx_left_in[19] cbx_6__8_/chanx_left_in[1] cbx_6__8_/chanx_left_in[2]
+ cbx_6__8_/chanx_left_in[3] cbx_6__8_/chanx_left_in[4] cbx_6__8_/chanx_left_in[5]
+ cbx_6__8_/chanx_left_in[6] cbx_6__8_/chanx_left_in[7] cbx_6__8_/chanx_left_in[8]
+ cbx_6__8_/chanx_left_in[9] cby_5__8_/chany_top_out[0] cby_5__8_/chany_top_out[10]
+ cby_5__8_/chany_top_out[11] cby_5__8_/chany_top_out[12] cby_5__8_/chany_top_out[13]
+ cby_5__8_/chany_top_out[14] cby_5__8_/chany_top_out[15] cby_5__8_/chany_top_out[16]
+ cby_5__8_/chany_top_out[17] cby_5__8_/chany_top_out[18] cby_5__8_/chany_top_out[19]
+ cby_5__8_/chany_top_out[1] cby_5__8_/chany_top_out[2] cby_5__8_/chany_top_out[3]
+ cby_5__8_/chany_top_out[4] cby_5__8_/chany_top_out[5] cby_5__8_/chany_top_out[6]
+ cby_5__8_/chany_top_out[7] cby_5__8_/chany_top_out[8] cby_5__8_/chany_top_out[9]
+ cby_5__8_/chany_top_in[0] cby_5__8_/chany_top_in[10] cby_5__8_/chany_top_in[11]
+ cby_5__8_/chany_top_in[12] cby_5__8_/chany_top_in[13] cby_5__8_/chany_top_in[14]
+ cby_5__8_/chany_top_in[15] cby_5__8_/chany_top_in[16] cby_5__8_/chany_top_in[17]
+ cby_5__8_/chany_top_in[18] cby_5__8_/chany_top_in[19] cby_5__8_/chany_top_in[1]
+ cby_5__8_/chany_top_in[2] cby_5__8_/chany_top_in[3] cby_5__8_/chany_top_in[4] cby_5__8_/chany_top_in[5]
+ cby_5__8_/chany_top_in[6] cby_5__8_/chany_top_in[7] cby_5__8_/chany_top_in[8] cby_5__8_/chany_top_in[9]
+ sb_5__8_/left_bottom_grid_pin_34_ sb_5__8_/left_bottom_grid_pin_35_ sb_5__8_/left_bottom_grid_pin_36_
+ sb_5__8_/left_bottom_grid_pin_37_ sb_5__8_/left_bottom_grid_pin_38_ sb_5__8_/left_bottom_grid_pin_39_
+ sb_5__8_/left_bottom_grid_pin_40_ sb_5__8_/left_bottom_grid_pin_41_ sb_5__8_/left_top_grid_pin_1_
+ sb_5__8_/prog_clk_0_S_in sb_5__8_/right_bottom_grid_pin_34_ sb_5__8_/right_bottom_grid_pin_35_
+ sb_5__8_/right_bottom_grid_pin_36_ sb_5__8_/right_bottom_grid_pin_37_ sb_5__8_/right_bottom_grid_pin_38_
+ sb_5__8_/right_bottom_grid_pin_39_ sb_5__8_/right_bottom_grid_pin_40_ sb_5__8_/right_bottom_grid_pin_41_
+ sb_5__8_/right_top_grid_pin_1_ sb_1__2_
Xsb_2__5_ sb_2__5_/Test_en_N_out sb_2__5_/Test_en_S_in VGND VPWR sb_2__5_/bottom_left_grid_pin_42_
+ sb_2__5_/bottom_left_grid_pin_43_ sb_2__5_/bottom_left_grid_pin_44_ sb_2__5_/bottom_left_grid_pin_45_
+ sb_2__5_/bottom_left_grid_pin_46_ sb_2__5_/bottom_left_grid_pin_47_ sb_2__5_/bottom_left_grid_pin_48_
+ sb_2__5_/bottom_left_grid_pin_49_ sb_2__5_/ccff_head sb_2__5_/ccff_tail sb_2__5_/chanx_left_in[0]
+ sb_2__5_/chanx_left_in[10] sb_2__5_/chanx_left_in[11] sb_2__5_/chanx_left_in[12]
+ sb_2__5_/chanx_left_in[13] sb_2__5_/chanx_left_in[14] sb_2__5_/chanx_left_in[15]
+ sb_2__5_/chanx_left_in[16] sb_2__5_/chanx_left_in[17] sb_2__5_/chanx_left_in[18]
+ sb_2__5_/chanx_left_in[19] sb_2__5_/chanx_left_in[1] sb_2__5_/chanx_left_in[2] sb_2__5_/chanx_left_in[3]
+ sb_2__5_/chanx_left_in[4] sb_2__5_/chanx_left_in[5] sb_2__5_/chanx_left_in[6] sb_2__5_/chanx_left_in[7]
+ sb_2__5_/chanx_left_in[8] sb_2__5_/chanx_left_in[9] sb_2__5_/chanx_left_out[0] sb_2__5_/chanx_left_out[10]
+ sb_2__5_/chanx_left_out[11] sb_2__5_/chanx_left_out[12] sb_2__5_/chanx_left_out[13]
+ sb_2__5_/chanx_left_out[14] sb_2__5_/chanx_left_out[15] sb_2__5_/chanx_left_out[16]
+ sb_2__5_/chanx_left_out[17] sb_2__5_/chanx_left_out[18] sb_2__5_/chanx_left_out[19]
+ sb_2__5_/chanx_left_out[1] sb_2__5_/chanx_left_out[2] sb_2__5_/chanx_left_out[3]
+ sb_2__5_/chanx_left_out[4] sb_2__5_/chanx_left_out[5] sb_2__5_/chanx_left_out[6]
+ sb_2__5_/chanx_left_out[7] sb_2__5_/chanx_left_out[8] sb_2__5_/chanx_left_out[9]
+ sb_2__5_/chanx_right_in[0] sb_2__5_/chanx_right_in[10] sb_2__5_/chanx_right_in[11]
+ sb_2__5_/chanx_right_in[12] sb_2__5_/chanx_right_in[13] sb_2__5_/chanx_right_in[14]
+ sb_2__5_/chanx_right_in[15] sb_2__5_/chanx_right_in[16] sb_2__5_/chanx_right_in[17]
+ sb_2__5_/chanx_right_in[18] sb_2__5_/chanx_right_in[19] sb_2__5_/chanx_right_in[1]
+ sb_2__5_/chanx_right_in[2] sb_2__5_/chanx_right_in[3] sb_2__5_/chanx_right_in[4]
+ sb_2__5_/chanx_right_in[5] sb_2__5_/chanx_right_in[6] sb_2__5_/chanx_right_in[7]
+ sb_2__5_/chanx_right_in[8] sb_2__5_/chanx_right_in[9] cbx_3__5_/chanx_left_in[0]
+ cbx_3__5_/chanx_left_in[10] cbx_3__5_/chanx_left_in[11] cbx_3__5_/chanx_left_in[12]
+ cbx_3__5_/chanx_left_in[13] cbx_3__5_/chanx_left_in[14] cbx_3__5_/chanx_left_in[15]
+ cbx_3__5_/chanx_left_in[16] cbx_3__5_/chanx_left_in[17] cbx_3__5_/chanx_left_in[18]
+ cbx_3__5_/chanx_left_in[19] cbx_3__5_/chanx_left_in[1] cbx_3__5_/chanx_left_in[2]
+ cbx_3__5_/chanx_left_in[3] cbx_3__5_/chanx_left_in[4] cbx_3__5_/chanx_left_in[5]
+ cbx_3__5_/chanx_left_in[6] cbx_3__5_/chanx_left_in[7] cbx_3__5_/chanx_left_in[8]
+ cbx_3__5_/chanx_left_in[9] cby_2__5_/chany_top_out[0] cby_2__5_/chany_top_out[10]
+ cby_2__5_/chany_top_out[11] cby_2__5_/chany_top_out[12] cby_2__5_/chany_top_out[13]
+ cby_2__5_/chany_top_out[14] cby_2__5_/chany_top_out[15] cby_2__5_/chany_top_out[16]
+ cby_2__5_/chany_top_out[17] cby_2__5_/chany_top_out[18] cby_2__5_/chany_top_out[19]
+ cby_2__5_/chany_top_out[1] cby_2__5_/chany_top_out[2] cby_2__5_/chany_top_out[3]
+ cby_2__5_/chany_top_out[4] cby_2__5_/chany_top_out[5] cby_2__5_/chany_top_out[6]
+ cby_2__5_/chany_top_out[7] cby_2__5_/chany_top_out[8] cby_2__5_/chany_top_out[9]
+ cby_2__5_/chany_top_in[0] cby_2__5_/chany_top_in[10] cby_2__5_/chany_top_in[11]
+ cby_2__5_/chany_top_in[12] cby_2__5_/chany_top_in[13] cby_2__5_/chany_top_in[14]
+ cby_2__5_/chany_top_in[15] cby_2__5_/chany_top_in[16] cby_2__5_/chany_top_in[17]
+ cby_2__5_/chany_top_in[18] cby_2__5_/chany_top_in[19] cby_2__5_/chany_top_in[1]
+ cby_2__5_/chany_top_in[2] cby_2__5_/chany_top_in[3] cby_2__5_/chany_top_in[4] cby_2__5_/chany_top_in[5]
+ cby_2__5_/chany_top_in[6] cby_2__5_/chany_top_in[7] cby_2__5_/chany_top_in[8] cby_2__5_/chany_top_in[9]
+ sb_2__5_/chany_top_in[0] sb_2__5_/chany_top_in[10] sb_2__5_/chany_top_in[11] sb_2__5_/chany_top_in[12]
+ sb_2__5_/chany_top_in[13] sb_2__5_/chany_top_in[14] sb_2__5_/chany_top_in[15] sb_2__5_/chany_top_in[16]
+ sb_2__5_/chany_top_in[17] sb_2__5_/chany_top_in[18] sb_2__5_/chany_top_in[19] sb_2__5_/chany_top_in[1]
+ sb_2__5_/chany_top_in[2] sb_2__5_/chany_top_in[3] sb_2__5_/chany_top_in[4] sb_2__5_/chany_top_in[5]
+ sb_2__5_/chany_top_in[6] sb_2__5_/chany_top_in[7] sb_2__5_/chany_top_in[8] sb_2__5_/chany_top_in[9]
+ sb_2__5_/chany_top_out[0] sb_2__5_/chany_top_out[10] sb_2__5_/chany_top_out[11]
+ sb_2__5_/chany_top_out[12] sb_2__5_/chany_top_out[13] sb_2__5_/chany_top_out[14]
+ sb_2__5_/chany_top_out[15] sb_2__5_/chany_top_out[16] sb_2__5_/chany_top_out[17]
+ sb_2__5_/chany_top_out[18] sb_2__5_/chany_top_out[19] sb_2__5_/chany_top_out[1]
+ sb_2__5_/chany_top_out[2] sb_2__5_/chany_top_out[3] sb_2__5_/chany_top_out[4] sb_2__5_/chany_top_out[5]
+ sb_2__5_/chany_top_out[6] sb_2__5_/chany_top_out[7] sb_2__5_/chany_top_out[8] sb_2__5_/chany_top_out[9]
+ sb_2__5_/clk_1_E_out sb_2__5_/clk_1_N_in sb_2__5_/clk_1_W_out sb_2__5_/clk_2_E_out
+ sb_2__5_/clk_2_N_in sb_2__5_/clk_2_N_out sb_2__5_/clk_2_S_out sb_2__5_/clk_2_W_out
+ sb_2__5_/clk_3_E_out sb_2__5_/clk_3_N_in sb_2__5_/clk_3_N_out sb_2__5_/clk_3_S_out
+ sb_2__5_/clk_3_W_out sb_2__5_/left_bottom_grid_pin_34_ sb_2__5_/left_bottom_grid_pin_35_
+ sb_2__5_/left_bottom_grid_pin_36_ sb_2__5_/left_bottom_grid_pin_37_ sb_2__5_/left_bottom_grid_pin_38_
+ sb_2__5_/left_bottom_grid_pin_39_ sb_2__5_/left_bottom_grid_pin_40_ sb_2__5_/left_bottom_grid_pin_41_
+ sb_2__5_/prog_clk_0_N_in sb_2__5_/prog_clk_1_E_out sb_2__5_/prog_clk_1_N_in sb_2__5_/prog_clk_1_W_out
+ sb_2__5_/prog_clk_2_E_out sb_2__5_/prog_clk_2_N_in sb_2__5_/prog_clk_2_N_out sb_2__5_/prog_clk_2_S_out
+ sb_2__5_/prog_clk_2_W_out sb_2__5_/prog_clk_3_E_out sb_2__5_/prog_clk_3_N_in sb_2__5_/prog_clk_3_N_out
+ sb_2__5_/prog_clk_3_S_out sb_2__5_/prog_clk_3_W_out sb_2__5_/right_bottom_grid_pin_34_
+ sb_2__5_/right_bottom_grid_pin_35_ sb_2__5_/right_bottom_grid_pin_36_ sb_2__5_/right_bottom_grid_pin_37_
+ sb_2__5_/right_bottom_grid_pin_38_ sb_2__5_/right_bottom_grid_pin_39_ sb_2__5_/right_bottom_grid_pin_40_
+ sb_2__5_/right_bottom_grid_pin_41_ sb_2__5_/top_left_grid_pin_42_ sb_2__5_/top_left_grid_pin_43_
+ sb_2__5_/top_left_grid_pin_44_ sb_2__5_/top_left_grid_pin_45_ sb_2__5_/top_left_grid_pin_46_
+ sb_2__5_/top_left_grid_pin_47_ sb_2__5_/top_left_grid_pin_48_ sb_2__5_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_8__4_ IO_ISOL_N VGND VPWR cby_8__4_/ccff_head sb_8__3_/ccff_head sb_8__3_/chany_top_out[0]
+ sb_8__3_/chany_top_out[10] sb_8__3_/chany_top_out[11] sb_8__3_/chany_top_out[12]
+ sb_8__3_/chany_top_out[13] sb_8__3_/chany_top_out[14] sb_8__3_/chany_top_out[15]
+ sb_8__3_/chany_top_out[16] sb_8__3_/chany_top_out[17] sb_8__3_/chany_top_out[18]
+ sb_8__3_/chany_top_out[19] sb_8__3_/chany_top_out[1] sb_8__3_/chany_top_out[2] sb_8__3_/chany_top_out[3]
+ sb_8__3_/chany_top_out[4] sb_8__3_/chany_top_out[5] sb_8__3_/chany_top_out[6] sb_8__3_/chany_top_out[7]
+ sb_8__3_/chany_top_out[8] sb_8__3_/chany_top_out[9] sb_8__3_/chany_top_in[0] sb_8__3_/chany_top_in[10]
+ sb_8__3_/chany_top_in[11] sb_8__3_/chany_top_in[12] sb_8__3_/chany_top_in[13] sb_8__3_/chany_top_in[14]
+ sb_8__3_/chany_top_in[15] sb_8__3_/chany_top_in[16] sb_8__3_/chany_top_in[17] sb_8__3_/chany_top_in[18]
+ sb_8__3_/chany_top_in[19] sb_8__3_/chany_top_in[1] sb_8__3_/chany_top_in[2] sb_8__3_/chany_top_in[3]
+ sb_8__3_/chany_top_in[4] sb_8__3_/chany_top_in[5] sb_8__3_/chany_top_in[6] sb_8__3_/chany_top_in[7]
+ sb_8__3_/chany_top_in[8] sb_8__3_/chany_top_in[9] cby_8__4_/chany_top_in[0] cby_8__4_/chany_top_in[10]
+ cby_8__4_/chany_top_in[11] cby_8__4_/chany_top_in[12] cby_8__4_/chany_top_in[13]
+ cby_8__4_/chany_top_in[14] cby_8__4_/chany_top_in[15] cby_8__4_/chany_top_in[16]
+ cby_8__4_/chany_top_in[17] cby_8__4_/chany_top_in[18] cby_8__4_/chany_top_in[19]
+ cby_8__4_/chany_top_in[1] cby_8__4_/chany_top_in[2] cby_8__4_/chany_top_in[3] cby_8__4_/chany_top_in[4]
+ cby_8__4_/chany_top_in[5] cby_8__4_/chany_top_in[6] cby_8__4_/chany_top_in[7] cby_8__4_/chany_top_in[8]
+ cby_8__4_/chany_top_in[9] cby_8__4_/chany_top_out[0] cby_8__4_/chany_top_out[10]
+ cby_8__4_/chany_top_out[11] cby_8__4_/chany_top_out[12] cby_8__4_/chany_top_out[13]
+ cby_8__4_/chany_top_out[14] cby_8__4_/chany_top_out[15] cby_8__4_/chany_top_out[16]
+ cby_8__4_/chany_top_out[17] cby_8__4_/chany_top_out[18] cby_8__4_/chany_top_out[19]
+ cby_8__4_/chany_top_out[1] cby_8__4_/chany_top_out[2] cby_8__4_/chany_top_out[3]
+ cby_8__4_/chany_top_out[4] cby_8__4_/chany_top_out[5] cby_8__4_/chany_top_out[6]
+ cby_8__4_/chany_top_out[7] cby_8__4_/chany_top_out[8] cby_8__4_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
+ cby_8__4_/left_grid_pin_16_ cby_8__4_/left_grid_pin_17_ cby_8__4_/left_grid_pin_18_
+ cby_8__4_/left_grid_pin_19_ cby_8__4_/left_grid_pin_20_ cby_8__4_/left_grid_pin_21_
+ cby_8__4_/left_grid_pin_22_ cby_8__4_/left_grid_pin_23_ cby_8__4_/left_grid_pin_24_
+ cby_8__4_/left_grid_pin_25_ cby_8__4_/left_grid_pin_26_ cby_8__4_/left_grid_pin_27_
+ cby_8__4_/left_grid_pin_28_ cby_8__4_/left_grid_pin_29_ cby_8__4_/left_grid_pin_30_
+ cby_8__4_/left_grid_pin_31_ cby_8__4_/right_grid_pin_0_ sb_8__3_/top_right_grid_pin_1_
+ sb_8__4_/bottom_right_grid_pin_1_ cby_8__4_/prog_clk_0_N_out sb_8__3_/prog_clk_0_N_in
+ cby_8__4_/prog_clk_0_W_in cby_8__4_/right_grid_pin_0_ cby_2__1_
Xcby_5__1_ cby_5__1_/Test_en_W_in cby_5__1_/Test_en_E_out cby_5__1_/Test_en_N_out
+ cby_5__1_/Test_en_W_in cby_5__1_/Test_en_W_in cby_5__1_/Test_en_W_out VGND VPWR
+ cby_5__1_/ccff_head cby_5__1_/ccff_tail sb_5__0_/chany_top_out[0] sb_5__0_/chany_top_out[10]
+ sb_5__0_/chany_top_out[11] sb_5__0_/chany_top_out[12] sb_5__0_/chany_top_out[13]
+ sb_5__0_/chany_top_out[14] sb_5__0_/chany_top_out[15] sb_5__0_/chany_top_out[16]
+ sb_5__0_/chany_top_out[17] sb_5__0_/chany_top_out[18] sb_5__0_/chany_top_out[19]
+ sb_5__0_/chany_top_out[1] sb_5__0_/chany_top_out[2] sb_5__0_/chany_top_out[3] sb_5__0_/chany_top_out[4]
+ sb_5__0_/chany_top_out[5] sb_5__0_/chany_top_out[6] sb_5__0_/chany_top_out[7] sb_5__0_/chany_top_out[8]
+ sb_5__0_/chany_top_out[9] sb_5__0_/chany_top_in[0] sb_5__0_/chany_top_in[10] sb_5__0_/chany_top_in[11]
+ sb_5__0_/chany_top_in[12] sb_5__0_/chany_top_in[13] sb_5__0_/chany_top_in[14] sb_5__0_/chany_top_in[15]
+ sb_5__0_/chany_top_in[16] sb_5__0_/chany_top_in[17] sb_5__0_/chany_top_in[18] sb_5__0_/chany_top_in[19]
+ sb_5__0_/chany_top_in[1] sb_5__0_/chany_top_in[2] sb_5__0_/chany_top_in[3] sb_5__0_/chany_top_in[4]
+ sb_5__0_/chany_top_in[5] sb_5__0_/chany_top_in[6] sb_5__0_/chany_top_in[7] sb_5__0_/chany_top_in[8]
+ sb_5__0_/chany_top_in[9] cby_5__1_/chany_top_in[0] cby_5__1_/chany_top_in[10] cby_5__1_/chany_top_in[11]
+ cby_5__1_/chany_top_in[12] cby_5__1_/chany_top_in[13] cby_5__1_/chany_top_in[14]
+ cby_5__1_/chany_top_in[15] cby_5__1_/chany_top_in[16] cby_5__1_/chany_top_in[17]
+ cby_5__1_/chany_top_in[18] cby_5__1_/chany_top_in[19] cby_5__1_/chany_top_in[1]
+ cby_5__1_/chany_top_in[2] cby_5__1_/chany_top_in[3] cby_5__1_/chany_top_in[4] cby_5__1_/chany_top_in[5]
+ cby_5__1_/chany_top_in[6] cby_5__1_/chany_top_in[7] cby_5__1_/chany_top_in[8] cby_5__1_/chany_top_in[9]
+ cby_5__1_/chany_top_out[0] cby_5__1_/chany_top_out[10] cby_5__1_/chany_top_out[11]
+ cby_5__1_/chany_top_out[12] cby_5__1_/chany_top_out[13] cby_5__1_/chany_top_out[14]
+ cby_5__1_/chany_top_out[15] cby_5__1_/chany_top_out[16] cby_5__1_/chany_top_out[17]
+ cby_5__1_/chany_top_out[18] cby_5__1_/chany_top_out[19] cby_5__1_/chany_top_out[1]
+ cby_5__1_/chany_top_out[2] cby_5__1_/chany_top_out[3] cby_5__1_/chany_top_out[4]
+ cby_5__1_/chany_top_out[5] cby_5__1_/chany_top_out[6] cby_5__1_/chany_top_out[7]
+ cby_5__1_/chany_top_out[8] cby_5__1_/chany_top_out[9] cby_5__1_/clk_2_N_out cby_5__1_/clk_2_S_in
+ cby_5__1_/clk_2_S_out cby_5__1_/clk_3_N_out cby_5__1_/clk_3_S_in cby_5__1_/clk_3_S_out
+ cby_5__1_/left_grid_pin_16_ cby_5__1_/left_grid_pin_17_ cby_5__1_/left_grid_pin_18_
+ cby_5__1_/left_grid_pin_19_ cby_5__1_/left_grid_pin_20_ cby_5__1_/left_grid_pin_21_
+ cby_5__1_/left_grid_pin_22_ cby_5__1_/left_grid_pin_23_ cby_5__1_/left_grid_pin_24_
+ cby_5__1_/left_grid_pin_25_ cby_5__1_/left_grid_pin_26_ cby_5__1_/left_grid_pin_27_
+ cby_5__1_/left_grid_pin_28_ cby_5__1_/left_grid_pin_29_ cby_5__1_/left_grid_pin_30_
+ cby_5__1_/left_grid_pin_31_ cby_5__1_/prog_clk_0_N_out sb_5__0_/prog_clk_0_N_in
+ cby_5__1_/prog_clk_0_W_in cby_5__1_/prog_clk_2_N_out cby_5__1_/prog_clk_2_S_in cby_5__1_/prog_clk_2_S_out
+ cby_5__1_/prog_clk_3_N_out cby_5__1_/prog_clk_3_S_in cby_5__1_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_8__5_ cbx_8__5_/REGIN_FEEDTHROUGH cbx_8__5_/REGOUT_FEEDTHROUGH cbx_8__5_/SC_IN_BOT
+ cbx_8__5_/SC_IN_TOP cbx_8__5_/SC_OUT_BOT cbx_8__5_/SC_OUT_TOP VGND VPWR cbx_8__5_/bottom_grid_pin_0_
+ cbx_8__5_/bottom_grid_pin_10_ cbx_8__5_/bottom_grid_pin_11_ cbx_8__5_/bottom_grid_pin_12_
+ cbx_8__5_/bottom_grid_pin_13_ cbx_8__5_/bottom_grid_pin_14_ cbx_8__5_/bottom_grid_pin_15_
+ cbx_8__5_/bottom_grid_pin_1_ cbx_8__5_/bottom_grid_pin_2_ cbx_8__5_/bottom_grid_pin_3_
+ cbx_8__5_/bottom_grid_pin_4_ cbx_8__5_/bottom_grid_pin_5_ cbx_8__5_/bottom_grid_pin_6_
+ cbx_8__5_/bottom_grid_pin_7_ cbx_8__5_/bottom_grid_pin_8_ cbx_8__5_/bottom_grid_pin_9_
+ sb_8__5_/ccff_tail sb_7__5_/ccff_head cbx_8__5_/chanx_left_in[0] cbx_8__5_/chanx_left_in[10]
+ cbx_8__5_/chanx_left_in[11] cbx_8__5_/chanx_left_in[12] cbx_8__5_/chanx_left_in[13]
+ cbx_8__5_/chanx_left_in[14] cbx_8__5_/chanx_left_in[15] cbx_8__5_/chanx_left_in[16]
+ cbx_8__5_/chanx_left_in[17] cbx_8__5_/chanx_left_in[18] cbx_8__5_/chanx_left_in[19]
+ cbx_8__5_/chanx_left_in[1] cbx_8__5_/chanx_left_in[2] cbx_8__5_/chanx_left_in[3]
+ cbx_8__5_/chanx_left_in[4] cbx_8__5_/chanx_left_in[5] cbx_8__5_/chanx_left_in[6]
+ cbx_8__5_/chanx_left_in[7] cbx_8__5_/chanx_left_in[8] cbx_8__5_/chanx_left_in[9]
+ sb_7__5_/chanx_right_in[0] sb_7__5_/chanx_right_in[10] sb_7__5_/chanx_right_in[11]
+ sb_7__5_/chanx_right_in[12] sb_7__5_/chanx_right_in[13] sb_7__5_/chanx_right_in[14]
+ sb_7__5_/chanx_right_in[15] sb_7__5_/chanx_right_in[16] sb_7__5_/chanx_right_in[17]
+ sb_7__5_/chanx_right_in[18] sb_7__5_/chanx_right_in[19] sb_7__5_/chanx_right_in[1]
+ sb_7__5_/chanx_right_in[2] sb_7__5_/chanx_right_in[3] sb_7__5_/chanx_right_in[4]
+ sb_7__5_/chanx_right_in[5] sb_7__5_/chanx_right_in[6] sb_7__5_/chanx_right_in[7]
+ sb_7__5_/chanx_right_in[8] sb_7__5_/chanx_right_in[9] sb_8__5_/chanx_left_out[0]
+ sb_8__5_/chanx_left_out[10] sb_8__5_/chanx_left_out[11] sb_8__5_/chanx_left_out[12]
+ sb_8__5_/chanx_left_out[13] sb_8__5_/chanx_left_out[14] sb_8__5_/chanx_left_out[15]
+ sb_8__5_/chanx_left_out[16] sb_8__5_/chanx_left_out[17] sb_8__5_/chanx_left_out[18]
+ sb_8__5_/chanx_left_out[19] sb_8__5_/chanx_left_out[1] sb_8__5_/chanx_left_out[2]
+ sb_8__5_/chanx_left_out[3] sb_8__5_/chanx_left_out[4] sb_8__5_/chanx_left_out[5]
+ sb_8__5_/chanx_left_out[6] sb_8__5_/chanx_left_out[7] sb_8__5_/chanx_left_out[8]
+ sb_8__5_/chanx_left_out[9] sb_8__5_/chanx_left_in[0] sb_8__5_/chanx_left_in[10]
+ sb_8__5_/chanx_left_in[11] sb_8__5_/chanx_left_in[12] sb_8__5_/chanx_left_in[13]
+ sb_8__5_/chanx_left_in[14] sb_8__5_/chanx_left_in[15] sb_8__5_/chanx_left_in[16]
+ sb_8__5_/chanx_left_in[17] sb_8__5_/chanx_left_in[18] sb_8__5_/chanx_left_in[19]
+ sb_8__5_/chanx_left_in[1] sb_8__5_/chanx_left_in[2] sb_8__5_/chanx_left_in[3] sb_8__5_/chanx_left_in[4]
+ sb_8__5_/chanx_left_in[5] sb_8__5_/chanx_left_in[6] sb_8__5_/chanx_left_in[7] sb_8__5_/chanx_left_in[8]
+ sb_8__5_/chanx_left_in[9] cbx_8__5_/clk_1_N_out cbx_8__5_/clk_1_S_out sb_7__5_/clk_1_E_out
+ cbx_8__5_/clk_2_E_out cbx_8__5_/clk_2_W_in cbx_8__5_/clk_2_W_out cbx_8__5_/clk_3_E_out
+ cbx_8__5_/clk_3_W_in cbx_8__5_/clk_3_W_out cbx_8__5_/prog_clk_0_N_in cbx_8__5_/prog_clk_0_W_out
+ cbx_8__5_/prog_clk_1_N_out cbx_8__5_/prog_clk_1_S_out sb_7__5_/prog_clk_1_E_out
+ cbx_8__5_/prog_clk_2_E_out cbx_8__5_/prog_clk_2_W_in cbx_8__5_/prog_clk_2_W_out
+ cbx_8__5_/prog_clk_3_E_out cbx_8__5_/prog_clk_3_W_in cbx_8__5_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_7__5_ cbx_7__5_/SC_OUT_BOT cbx_7__4_/SC_IN_TOP grid_clb_7__5_/SC_OUT_TOP
+ cby_6__5_/Test_en_E_out cby_7__5_/Test_en_W_in cby_6__5_/Test_en_E_out grid_clb_7__5_/Test_en_W_out
+ VGND VPWR cbx_7__4_/REGIN_FEEDTHROUGH grid_clb_7__5_/bottom_width_0_height_0__pin_51_
+ cby_6__5_/ccff_tail cby_7__5_/ccff_head cbx_7__5_/clk_1_S_out cbx_7__5_/clk_1_S_out
+ cby_7__5_/prog_clk_0_W_in cbx_7__5_/prog_clk_1_S_out grid_clb_7__5_/prog_clk_0_N_out
+ cbx_7__5_/prog_clk_1_S_out cbx_7__4_/prog_clk_0_N_in grid_clb_7__5_/prog_clk_0_W_out
+ cby_7__5_/left_grid_pin_16_ cby_7__5_/left_grid_pin_17_ cby_7__5_/left_grid_pin_18_
+ cby_7__5_/left_grid_pin_19_ cby_7__5_/left_grid_pin_20_ cby_7__5_/left_grid_pin_21_
+ cby_7__5_/left_grid_pin_22_ cby_7__5_/left_grid_pin_23_ cby_7__5_/left_grid_pin_24_
+ cby_7__5_/left_grid_pin_25_ cby_7__5_/left_grid_pin_26_ cby_7__5_/left_grid_pin_27_
+ cby_7__5_/left_grid_pin_28_ cby_7__5_/left_grid_pin_29_ cby_7__5_/left_grid_pin_30_
+ cby_7__5_/left_grid_pin_31_ sb_7__4_/top_left_grid_pin_42_ sb_7__5_/bottom_left_grid_pin_42_
+ sb_7__4_/top_left_grid_pin_43_ sb_7__5_/bottom_left_grid_pin_43_ sb_7__4_/top_left_grid_pin_44_
+ sb_7__5_/bottom_left_grid_pin_44_ sb_7__4_/top_left_grid_pin_45_ sb_7__5_/bottom_left_grid_pin_45_
+ sb_7__4_/top_left_grid_pin_46_ sb_7__5_/bottom_left_grid_pin_46_ sb_7__4_/top_left_grid_pin_47_
+ sb_7__5_/bottom_left_grid_pin_47_ sb_7__4_/top_left_grid_pin_48_ sb_7__5_/bottom_left_grid_pin_48_
+ sb_7__4_/top_left_grid_pin_49_ sb_7__5_/bottom_left_grid_pin_49_ cbx_7__5_/bottom_grid_pin_0_
+ cbx_7__5_/bottom_grid_pin_10_ cbx_7__5_/bottom_grid_pin_11_ cbx_7__5_/bottom_grid_pin_12_
+ cbx_7__5_/bottom_grid_pin_13_ cbx_7__5_/bottom_grid_pin_14_ cbx_7__5_/bottom_grid_pin_15_
+ cbx_7__5_/bottom_grid_pin_1_ cbx_7__5_/bottom_grid_pin_2_ cbx_7__5_/REGOUT_FEEDTHROUGH
+ grid_clb_7__5_/top_width_0_height_0__pin_33_ sb_7__5_/left_bottom_grid_pin_34_ sb_6__5_/right_bottom_grid_pin_34_
+ sb_7__5_/left_bottom_grid_pin_35_ sb_6__5_/right_bottom_grid_pin_35_ sb_7__5_/left_bottom_grid_pin_36_
+ sb_6__5_/right_bottom_grid_pin_36_ sb_7__5_/left_bottom_grid_pin_37_ sb_6__5_/right_bottom_grid_pin_37_
+ sb_7__5_/left_bottom_grid_pin_38_ sb_6__5_/right_bottom_grid_pin_38_ sb_7__5_/left_bottom_grid_pin_39_
+ sb_6__5_/right_bottom_grid_pin_39_ cbx_7__5_/bottom_grid_pin_3_ sb_7__5_/left_bottom_grid_pin_40_
+ sb_6__5_/right_bottom_grid_pin_40_ sb_7__5_/left_bottom_grid_pin_41_ sb_6__5_/right_bottom_grid_pin_41_
+ cbx_7__5_/bottom_grid_pin_4_ cbx_7__5_/bottom_grid_pin_5_ cbx_7__5_/bottom_grid_pin_6_
+ cbx_7__5_/bottom_grid_pin_7_ cbx_7__5_/bottom_grid_pin_8_ cbx_7__5_/bottom_grid_pin_9_
+ grid_clb
Xcbx_5__2_ cbx_5__2_/REGIN_FEEDTHROUGH cbx_5__2_/REGOUT_FEEDTHROUGH cbx_5__2_/SC_IN_BOT
+ cbx_5__2_/SC_IN_TOP cbx_5__2_/SC_OUT_BOT cbx_5__2_/SC_OUT_TOP VGND VPWR cbx_5__2_/bottom_grid_pin_0_
+ cbx_5__2_/bottom_grid_pin_10_ cbx_5__2_/bottom_grid_pin_11_ cbx_5__2_/bottom_grid_pin_12_
+ cbx_5__2_/bottom_grid_pin_13_ cbx_5__2_/bottom_grid_pin_14_ cbx_5__2_/bottom_grid_pin_15_
+ cbx_5__2_/bottom_grid_pin_1_ cbx_5__2_/bottom_grid_pin_2_ cbx_5__2_/bottom_grid_pin_3_
+ cbx_5__2_/bottom_grid_pin_4_ cbx_5__2_/bottom_grid_pin_5_ cbx_5__2_/bottom_grid_pin_6_
+ cbx_5__2_/bottom_grid_pin_7_ cbx_5__2_/bottom_grid_pin_8_ cbx_5__2_/bottom_grid_pin_9_
+ sb_5__2_/ccff_tail sb_4__2_/ccff_head cbx_5__2_/chanx_left_in[0] cbx_5__2_/chanx_left_in[10]
+ cbx_5__2_/chanx_left_in[11] cbx_5__2_/chanx_left_in[12] cbx_5__2_/chanx_left_in[13]
+ cbx_5__2_/chanx_left_in[14] cbx_5__2_/chanx_left_in[15] cbx_5__2_/chanx_left_in[16]
+ cbx_5__2_/chanx_left_in[17] cbx_5__2_/chanx_left_in[18] cbx_5__2_/chanx_left_in[19]
+ cbx_5__2_/chanx_left_in[1] cbx_5__2_/chanx_left_in[2] cbx_5__2_/chanx_left_in[3]
+ cbx_5__2_/chanx_left_in[4] cbx_5__2_/chanx_left_in[5] cbx_5__2_/chanx_left_in[6]
+ cbx_5__2_/chanx_left_in[7] cbx_5__2_/chanx_left_in[8] cbx_5__2_/chanx_left_in[9]
+ sb_4__2_/chanx_right_in[0] sb_4__2_/chanx_right_in[10] sb_4__2_/chanx_right_in[11]
+ sb_4__2_/chanx_right_in[12] sb_4__2_/chanx_right_in[13] sb_4__2_/chanx_right_in[14]
+ sb_4__2_/chanx_right_in[15] sb_4__2_/chanx_right_in[16] sb_4__2_/chanx_right_in[17]
+ sb_4__2_/chanx_right_in[18] sb_4__2_/chanx_right_in[19] sb_4__2_/chanx_right_in[1]
+ sb_4__2_/chanx_right_in[2] sb_4__2_/chanx_right_in[3] sb_4__2_/chanx_right_in[4]
+ sb_4__2_/chanx_right_in[5] sb_4__2_/chanx_right_in[6] sb_4__2_/chanx_right_in[7]
+ sb_4__2_/chanx_right_in[8] sb_4__2_/chanx_right_in[9] sb_5__2_/chanx_left_out[0]
+ sb_5__2_/chanx_left_out[10] sb_5__2_/chanx_left_out[11] sb_5__2_/chanx_left_out[12]
+ sb_5__2_/chanx_left_out[13] sb_5__2_/chanx_left_out[14] sb_5__2_/chanx_left_out[15]
+ sb_5__2_/chanx_left_out[16] sb_5__2_/chanx_left_out[17] sb_5__2_/chanx_left_out[18]
+ sb_5__2_/chanx_left_out[19] sb_5__2_/chanx_left_out[1] sb_5__2_/chanx_left_out[2]
+ sb_5__2_/chanx_left_out[3] sb_5__2_/chanx_left_out[4] sb_5__2_/chanx_left_out[5]
+ sb_5__2_/chanx_left_out[6] sb_5__2_/chanx_left_out[7] sb_5__2_/chanx_left_out[8]
+ sb_5__2_/chanx_left_out[9] sb_5__2_/chanx_left_in[0] sb_5__2_/chanx_left_in[10]
+ sb_5__2_/chanx_left_in[11] sb_5__2_/chanx_left_in[12] sb_5__2_/chanx_left_in[13]
+ sb_5__2_/chanx_left_in[14] sb_5__2_/chanx_left_in[15] sb_5__2_/chanx_left_in[16]
+ sb_5__2_/chanx_left_in[17] sb_5__2_/chanx_left_in[18] sb_5__2_/chanx_left_in[19]
+ sb_5__2_/chanx_left_in[1] sb_5__2_/chanx_left_in[2] sb_5__2_/chanx_left_in[3] sb_5__2_/chanx_left_in[4]
+ sb_5__2_/chanx_left_in[5] sb_5__2_/chanx_left_in[6] sb_5__2_/chanx_left_in[7] sb_5__2_/chanx_left_in[8]
+ sb_5__2_/chanx_left_in[9] cbx_5__2_/clk_1_N_out cbx_5__2_/clk_1_S_out cbx_5__2_/clk_1_W_in
+ cbx_5__2_/clk_2_E_out cbx_5__2_/clk_2_W_in cbx_5__2_/clk_2_W_out cbx_5__2_/clk_3_E_out
+ cbx_5__2_/clk_3_W_in cbx_5__2_/clk_3_W_out cbx_5__2_/prog_clk_0_N_in cbx_5__2_/prog_clk_0_W_out
+ cbx_5__2_/prog_clk_1_N_out cbx_5__2_/prog_clk_1_S_out cbx_5__2_/prog_clk_1_W_in
+ cbx_5__2_/prog_clk_2_E_out cbx_5__2_/prog_clk_2_W_in cbx_5__2_/prog_clk_2_W_out
+ cbx_5__2_/prog_clk_3_E_out cbx_5__2_/prog_clk_3_W_in cbx_5__2_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_5__7_ sb_5__7_/Test_en_N_out sb_5__7_/Test_en_S_in VGND VPWR sb_5__7_/bottom_left_grid_pin_42_
+ sb_5__7_/bottom_left_grid_pin_43_ sb_5__7_/bottom_left_grid_pin_44_ sb_5__7_/bottom_left_grid_pin_45_
+ sb_5__7_/bottom_left_grid_pin_46_ sb_5__7_/bottom_left_grid_pin_47_ sb_5__7_/bottom_left_grid_pin_48_
+ sb_5__7_/bottom_left_grid_pin_49_ sb_5__7_/ccff_head sb_5__7_/ccff_tail sb_5__7_/chanx_left_in[0]
+ sb_5__7_/chanx_left_in[10] sb_5__7_/chanx_left_in[11] sb_5__7_/chanx_left_in[12]
+ sb_5__7_/chanx_left_in[13] sb_5__7_/chanx_left_in[14] sb_5__7_/chanx_left_in[15]
+ sb_5__7_/chanx_left_in[16] sb_5__7_/chanx_left_in[17] sb_5__7_/chanx_left_in[18]
+ sb_5__7_/chanx_left_in[19] sb_5__7_/chanx_left_in[1] sb_5__7_/chanx_left_in[2] sb_5__7_/chanx_left_in[3]
+ sb_5__7_/chanx_left_in[4] sb_5__7_/chanx_left_in[5] sb_5__7_/chanx_left_in[6] sb_5__7_/chanx_left_in[7]
+ sb_5__7_/chanx_left_in[8] sb_5__7_/chanx_left_in[9] sb_5__7_/chanx_left_out[0] sb_5__7_/chanx_left_out[10]
+ sb_5__7_/chanx_left_out[11] sb_5__7_/chanx_left_out[12] sb_5__7_/chanx_left_out[13]
+ sb_5__7_/chanx_left_out[14] sb_5__7_/chanx_left_out[15] sb_5__7_/chanx_left_out[16]
+ sb_5__7_/chanx_left_out[17] sb_5__7_/chanx_left_out[18] sb_5__7_/chanx_left_out[19]
+ sb_5__7_/chanx_left_out[1] sb_5__7_/chanx_left_out[2] sb_5__7_/chanx_left_out[3]
+ sb_5__7_/chanx_left_out[4] sb_5__7_/chanx_left_out[5] sb_5__7_/chanx_left_out[6]
+ sb_5__7_/chanx_left_out[7] sb_5__7_/chanx_left_out[8] sb_5__7_/chanx_left_out[9]
+ sb_5__7_/chanx_right_in[0] sb_5__7_/chanx_right_in[10] sb_5__7_/chanx_right_in[11]
+ sb_5__7_/chanx_right_in[12] sb_5__7_/chanx_right_in[13] sb_5__7_/chanx_right_in[14]
+ sb_5__7_/chanx_right_in[15] sb_5__7_/chanx_right_in[16] sb_5__7_/chanx_right_in[17]
+ sb_5__7_/chanx_right_in[18] sb_5__7_/chanx_right_in[19] sb_5__7_/chanx_right_in[1]
+ sb_5__7_/chanx_right_in[2] sb_5__7_/chanx_right_in[3] sb_5__7_/chanx_right_in[4]
+ sb_5__7_/chanx_right_in[5] sb_5__7_/chanx_right_in[6] sb_5__7_/chanx_right_in[7]
+ sb_5__7_/chanx_right_in[8] sb_5__7_/chanx_right_in[9] cbx_6__7_/chanx_left_in[0]
+ cbx_6__7_/chanx_left_in[10] cbx_6__7_/chanx_left_in[11] cbx_6__7_/chanx_left_in[12]
+ cbx_6__7_/chanx_left_in[13] cbx_6__7_/chanx_left_in[14] cbx_6__7_/chanx_left_in[15]
+ cbx_6__7_/chanx_left_in[16] cbx_6__7_/chanx_left_in[17] cbx_6__7_/chanx_left_in[18]
+ cbx_6__7_/chanx_left_in[19] cbx_6__7_/chanx_left_in[1] cbx_6__7_/chanx_left_in[2]
+ cbx_6__7_/chanx_left_in[3] cbx_6__7_/chanx_left_in[4] cbx_6__7_/chanx_left_in[5]
+ cbx_6__7_/chanx_left_in[6] cbx_6__7_/chanx_left_in[7] cbx_6__7_/chanx_left_in[8]
+ cbx_6__7_/chanx_left_in[9] cby_5__7_/chany_top_out[0] cby_5__7_/chany_top_out[10]
+ cby_5__7_/chany_top_out[11] cby_5__7_/chany_top_out[12] cby_5__7_/chany_top_out[13]
+ cby_5__7_/chany_top_out[14] cby_5__7_/chany_top_out[15] cby_5__7_/chany_top_out[16]
+ cby_5__7_/chany_top_out[17] cby_5__7_/chany_top_out[18] cby_5__7_/chany_top_out[19]
+ cby_5__7_/chany_top_out[1] cby_5__7_/chany_top_out[2] cby_5__7_/chany_top_out[3]
+ cby_5__7_/chany_top_out[4] cby_5__7_/chany_top_out[5] cby_5__7_/chany_top_out[6]
+ cby_5__7_/chany_top_out[7] cby_5__7_/chany_top_out[8] cby_5__7_/chany_top_out[9]
+ cby_5__7_/chany_top_in[0] cby_5__7_/chany_top_in[10] cby_5__7_/chany_top_in[11]
+ cby_5__7_/chany_top_in[12] cby_5__7_/chany_top_in[13] cby_5__7_/chany_top_in[14]
+ cby_5__7_/chany_top_in[15] cby_5__7_/chany_top_in[16] cby_5__7_/chany_top_in[17]
+ cby_5__7_/chany_top_in[18] cby_5__7_/chany_top_in[19] cby_5__7_/chany_top_in[1]
+ cby_5__7_/chany_top_in[2] cby_5__7_/chany_top_in[3] cby_5__7_/chany_top_in[4] cby_5__7_/chany_top_in[5]
+ cby_5__7_/chany_top_in[6] cby_5__7_/chany_top_in[7] cby_5__7_/chany_top_in[8] cby_5__7_/chany_top_in[9]
+ sb_5__7_/chany_top_in[0] sb_5__7_/chany_top_in[10] sb_5__7_/chany_top_in[11] sb_5__7_/chany_top_in[12]
+ sb_5__7_/chany_top_in[13] sb_5__7_/chany_top_in[14] sb_5__7_/chany_top_in[15] sb_5__7_/chany_top_in[16]
+ sb_5__7_/chany_top_in[17] sb_5__7_/chany_top_in[18] sb_5__7_/chany_top_in[19] sb_5__7_/chany_top_in[1]
+ sb_5__7_/chany_top_in[2] sb_5__7_/chany_top_in[3] sb_5__7_/chany_top_in[4] sb_5__7_/chany_top_in[5]
+ sb_5__7_/chany_top_in[6] sb_5__7_/chany_top_in[7] sb_5__7_/chany_top_in[8] sb_5__7_/chany_top_in[9]
+ sb_5__7_/chany_top_out[0] sb_5__7_/chany_top_out[10] sb_5__7_/chany_top_out[11]
+ sb_5__7_/chany_top_out[12] sb_5__7_/chany_top_out[13] sb_5__7_/chany_top_out[14]
+ sb_5__7_/chany_top_out[15] sb_5__7_/chany_top_out[16] sb_5__7_/chany_top_out[17]
+ sb_5__7_/chany_top_out[18] sb_5__7_/chany_top_out[19] sb_5__7_/chany_top_out[1]
+ sb_5__7_/chany_top_out[2] sb_5__7_/chany_top_out[3] sb_5__7_/chany_top_out[4] sb_5__7_/chany_top_out[5]
+ sb_5__7_/chany_top_out[6] sb_5__7_/chany_top_out[7] sb_5__7_/chany_top_out[8] sb_5__7_/chany_top_out[9]
+ sb_5__7_/clk_1_E_out sb_5__7_/clk_1_N_in sb_5__7_/clk_1_W_out sb_5__7_/clk_2_E_out
+ sb_5__7_/clk_2_N_in sb_5__7_/clk_2_N_out sb_5__7_/clk_2_S_out sb_5__7_/clk_2_W_out
+ sb_5__7_/clk_3_E_out sb_5__7_/clk_3_N_in sb_5__7_/clk_3_N_out sb_5__7_/clk_3_S_out
+ sb_5__7_/clk_3_W_out sb_5__7_/left_bottom_grid_pin_34_ sb_5__7_/left_bottom_grid_pin_35_
+ sb_5__7_/left_bottom_grid_pin_36_ sb_5__7_/left_bottom_grid_pin_37_ sb_5__7_/left_bottom_grid_pin_38_
+ sb_5__7_/left_bottom_grid_pin_39_ sb_5__7_/left_bottom_grid_pin_40_ sb_5__7_/left_bottom_grid_pin_41_
+ sb_5__7_/prog_clk_0_N_in sb_5__7_/prog_clk_1_E_out sb_5__7_/prog_clk_1_N_in sb_5__7_/prog_clk_1_W_out
+ sb_5__7_/prog_clk_2_E_out sb_5__7_/prog_clk_2_N_in sb_5__7_/prog_clk_2_N_out sb_5__7_/prog_clk_2_S_out
+ sb_5__7_/prog_clk_2_W_out sb_5__7_/prog_clk_3_E_out sb_5__7_/prog_clk_3_N_in sb_5__7_/prog_clk_3_N_out
+ sb_5__7_/prog_clk_3_S_out sb_5__7_/prog_clk_3_W_out sb_5__7_/right_bottom_grid_pin_34_
+ sb_5__7_/right_bottom_grid_pin_35_ sb_5__7_/right_bottom_grid_pin_36_ sb_5__7_/right_bottom_grid_pin_37_
+ sb_5__7_/right_bottom_grid_pin_38_ sb_5__7_/right_bottom_grid_pin_39_ sb_5__7_/right_bottom_grid_pin_40_
+ sb_5__7_/right_bottom_grid_pin_41_ sb_5__7_/top_left_grid_pin_42_ sb_5__7_/top_left_grid_pin_43_
+ sb_5__7_/top_left_grid_pin_44_ sb_5__7_/top_left_grid_pin_45_ sb_5__7_/top_left_grid_pin_46_
+ sb_5__7_/top_left_grid_pin_47_ sb_5__7_/top_left_grid_pin_48_ sb_5__7_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_4__2_ cbx_4__1_/SC_OUT_TOP grid_clb_4__2_/SC_OUT_BOT cbx_4__2_/SC_IN_BOT
+ cby_4__2_/Test_en_W_out grid_clb_4__2_/Test_en_E_out cby_4__2_/Test_en_W_out cby_3__2_/Test_en_W_in
+ VGND VPWR cbx_4__1_/REGIN_FEEDTHROUGH grid_clb_4__2_/bottom_width_0_height_0__pin_51_
+ cby_3__2_/ccff_tail cby_4__2_/ccff_head cbx_4__1_/clk_1_N_out cbx_4__1_/clk_1_N_out
+ cby_4__2_/prog_clk_0_W_in cbx_4__1_/prog_clk_1_N_out grid_clb_4__2_/prog_clk_0_N_out
+ cbx_4__1_/prog_clk_1_N_out cbx_4__1_/prog_clk_0_N_in grid_clb_4__2_/prog_clk_0_W_out
+ cby_4__2_/left_grid_pin_16_ cby_4__2_/left_grid_pin_17_ cby_4__2_/left_grid_pin_18_
+ cby_4__2_/left_grid_pin_19_ cby_4__2_/left_grid_pin_20_ cby_4__2_/left_grid_pin_21_
+ cby_4__2_/left_grid_pin_22_ cby_4__2_/left_grid_pin_23_ cby_4__2_/left_grid_pin_24_
+ cby_4__2_/left_grid_pin_25_ cby_4__2_/left_grid_pin_26_ cby_4__2_/left_grid_pin_27_
+ cby_4__2_/left_grid_pin_28_ cby_4__2_/left_grid_pin_29_ cby_4__2_/left_grid_pin_30_
+ cby_4__2_/left_grid_pin_31_ sb_4__1_/top_left_grid_pin_42_ sb_4__2_/bottom_left_grid_pin_42_
+ sb_4__1_/top_left_grid_pin_43_ sb_4__2_/bottom_left_grid_pin_43_ sb_4__1_/top_left_grid_pin_44_
+ sb_4__2_/bottom_left_grid_pin_44_ sb_4__1_/top_left_grid_pin_45_ sb_4__2_/bottom_left_grid_pin_45_
+ sb_4__1_/top_left_grid_pin_46_ sb_4__2_/bottom_left_grid_pin_46_ sb_4__1_/top_left_grid_pin_47_
+ sb_4__2_/bottom_left_grid_pin_47_ sb_4__1_/top_left_grid_pin_48_ sb_4__2_/bottom_left_grid_pin_48_
+ sb_4__1_/top_left_grid_pin_49_ sb_4__2_/bottom_left_grid_pin_49_ cbx_4__2_/bottom_grid_pin_0_
+ cbx_4__2_/bottom_grid_pin_10_ cbx_4__2_/bottom_grid_pin_11_ cbx_4__2_/bottom_grid_pin_12_
+ cbx_4__2_/bottom_grid_pin_13_ cbx_4__2_/bottom_grid_pin_14_ cbx_4__2_/bottom_grid_pin_15_
+ cbx_4__2_/bottom_grid_pin_1_ cbx_4__2_/bottom_grid_pin_2_ cbx_4__2_/REGOUT_FEEDTHROUGH
+ grid_clb_4__2_/top_width_0_height_0__pin_33_ sb_4__2_/left_bottom_grid_pin_34_ sb_3__2_/right_bottom_grid_pin_34_
+ sb_4__2_/left_bottom_grid_pin_35_ sb_3__2_/right_bottom_grid_pin_35_ sb_4__2_/left_bottom_grid_pin_36_
+ sb_3__2_/right_bottom_grid_pin_36_ sb_4__2_/left_bottom_grid_pin_37_ sb_3__2_/right_bottom_grid_pin_37_
+ sb_4__2_/left_bottom_grid_pin_38_ sb_3__2_/right_bottom_grid_pin_38_ sb_4__2_/left_bottom_grid_pin_39_
+ sb_3__2_/right_bottom_grid_pin_39_ cbx_4__2_/bottom_grid_pin_3_ sb_4__2_/left_bottom_grid_pin_40_
+ sb_3__2_/right_bottom_grid_pin_40_ sb_4__2_/left_bottom_grid_pin_41_ sb_3__2_/right_bottom_grid_pin_41_
+ cbx_4__2_/bottom_grid_pin_4_ cbx_4__2_/bottom_grid_pin_5_ cbx_4__2_/bottom_grid_pin_6_
+ cbx_4__2_/bottom_grid_pin_7_ cbx_4__2_/bottom_grid_pin_8_ cbx_4__2_/bottom_grid_pin_9_
+ grid_clb
Xsb_2__4_ sb_2__4_/Test_en_N_out sb_2__4_/Test_en_S_in VGND VPWR sb_2__4_/bottom_left_grid_pin_42_
+ sb_2__4_/bottom_left_grid_pin_43_ sb_2__4_/bottom_left_grid_pin_44_ sb_2__4_/bottom_left_grid_pin_45_
+ sb_2__4_/bottom_left_grid_pin_46_ sb_2__4_/bottom_left_grid_pin_47_ sb_2__4_/bottom_left_grid_pin_48_
+ sb_2__4_/bottom_left_grid_pin_49_ sb_2__4_/ccff_head sb_2__4_/ccff_tail sb_2__4_/chanx_left_in[0]
+ sb_2__4_/chanx_left_in[10] sb_2__4_/chanx_left_in[11] sb_2__4_/chanx_left_in[12]
+ sb_2__4_/chanx_left_in[13] sb_2__4_/chanx_left_in[14] sb_2__4_/chanx_left_in[15]
+ sb_2__4_/chanx_left_in[16] sb_2__4_/chanx_left_in[17] sb_2__4_/chanx_left_in[18]
+ sb_2__4_/chanx_left_in[19] sb_2__4_/chanx_left_in[1] sb_2__4_/chanx_left_in[2] sb_2__4_/chanx_left_in[3]
+ sb_2__4_/chanx_left_in[4] sb_2__4_/chanx_left_in[5] sb_2__4_/chanx_left_in[6] sb_2__4_/chanx_left_in[7]
+ sb_2__4_/chanx_left_in[8] sb_2__4_/chanx_left_in[9] sb_2__4_/chanx_left_out[0] sb_2__4_/chanx_left_out[10]
+ sb_2__4_/chanx_left_out[11] sb_2__4_/chanx_left_out[12] sb_2__4_/chanx_left_out[13]
+ sb_2__4_/chanx_left_out[14] sb_2__4_/chanx_left_out[15] sb_2__4_/chanx_left_out[16]
+ sb_2__4_/chanx_left_out[17] sb_2__4_/chanx_left_out[18] sb_2__4_/chanx_left_out[19]
+ sb_2__4_/chanx_left_out[1] sb_2__4_/chanx_left_out[2] sb_2__4_/chanx_left_out[3]
+ sb_2__4_/chanx_left_out[4] sb_2__4_/chanx_left_out[5] sb_2__4_/chanx_left_out[6]
+ sb_2__4_/chanx_left_out[7] sb_2__4_/chanx_left_out[8] sb_2__4_/chanx_left_out[9]
+ sb_2__4_/chanx_right_in[0] sb_2__4_/chanx_right_in[10] sb_2__4_/chanx_right_in[11]
+ sb_2__4_/chanx_right_in[12] sb_2__4_/chanx_right_in[13] sb_2__4_/chanx_right_in[14]
+ sb_2__4_/chanx_right_in[15] sb_2__4_/chanx_right_in[16] sb_2__4_/chanx_right_in[17]
+ sb_2__4_/chanx_right_in[18] sb_2__4_/chanx_right_in[19] sb_2__4_/chanx_right_in[1]
+ sb_2__4_/chanx_right_in[2] sb_2__4_/chanx_right_in[3] sb_2__4_/chanx_right_in[4]
+ sb_2__4_/chanx_right_in[5] sb_2__4_/chanx_right_in[6] sb_2__4_/chanx_right_in[7]
+ sb_2__4_/chanx_right_in[8] sb_2__4_/chanx_right_in[9] cbx_3__4_/chanx_left_in[0]
+ cbx_3__4_/chanx_left_in[10] cbx_3__4_/chanx_left_in[11] cbx_3__4_/chanx_left_in[12]
+ cbx_3__4_/chanx_left_in[13] cbx_3__4_/chanx_left_in[14] cbx_3__4_/chanx_left_in[15]
+ cbx_3__4_/chanx_left_in[16] cbx_3__4_/chanx_left_in[17] cbx_3__4_/chanx_left_in[18]
+ cbx_3__4_/chanx_left_in[19] cbx_3__4_/chanx_left_in[1] cbx_3__4_/chanx_left_in[2]
+ cbx_3__4_/chanx_left_in[3] cbx_3__4_/chanx_left_in[4] cbx_3__4_/chanx_left_in[5]
+ cbx_3__4_/chanx_left_in[6] cbx_3__4_/chanx_left_in[7] cbx_3__4_/chanx_left_in[8]
+ cbx_3__4_/chanx_left_in[9] cby_2__4_/chany_top_out[0] cby_2__4_/chany_top_out[10]
+ cby_2__4_/chany_top_out[11] cby_2__4_/chany_top_out[12] cby_2__4_/chany_top_out[13]
+ cby_2__4_/chany_top_out[14] cby_2__4_/chany_top_out[15] cby_2__4_/chany_top_out[16]
+ cby_2__4_/chany_top_out[17] cby_2__4_/chany_top_out[18] cby_2__4_/chany_top_out[19]
+ cby_2__4_/chany_top_out[1] cby_2__4_/chany_top_out[2] cby_2__4_/chany_top_out[3]
+ cby_2__4_/chany_top_out[4] cby_2__4_/chany_top_out[5] cby_2__4_/chany_top_out[6]
+ cby_2__4_/chany_top_out[7] cby_2__4_/chany_top_out[8] cby_2__4_/chany_top_out[9]
+ cby_2__4_/chany_top_in[0] cby_2__4_/chany_top_in[10] cby_2__4_/chany_top_in[11]
+ cby_2__4_/chany_top_in[12] cby_2__4_/chany_top_in[13] cby_2__4_/chany_top_in[14]
+ cby_2__4_/chany_top_in[15] cby_2__4_/chany_top_in[16] cby_2__4_/chany_top_in[17]
+ cby_2__4_/chany_top_in[18] cby_2__4_/chany_top_in[19] cby_2__4_/chany_top_in[1]
+ cby_2__4_/chany_top_in[2] cby_2__4_/chany_top_in[3] cby_2__4_/chany_top_in[4] cby_2__4_/chany_top_in[5]
+ cby_2__4_/chany_top_in[6] cby_2__4_/chany_top_in[7] cby_2__4_/chany_top_in[8] cby_2__4_/chany_top_in[9]
+ sb_2__4_/chany_top_in[0] sb_2__4_/chany_top_in[10] sb_2__4_/chany_top_in[11] sb_2__4_/chany_top_in[12]
+ sb_2__4_/chany_top_in[13] sb_2__4_/chany_top_in[14] sb_2__4_/chany_top_in[15] sb_2__4_/chany_top_in[16]
+ sb_2__4_/chany_top_in[17] sb_2__4_/chany_top_in[18] sb_2__4_/chany_top_in[19] sb_2__4_/chany_top_in[1]
+ sb_2__4_/chany_top_in[2] sb_2__4_/chany_top_in[3] sb_2__4_/chany_top_in[4] sb_2__4_/chany_top_in[5]
+ sb_2__4_/chany_top_in[6] sb_2__4_/chany_top_in[7] sb_2__4_/chany_top_in[8] sb_2__4_/chany_top_in[9]
+ sb_2__4_/chany_top_out[0] sb_2__4_/chany_top_out[10] sb_2__4_/chany_top_out[11]
+ sb_2__4_/chany_top_out[12] sb_2__4_/chany_top_out[13] sb_2__4_/chany_top_out[14]
+ sb_2__4_/chany_top_out[15] sb_2__4_/chany_top_out[16] sb_2__4_/chany_top_out[17]
+ sb_2__4_/chany_top_out[18] sb_2__4_/chany_top_out[19] sb_2__4_/chany_top_out[1]
+ sb_2__4_/chany_top_out[2] sb_2__4_/chany_top_out[3] sb_2__4_/chany_top_out[4] sb_2__4_/chany_top_out[5]
+ sb_2__4_/chany_top_out[6] sb_2__4_/chany_top_out[7] sb_2__4_/chany_top_out[8] sb_2__4_/chany_top_out[9]
+ sb_2__4_/clk_1_E_out sb_2__4_/clk_1_N_in sb_2__4_/clk_1_W_out sb_2__4_/clk_2_E_out
+ sb_2__4_/clk_2_N_in sb_2__4_/clk_2_N_out sb_2__4_/clk_2_S_out sb_2__4_/clk_2_W_out
+ sb_2__4_/clk_3_E_out sb_2__4_/clk_3_N_in sb_2__4_/clk_3_N_out sb_2__4_/clk_3_S_out
+ sb_2__4_/clk_3_W_out sb_2__4_/left_bottom_grid_pin_34_ sb_2__4_/left_bottom_grid_pin_35_
+ sb_2__4_/left_bottom_grid_pin_36_ sb_2__4_/left_bottom_grid_pin_37_ sb_2__4_/left_bottom_grid_pin_38_
+ sb_2__4_/left_bottom_grid_pin_39_ sb_2__4_/left_bottom_grid_pin_40_ sb_2__4_/left_bottom_grid_pin_41_
+ sb_2__4_/prog_clk_0_N_in sb_2__4_/prog_clk_1_E_out sb_2__4_/prog_clk_1_N_in sb_2__4_/prog_clk_1_W_out
+ sb_2__4_/prog_clk_2_E_out sb_2__4_/prog_clk_2_N_in sb_2__4_/prog_clk_2_N_out sb_2__4_/prog_clk_2_S_out
+ sb_2__4_/prog_clk_2_W_out sb_2__4_/prog_clk_3_E_out sb_2__4_/prog_clk_3_N_in sb_2__4_/prog_clk_3_N_out
+ sb_2__4_/prog_clk_3_S_out sb_2__4_/prog_clk_3_W_out sb_2__4_/right_bottom_grid_pin_34_
+ sb_2__4_/right_bottom_grid_pin_35_ sb_2__4_/right_bottom_grid_pin_36_ sb_2__4_/right_bottom_grid_pin_37_
+ sb_2__4_/right_bottom_grid_pin_38_ sb_2__4_/right_bottom_grid_pin_39_ sb_2__4_/right_bottom_grid_pin_40_
+ sb_2__4_/right_bottom_grid_pin_41_ sb_2__4_/top_left_grid_pin_42_ sb_2__4_/top_left_grid_pin_43_
+ sb_2__4_/top_left_grid_pin_44_ sb_2__4_/top_left_grid_pin_45_ sb_2__4_/top_left_grid_pin_46_
+ sb_2__4_/top_left_grid_pin_47_ sb_2__4_/top_left_grid_pin_48_ sb_2__4_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_8__3_ IO_ISOL_N VGND VPWR cby_8__3_/ccff_head sb_8__2_/ccff_head sb_8__2_/chany_top_out[0]
+ sb_8__2_/chany_top_out[10] sb_8__2_/chany_top_out[11] sb_8__2_/chany_top_out[12]
+ sb_8__2_/chany_top_out[13] sb_8__2_/chany_top_out[14] sb_8__2_/chany_top_out[15]
+ sb_8__2_/chany_top_out[16] sb_8__2_/chany_top_out[17] sb_8__2_/chany_top_out[18]
+ sb_8__2_/chany_top_out[19] sb_8__2_/chany_top_out[1] sb_8__2_/chany_top_out[2] sb_8__2_/chany_top_out[3]
+ sb_8__2_/chany_top_out[4] sb_8__2_/chany_top_out[5] sb_8__2_/chany_top_out[6] sb_8__2_/chany_top_out[7]
+ sb_8__2_/chany_top_out[8] sb_8__2_/chany_top_out[9] sb_8__2_/chany_top_in[0] sb_8__2_/chany_top_in[10]
+ sb_8__2_/chany_top_in[11] sb_8__2_/chany_top_in[12] sb_8__2_/chany_top_in[13] sb_8__2_/chany_top_in[14]
+ sb_8__2_/chany_top_in[15] sb_8__2_/chany_top_in[16] sb_8__2_/chany_top_in[17] sb_8__2_/chany_top_in[18]
+ sb_8__2_/chany_top_in[19] sb_8__2_/chany_top_in[1] sb_8__2_/chany_top_in[2] sb_8__2_/chany_top_in[3]
+ sb_8__2_/chany_top_in[4] sb_8__2_/chany_top_in[5] sb_8__2_/chany_top_in[6] sb_8__2_/chany_top_in[7]
+ sb_8__2_/chany_top_in[8] sb_8__2_/chany_top_in[9] cby_8__3_/chany_top_in[0] cby_8__3_/chany_top_in[10]
+ cby_8__3_/chany_top_in[11] cby_8__3_/chany_top_in[12] cby_8__3_/chany_top_in[13]
+ cby_8__3_/chany_top_in[14] cby_8__3_/chany_top_in[15] cby_8__3_/chany_top_in[16]
+ cby_8__3_/chany_top_in[17] cby_8__3_/chany_top_in[18] cby_8__3_/chany_top_in[19]
+ cby_8__3_/chany_top_in[1] cby_8__3_/chany_top_in[2] cby_8__3_/chany_top_in[3] cby_8__3_/chany_top_in[4]
+ cby_8__3_/chany_top_in[5] cby_8__3_/chany_top_in[6] cby_8__3_/chany_top_in[7] cby_8__3_/chany_top_in[8]
+ cby_8__3_/chany_top_in[9] cby_8__3_/chany_top_out[0] cby_8__3_/chany_top_out[10]
+ cby_8__3_/chany_top_out[11] cby_8__3_/chany_top_out[12] cby_8__3_/chany_top_out[13]
+ cby_8__3_/chany_top_out[14] cby_8__3_/chany_top_out[15] cby_8__3_/chany_top_out[16]
+ cby_8__3_/chany_top_out[17] cby_8__3_/chany_top_out[18] cby_8__3_/chany_top_out[19]
+ cby_8__3_/chany_top_out[1] cby_8__3_/chany_top_out[2] cby_8__3_/chany_top_out[3]
+ cby_8__3_/chany_top_out[4] cby_8__3_/chany_top_out[5] cby_8__3_/chany_top_out[6]
+ cby_8__3_/chany_top_out[7] cby_8__3_/chany_top_out[8] cby_8__3_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
+ cby_8__3_/left_grid_pin_16_ cby_8__3_/left_grid_pin_17_ cby_8__3_/left_grid_pin_18_
+ cby_8__3_/left_grid_pin_19_ cby_8__3_/left_grid_pin_20_ cby_8__3_/left_grid_pin_21_
+ cby_8__3_/left_grid_pin_22_ cby_8__3_/left_grid_pin_23_ cby_8__3_/left_grid_pin_24_
+ cby_8__3_/left_grid_pin_25_ cby_8__3_/left_grid_pin_26_ cby_8__3_/left_grid_pin_27_
+ cby_8__3_/left_grid_pin_28_ cby_8__3_/left_grid_pin_29_ cby_8__3_/left_grid_pin_30_
+ cby_8__3_/left_grid_pin_31_ cby_8__3_/right_grid_pin_0_ sb_8__2_/top_right_grid_pin_1_
+ sb_8__3_/bottom_right_grid_pin_1_ cby_8__3_/prog_clk_0_N_out sb_8__2_/prog_clk_0_N_in
+ cby_8__3_/prog_clk_0_W_in cby_8__3_/right_grid_pin_0_ cby_2__1_
Xcbx_8__4_ cbx_8__4_/REGIN_FEEDTHROUGH cbx_8__4_/REGOUT_FEEDTHROUGH cbx_8__4_/SC_IN_BOT
+ cbx_8__4_/SC_IN_TOP cbx_8__4_/SC_OUT_BOT cbx_8__4_/SC_OUT_TOP VGND VPWR cbx_8__4_/bottom_grid_pin_0_
+ cbx_8__4_/bottom_grid_pin_10_ cbx_8__4_/bottom_grid_pin_11_ cbx_8__4_/bottom_grid_pin_12_
+ cbx_8__4_/bottom_grid_pin_13_ cbx_8__4_/bottom_grid_pin_14_ cbx_8__4_/bottom_grid_pin_15_
+ cbx_8__4_/bottom_grid_pin_1_ cbx_8__4_/bottom_grid_pin_2_ cbx_8__4_/bottom_grid_pin_3_
+ cbx_8__4_/bottom_grid_pin_4_ cbx_8__4_/bottom_grid_pin_5_ cbx_8__4_/bottom_grid_pin_6_
+ cbx_8__4_/bottom_grid_pin_7_ cbx_8__4_/bottom_grid_pin_8_ cbx_8__4_/bottom_grid_pin_9_
+ sb_8__4_/ccff_tail sb_7__4_/ccff_head cbx_8__4_/chanx_left_in[0] cbx_8__4_/chanx_left_in[10]
+ cbx_8__4_/chanx_left_in[11] cbx_8__4_/chanx_left_in[12] cbx_8__4_/chanx_left_in[13]
+ cbx_8__4_/chanx_left_in[14] cbx_8__4_/chanx_left_in[15] cbx_8__4_/chanx_left_in[16]
+ cbx_8__4_/chanx_left_in[17] cbx_8__4_/chanx_left_in[18] cbx_8__4_/chanx_left_in[19]
+ cbx_8__4_/chanx_left_in[1] cbx_8__4_/chanx_left_in[2] cbx_8__4_/chanx_left_in[3]
+ cbx_8__4_/chanx_left_in[4] cbx_8__4_/chanx_left_in[5] cbx_8__4_/chanx_left_in[6]
+ cbx_8__4_/chanx_left_in[7] cbx_8__4_/chanx_left_in[8] cbx_8__4_/chanx_left_in[9]
+ sb_7__4_/chanx_right_in[0] sb_7__4_/chanx_right_in[10] sb_7__4_/chanx_right_in[11]
+ sb_7__4_/chanx_right_in[12] sb_7__4_/chanx_right_in[13] sb_7__4_/chanx_right_in[14]
+ sb_7__4_/chanx_right_in[15] sb_7__4_/chanx_right_in[16] sb_7__4_/chanx_right_in[17]
+ sb_7__4_/chanx_right_in[18] sb_7__4_/chanx_right_in[19] sb_7__4_/chanx_right_in[1]
+ sb_7__4_/chanx_right_in[2] sb_7__4_/chanx_right_in[3] sb_7__4_/chanx_right_in[4]
+ sb_7__4_/chanx_right_in[5] sb_7__4_/chanx_right_in[6] sb_7__4_/chanx_right_in[7]
+ sb_7__4_/chanx_right_in[8] sb_7__4_/chanx_right_in[9] sb_8__4_/chanx_left_out[0]
+ sb_8__4_/chanx_left_out[10] sb_8__4_/chanx_left_out[11] sb_8__4_/chanx_left_out[12]
+ sb_8__4_/chanx_left_out[13] sb_8__4_/chanx_left_out[14] sb_8__4_/chanx_left_out[15]
+ sb_8__4_/chanx_left_out[16] sb_8__4_/chanx_left_out[17] sb_8__4_/chanx_left_out[18]
+ sb_8__4_/chanx_left_out[19] sb_8__4_/chanx_left_out[1] sb_8__4_/chanx_left_out[2]
+ sb_8__4_/chanx_left_out[3] sb_8__4_/chanx_left_out[4] sb_8__4_/chanx_left_out[5]
+ sb_8__4_/chanx_left_out[6] sb_8__4_/chanx_left_out[7] sb_8__4_/chanx_left_out[8]
+ sb_8__4_/chanx_left_out[9] sb_8__4_/chanx_left_in[0] sb_8__4_/chanx_left_in[10]
+ sb_8__4_/chanx_left_in[11] sb_8__4_/chanx_left_in[12] sb_8__4_/chanx_left_in[13]
+ sb_8__4_/chanx_left_in[14] sb_8__4_/chanx_left_in[15] sb_8__4_/chanx_left_in[16]
+ sb_8__4_/chanx_left_in[17] sb_8__4_/chanx_left_in[18] sb_8__4_/chanx_left_in[19]
+ sb_8__4_/chanx_left_in[1] sb_8__4_/chanx_left_in[2] sb_8__4_/chanx_left_in[3] sb_8__4_/chanx_left_in[4]
+ sb_8__4_/chanx_left_in[5] sb_8__4_/chanx_left_in[6] sb_8__4_/chanx_left_in[7] sb_8__4_/chanx_left_in[8]
+ sb_8__4_/chanx_left_in[9] cbx_8__4_/clk_1_N_out cbx_8__4_/clk_1_S_out cbx_8__4_/clk_1_W_in
+ cbx_8__4_/clk_2_E_out cbx_8__4_/clk_2_W_in cbx_8__4_/clk_2_W_out cbx_8__4_/clk_3_E_out
+ cbx_8__4_/clk_3_W_in cbx_8__4_/clk_3_W_out cbx_8__4_/prog_clk_0_N_in cbx_8__4_/prog_clk_0_W_out
+ cbx_8__4_/prog_clk_1_N_out cbx_8__4_/prog_clk_1_S_out cbx_8__4_/prog_clk_1_W_in
+ cbx_8__4_/prog_clk_2_E_out cbx_8__4_/prog_clk_2_W_in cbx_8__4_/prog_clk_2_W_out
+ cbx_8__4_/prog_clk_3_E_out cbx_8__4_/prog_clk_3_W_in cbx_8__4_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_1__8_ cby_1__8_/Test_en_W_in cby_1__8_/Test_en_E_out cby_1__8_/Test_en_N_out
+ cby_1__8_/Test_en_W_in cby_1__8_/Test_en_W_in cby_1__8_/Test_en_W_out VGND VPWR
+ cby_1__8_/ccff_head cby_1__8_/ccff_tail sb_1__7_/chany_top_out[0] sb_1__7_/chany_top_out[10]
+ sb_1__7_/chany_top_out[11] sb_1__7_/chany_top_out[12] sb_1__7_/chany_top_out[13]
+ sb_1__7_/chany_top_out[14] sb_1__7_/chany_top_out[15] sb_1__7_/chany_top_out[16]
+ sb_1__7_/chany_top_out[17] sb_1__7_/chany_top_out[18] sb_1__7_/chany_top_out[19]
+ sb_1__7_/chany_top_out[1] sb_1__7_/chany_top_out[2] sb_1__7_/chany_top_out[3] sb_1__7_/chany_top_out[4]
+ sb_1__7_/chany_top_out[5] sb_1__7_/chany_top_out[6] sb_1__7_/chany_top_out[7] sb_1__7_/chany_top_out[8]
+ sb_1__7_/chany_top_out[9] sb_1__7_/chany_top_in[0] sb_1__7_/chany_top_in[10] sb_1__7_/chany_top_in[11]
+ sb_1__7_/chany_top_in[12] sb_1__7_/chany_top_in[13] sb_1__7_/chany_top_in[14] sb_1__7_/chany_top_in[15]
+ sb_1__7_/chany_top_in[16] sb_1__7_/chany_top_in[17] sb_1__7_/chany_top_in[18] sb_1__7_/chany_top_in[19]
+ sb_1__7_/chany_top_in[1] sb_1__7_/chany_top_in[2] sb_1__7_/chany_top_in[3] sb_1__7_/chany_top_in[4]
+ sb_1__7_/chany_top_in[5] sb_1__7_/chany_top_in[6] sb_1__7_/chany_top_in[7] sb_1__7_/chany_top_in[8]
+ sb_1__7_/chany_top_in[9] cby_1__8_/chany_top_in[0] cby_1__8_/chany_top_in[10] cby_1__8_/chany_top_in[11]
+ cby_1__8_/chany_top_in[12] cby_1__8_/chany_top_in[13] cby_1__8_/chany_top_in[14]
+ cby_1__8_/chany_top_in[15] cby_1__8_/chany_top_in[16] cby_1__8_/chany_top_in[17]
+ cby_1__8_/chany_top_in[18] cby_1__8_/chany_top_in[19] cby_1__8_/chany_top_in[1]
+ cby_1__8_/chany_top_in[2] cby_1__8_/chany_top_in[3] cby_1__8_/chany_top_in[4] cby_1__8_/chany_top_in[5]
+ cby_1__8_/chany_top_in[6] cby_1__8_/chany_top_in[7] cby_1__8_/chany_top_in[8] cby_1__8_/chany_top_in[9]
+ cby_1__8_/chany_top_out[0] cby_1__8_/chany_top_out[10] cby_1__8_/chany_top_out[11]
+ cby_1__8_/chany_top_out[12] cby_1__8_/chany_top_out[13] cby_1__8_/chany_top_out[14]
+ cby_1__8_/chany_top_out[15] cby_1__8_/chany_top_out[16] cby_1__8_/chany_top_out[17]
+ cby_1__8_/chany_top_out[18] cby_1__8_/chany_top_out[19] cby_1__8_/chany_top_out[1]
+ cby_1__8_/chany_top_out[2] cby_1__8_/chany_top_out[3] cby_1__8_/chany_top_out[4]
+ cby_1__8_/chany_top_out[5] cby_1__8_/chany_top_out[6] cby_1__8_/chany_top_out[7]
+ cby_1__8_/chany_top_out[8] cby_1__8_/chany_top_out[9] cby_1__8_/clk_2_N_out cby_1__8_/clk_2_S_in
+ cby_1__8_/clk_2_S_out cby_1__8_/clk_3_N_out cby_1__8_/clk_3_S_in cby_1__8_/clk_3_S_out
+ cby_1__8_/left_grid_pin_16_ cby_1__8_/left_grid_pin_17_ cby_1__8_/left_grid_pin_18_
+ cby_1__8_/left_grid_pin_19_ cby_1__8_/left_grid_pin_20_ cby_1__8_/left_grid_pin_21_
+ cby_1__8_/left_grid_pin_22_ cby_1__8_/left_grid_pin_23_ cby_1__8_/left_grid_pin_24_
+ cby_1__8_/left_grid_pin_25_ cby_1__8_/left_grid_pin_26_ cby_1__8_/left_grid_pin_27_
+ cby_1__8_/left_grid_pin_28_ cby_1__8_/left_grid_pin_29_ cby_1__8_/left_grid_pin_30_
+ cby_1__8_/left_grid_pin_31_ sb_1__8_/prog_clk_0_S_in sb_1__7_/prog_clk_0_N_in cby_1__8_/prog_clk_0_W_in
+ cby_1__8_/prog_clk_2_N_out cby_1__8_/prog_clk_2_S_in cby_1__8_/prog_clk_2_S_out
+ cby_1__8_/prog_clk_3_N_out cby_1__8_/prog_clk_3_S_in cby_1__8_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_7__4_ cbx_7__4_/SC_OUT_BOT cbx_7__3_/SC_IN_TOP grid_clb_7__4_/SC_OUT_TOP
+ cby_6__4_/Test_en_E_out cby_7__4_/Test_en_W_in cby_6__4_/Test_en_E_out grid_clb_7__4_/Test_en_W_out
+ VGND VPWR cbx_7__3_/REGIN_FEEDTHROUGH grid_clb_7__4_/bottom_width_0_height_0__pin_51_
+ cby_6__4_/ccff_tail cby_7__4_/ccff_head cbx_7__3_/clk_1_N_out cbx_7__3_/clk_1_N_out
+ cby_7__4_/prog_clk_0_W_in cbx_7__3_/prog_clk_1_N_out grid_clb_7__4_/prog_clk_0_N_out
+ cbx_7__3_/prog_clk_1_N_out cbx_7__3_/prog_clk_0_N_in grid_clb_7__4_/prog_clk_0_W_out
+ cby_7__4_/left_grid_pin_16_ cby_7__4_/left_grid_pin_17_ cby_7__4_/left_grid_pin_18_
+ cby_7__4_/left_grid_pin_19_ cby_7__4_/left_grid_pin_20_ cby_7__4_/left_grid_pin_21_
+ cby_7__4_/left_grid_pin_22_ cby_7__4_/left_grid_pin_23_ cby_7__4_/left_grid_pin_24_
+ cby_7__4_/left_grid_pin_25_ cby_7__4_/left_grid_pin_26_ cby_7__4_/left_grid_pin_27_
+ cby_7__4_/left_grid_pin_28_ cby_7__4_/left_grid_pin_29_ cby_7__4_/left_grid_pin_30_
+ cby_7__4_/left_grid_pin_31_ sb_7__3_/top_left_grid_pin_42_ sb_7__4_/bottom_left_grid_pin_42_
+ sb_7__3_/top_left_grid_pin_43_ sb_7__4_/bottom_left_grid_pin_43_ sb_7__3_/top_left_grid_pin_44_
+ sb_7__4_/bottom_left_grid_pin_44_ sb_7__3_/top_left_grid_pin_45_ sb_7__4_/bottom_left_grid_pin_45_
+ sb_7__3_/top_left_grid_pin_46_ sb_7__4_/bottom_left_grid_pin_46_ sb_7__3_/top_left_grid_pin_47_
+ sb_7__4_/bottom_left_grid_pin_47_ sb_7__3_/top_left_grid_pin_48_ sb_7__4_/bottom_left_grid_pin_48_
+ sb_7__3_/top_left_grid_pin_49_ sb_7__4_/bottom_left_grid_pin_49_ cbx_7__4_/bottom_grid_pin_0_
+ cbx_7__4_/bottom_grid_pin_10_ cbx_7__4_/bottom_grid_pin_11_ cbx_7__4_/bottom_grid_pin_12_
+ cbx_7__4_/bottom_grid_pin_13_ cbx_7__4_/bottom_grid_pin_14_ cbx_7__4_/bottom_grid_pin_15_
+ cbx_7__4_/bottom_grid_pin_1_ cbx_7__4_/bottom_grid_pin_2_ cbx_7__4_/REGOUT_FEEDTHROUGH
+ grid_clb_7__4_/top_width_0_height_0__pin_33_ sb_7__4_/left_bottom_grid_pin_34_ sb_6__4_/right_bottom_grid_pin_34_
+ sb_7__4_/left_bottom_grid_pin_35_ sb_6__4_/right_bottom_grid_pin_35_ sb_7__4_/left_bottom_grid_pin_36_
+ sb_6__4_/right_bottom_grid_pin_36_ sb_7__4_/left_bottom_grid_pin_37_ sb_6__4_/right_bottom_grid_pin_37_
+ sb_7__4_/left_bottom_grid_pin_38_ sb_6__4_/right_bottom_grid_pin_38_ sb_7__4_/left_bottom_grid_pin_39_
+ sb_6__4_/right_bottom_grid_pin_39_ cbx_7__4_/bottom_grid_pin_3_ sb_7__4_/left_bottom_grid_pin_40_
+ sb_6__4_/right_bottom_grid_pin_40_ sb_7__4_/left_bottom_grid_pin_41_ sb_6__4_/right_bottom_grid_pin_41_
+ cbx_7__4_/bottom_grid_pin_4_ cbx_7__4_/bottom_grid_pin_5_ cbx_7__4_/bottom_grid_pin_6_
+ cbx_7__4_/bottom_grid_pin_7_ cbx_7__4_/bottom_grid_pin_8_ cbx_7__4_/bottom_grid_pin_9_
+ grid_clb
Xgrid_clb_4__1_ cbx_4__0_/SC_OUT_TOP grid_clb_4__1_/SC_OUT_BOT cbx_4__1_/SC_IN_BOT
+ cby_4__1_/Test_en_W_out grid_clb_4__1_/Test_en_E_out cby_4__1_/Test_en_W_out cby_3__1_/Test_en_W_in
+ VGND VPWR grid_clb_4__1_/bottom_width_0_height_0__pin_50_ grid_clb_4__1_/bottom_width_0_height_0__pin_51_
+ cby_3__1_/ccff_tail cby_4__1_/ccff_head cbx_4__1_/clk_1_S_out cbx_4__1_/clk_1_S_out
+ cby_4__1_/prog_clk_0_W_in cbx_4__1_/prog_clk_1_S_out grid_clb_4__1_/prog_clk_0_N_out
+ cbx_4__1_/prog_clk_1_S_out cbx_4__0_/prog_clk_0_N_in grid_clb_4__1_/prog_clk_0_W_out
+ cby_4__1_/left_grid_pin_16_ cby_4__1_/left_grid_pin_17_ cby_4__1_/left_grid_pin_18_
+ cby_4__1_/left_grid_pin_19_ cby_4__1_/left_grid_pin_20_ cby_4__1_/left_grid_pin_21_
+ cby_4__1_/left_grid_pin_22_ cby_4__1_/left_grid_pin_23_ cby_4__1_/left_grid_pin_24_
+ cby_4__1_/left_grid_pin_25_ cby_4__1_/left_grid_pin_26_ cby_4__1_/left_grid_pin_27_
+ cby_4__1_/left_grid_pin_28_ cby_4__1_/left_grid_pin_29_ cby_4__1_/left_grid_pin_30_
+ cby_4__1_/left_grid_pin_31_ sb_4__0_/top_left_grid_pin_42_ sb_4__1_/bottom_left_grid_pin_42_
+ sb_4__0_/top_left_grid_pin_43_ sb_4__1_/bottom_left_grid_pin_43_ sb_4__0_/top_left_grid_pin_44_
+ sb_4__1_/bottom_left_grid_pin_44_ sb_4__0_/top_left_grid_pin_45_ sb_4__1_/bottom_left_grid_pin_45_
+ sb_4__0_/top_left_grid_pin_46_ sb_4__1_/bottom_left_grid_pin_46_ sb_4__0_/top_left_grid_pin_47_
+ sb_4__1_/bottom_left_grid_pin_47_ sb_4__0_/top_left_grid_pin_48_ sb_4__1_/bottom_left_grid_pin_48_
+ sb_4__0_/top_left_grid_pin_49_ sb_4__1_/bottom_left_grid_pin_49_ cbx_4__1_/bottom_grid_pin_0_
+ cbx_4__1_/bottom_grid_pin_10_ cbx_4__1_/bottom_grid_pin_11_ cbx_4__1_/bottom_grid_pin_12_
+ cbx_4__1_/bottom_grid_pin_13_ cbx_4__1_/bottom_grid_pin_14_ cbx_4__1_/bottom_grid_pin_15_
+ cbx_4__1_/bottom_grid_pin_1_ cbx_4__1_/bottom_grid_pin_2_ cbx_4__1_/REGOUT_FEEDTHROUGH
+ grid_clb_4__1_/top_width_0_height_0__pin_33_ sb_4__1_/left_bottom_grid_pin_34_ sb_3__1_/right_bottom_grid_pin_34_
+ sb_4__1_/left_bottom_grid_pin_35_ sb_3__1_/right_bottom_grid_pin_35_ sb_4__1_/left_bottom_grid_pin_36_
+ sb_3__1_/right_bottom_grid_pin_36_ sb_4__1_/left_bottom_grid_pin_37_ sb_3__1_/right_bottom_grid_pin_37_
+ sb_4__1_/left_bottom_grid_pin_38_ sb_3__1_/right_bottom_grid_pin_38_ sb_4__1_/left_bottom_grid_pin_39_
+ sb_3__1_/right_bottom_grid_pin_39_ cbx_4__1_/bottom_grid_pin_3_ sb_4__1_/left_bottom_grid_pin_40_
+ sb_3__1_/right_bottom_grid_pin_40_ sb_4__1_/left_bottom_grid_pin_41_ sb_3__1_/right_bottom_grid_pin_41_
+ cbx_4__1_/bottom_grid_pin_4_ cbx_4__1_/bottom_grid_pin_5_ cbx_4__1_/bottom_grid_pin_6_
+ cbx_4__1_/bottom_grid_pin_7_ cbx_4__1_/bottom_grid_pin_8_ cbx_4__1_/bottom_grid_pin_9_
+ grid_clb
Xcbx_5__1_ cbx_5__1_/REGIN_FEEDTHROUGH cbx_5__1_/REGOUT_FEEDTHROUGH cbx_5__1_/SC_IN_BOT
+ cbx_5__1_/SC_IN_TOP cbx_5__1_/SC_OUT_BOT cbx_5__1_/SC_OUT_TOP VGND VPWR cbx_5__1_/bottom_grid_pin_0_
+ cbx_5__1_/bottom_grid_pin_10_ cbx_5__1_/bottom_grid_pin_11_ cbx_5__1_/bottom_grid_pin_12_
+ cbx_5__1_/bottom_grid_pin_13_ cbx_5__1_/bottom_grid_pin_14_ cbx_5__1_/bottom_grid_pin_15_
+ cbx_5__1_/bottom_grid_pin_1_ cbx_5__1_/bottom_grid_pin_2_ cbx_5__1_/bottom_grid_pin_3_
+ cbx_5__1_/bottom_grid_pin_4_ cbx_5__1_/bottom_grid_pin_5_ cbx_5__1_/bottom_grid_pin_6_
+ cbx_5__1_/bottom_grid_pin_7_ cbx_5__1_/bottom_grid_pin_8_ cbx_5__1_/bottom_grid_pin_9_
+ sb_5__1_/ccff_tail sb_4__1_/ccff_head cbx_5__1_/chanx_left_in[0] cbx_5__1_/chanx_left_in[10]
+ cbx_5__1_/chanx_left_in[11] cbx_5__1_/chanx_left_in[12] cbx_5__1_/chanx_left_in[13]
+ cbx_5__1_/chanx_left_in[14] cbx_5__1_/chanx_left_in[15] cbx_5__1_/chanx_left_in[16]
+ cbx_5__1_/chanx_left_in[17] cbx_5__1_/chanx_left_in[18] cbx_5__1_/chanx_left_in[19]
+ cbx_5__1_/chanx_left_in[1] cbx_5__1_/chanx_left_in[2] cbx_5__1_/chanx_left_in[3]
+ cbx_5__1_/chanx_left_in[4] cbx_5__1_/chanx_left_in[5] cbx_5__1_/chanx_left_in[6]
+ cbx_5__1_/chanx_left_in[7] cbx_5__1_/chanx_left_in[8] cbx_5__1_/chanx_left_in[9]
+ sb_4__1_/chanx_right_in[0] sb_4__1_/chanx_right_in[10] sb_4__1_/chanx_right_in[11]
+ sb_4__1_/chanx_right_in[12] sb_4__1_/chanx_right_in[13] sb_4__1_/chanx_right_in[14]
+ sb_4__1_/chanx_right_in[15] sb_4__1_/chanx_right_in[16] sb_4__1_/chanx_right_in[17]
+ sb_4__1_/chanx_right_in[18] sb_4__1_/chanx_right_in[19] sb_4__1_/chanx_right_in[1]
+ sb_4__1_/chanx_right_in[2] sb_4__1_/chanx_right_in[3] sb_4__1_/chanx_right_in[4]
+ sb_4__1_/chanx_right_in[5] sb_4__1_/chanx_right_in[6] sb_4__1_/chanx_right_in[7]
+ sb_4__1_/chanx_right_in[8] sb_4__1_/chanx_right_in[9] sb_5__1_/chanx_left_out[0]
+ sb_5__1_/chanx_left_out[10] sb_5__1_/chanx_left_out[11] sb_5__1_/chanx_left_out[12]
+ sb_5__1_/chanx_left_out[13] sb_5__1_/chanx_left_out[14] sb_5__1_/chanx_left_out[15]
+ sb_5__1_/chanx_left_out[16] sb_5__1_/chanx_left_out[17] sb_5__1_/chanx_left_out[18]
+ sb_5__1_/chanx_left_out[19] sb_5__1_/chanx_left_out[1] sb_5__1_/chanx_left_out[2]
+ sb_5__1_/chanx_left_out[3] sb_5__1_/chanx_left_out[4] sb_5__1_/chanx_left_out[5]
+ sb_5__1_/chanx_left_out[6] sb_5__1_/chanx_left_out[7] sb_5__1_/chanx_left_out[8]
+ sb_5__1_/chanx_left_out[9] sb_5__1_/chanx_left_in[0] sb_5__1_/chanx_left_in[10]
+ sb_5__1_/chanx_left_in[11] sb_5__1_/chanx_left_in[12] sb_5__1_/chanx_left_in[13]
+ sb_5__1_/chanx_left_in[14] sb_5__1_/chanx_left_in[15] sb_5__1_/chanx_left_in[16]
+ sb_5__1_/chanx_left_in[17] sb_5__1_/chanx_left_in[18] sb_5__1_/chanx_left_in[19]
+ sb_5__1_/chanx_left_in[1] sb_5__1_/chanx_left_in[2] sb_5__1_/chanx_left_in[3] sb_5__1_/chanx_left_in[4]
+ sb_5__1_/chanx_left_in[5] sb_5__1_/chanx_left_in[6] sb_5__1_/chanx_left_in[7] sb_5__1_/chanx_left_in[8]
+ sb_5__1_/chanx_left_in[9] cbx_5__1_/clk_1_N_out cbx_5__1_/clk_1_S_out sb_5__1_/clk_1_W_out
+ cbx_5__1_/clk_2_E_out cbx_5__1_/clk_2_W_in cbx_5__1_/clk_2_W_out cbx_5__1_/clk_3_E_out
+ cbx_5__1_/clk_3_W_in cbx_5__1_/clk_3_W_out cbx_5__1_/prog_clk_0_N_in cbx_5__1_/prog_clk_0_W_out
+ cbx_5__1_/prog_clk_1_N_out cbx_5__1_/prog_clk_1_S_out sb_5__1_/prog_clk_1_W_out
+ cbx_5__1_/prog_clk_2_E_out cbx_5__1_/prog_clk_2_W_in cbx_5__1_/prog_clk_2_W_out
+ cbx_5__1_/prog_clk_3_E_out cbx_5__1_/prog_clk_3_W_in cbx_5__1_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_5__6_ sb_5__6_/Test_en_N_out sb_5__6_/Test_en_S_in VGND VPWR sb_5__6_/bottom_left_grid_pin_42_
+ sb_5__6_/bottom_left_grid_pin_43_ sb_5__6_/bottom_left_grid_pin_44_ sb_5__6_/bottom_left_grid_pin_45_
+ sb_5__6_/bottom_left_grid_pin_46_ sb_5__6_/bottom_left_grid_pin_47_ sb_5__6_/bottom_left_grid_pin_48_
+ sb_5__6_/bottom_left_grid_pin_49_ sb_5__6_/ccff_head sb_5__6_/ccff_tail sb_5__6_/chanx_left_in[0]
+ sb_5__6_/chanx_left_in[10] sb_5__6_/chanx_left_in[11] sb_5__6_/chanx_left_in[12]
+ sb_5__6_/chanx_left_in[13] sb_5__6_/chanx_left_in[14] sb_5__6_/chanx_left_in[15]
+ sb_5__6_/chanx_left_in[16] sb_5__6_/chanx_left_in[17] sb_5__6_/chanx_left_in[18]
+ sb_5__6_/chanx_left_in[19] sb_5__6_/chanx_left_in[1] sb_5__6_/chanx_left_in[2] sb_5__6_/chanx_left_in[3]
+ sb_5__6_/chanx_left_in[4] sb_5__6_/chanx_left_in[5] sb_5__6_/chanx_left_in[6] sb_5__6_/chanx_left_in[7]
+ sb_5__6_/chanx_left_in[8] sb_5__6_/chanx_left_in[9] sb_5__6_/chanx_left_out[0] sb_5__6_/chanx_left_out[10]
+ sb_5__6_/chanx_left_out[11] sb_5__6_/chanx_left_out[12] sb_5__6_/chanx_left_out[13]
+ sb_5__6_/chanx_left_out[14] sb_5__6_/chanx_left_out[15] sb_5__6_/chanx_left_out[16]
+ sb_5__6_/chanx_left_out[17] sb_5__6_/chanx_left_out[18] sb_5__6_/chanx_left_out[19]
+ sb_5__6_/chanx_left_out[1] sb_5__6_/chanx_left_out[2] sb_5__6_/chanx_left_out[3]
+ sb_5__6_/chanx_left_out[4] sb_5__6_/chanx_left_out[5] sb_5__6_/chanx_left_out[6]
+ sb_5__6_/chanx_left_out[7] sb_5__6_/chanx_left_out[8] sb_5__6_/chanx_left_out[9]
+ sb_5__6_/chanx_right_in[0] sb_5__6_/chanx_right_in[10] sb_5__6_/chanx_right_in[11]
+ sb_5__6_/chanx_right_in[12] sb_5__6_/chanx_right_in[13] sb_5__6_/chanx_right_in[14]
+ sb_5__6_/chanx_right_in[15] sb_5__6_/chanx_right_in[16] sb_5__6_/chanx_right_in[17]
+ sb_5__6_/chanx_right_in[18] sb_5__6_/chanx_right_in[19] sb_5__6_/chanx_right_in[1]
+ sb_5__6_/chanx_right_in[2] sb_5__6_/chanx_right_in[3] sb_5__6_/chanx_right_in[4]
+ sb_5__6_/chanx_right_in[5] sb_5__6_/chanx_right_in[6] sb_5__6_/chanx_right_in[7]
+ sb_5__6_/chanx_right_in[8] sb_5__6_/chanx_right_in[9] cbx_6__6_/chanx_left_in[0]
+ cbx_6__6_/chanx_left_in[10] cbx_6__6_/chanx_left_in[11] cbx_6__6_/chanx_left_in[12]
+ cbx_6__6_/chanx_left_in[13] cbx_6__6_/chanx_left_in[14] cbx_6__6_/chanx_left_in[15]
+ cbx_6__6_/chanx_left_in[16] cbx_6__6_/chanx_left_in[17] cbx_6__6_/chanx_left_in[18]
+ cbx_6__6_/chanx_left_in[19] cbx_6__6_/chanx_left_in[1] cbx_6__6_/chanx_left_in[2]
+ cbx_6__6_/chanx_left_in[3] cbx_6__6_/chanx_left_in[4] cbx_6__6_/chanx_left_in[5]
+ cbx_6__6_/chanx_left_in[6] cbx_6__6_/chanx_left_in[7] cbx_6__6_/chanx_left_in[8]
+ cbx_6__6_/chanx_left_in[9] cby_5__6_/chany_top_out[0] cby_5__6_/chany_top_out[10]
+ cby_5__6_/chany_top_out[11] cby_5__6_/chany_top_out[12] cby_5__6_/chany_top_out[13]
+ cby_5__6_/chany_top_out[14] cby_5__6_/chany_top_out[15] cby_5__6_/chany_top_out[16]
+ cby_5__6_/chany_top_out[17] cby_5__6_/chany_top_out[18] cby_5__6_/chany_top_out[19]
+ cby_5__6_/chany_top_out[1] cby_5__6_/chany_top_out[2] cby_5__6_/chany_top_out[3]
+ cby_5__6_/chany_top_out[4] cby_5__6_/chany_top_out[5] cby_5__6_/chany_top_out[6]
+ cby_5__6_/chany_top_out[7] cby_5__6_/chany_top_out[8] cby_5__6_/chany_top_out[9]
+ cby_5__6_/chany_top_in[0] cby_5__6_/chany_top_in[10] cby_5__6_/chany_top_in[11]
+ cby_5__6_/chany_top_in[12] cby_5__6_/chany_top_in[13] cby_5__6_/chany_top_in[14]
+ cby_5__6_/chany_top_in[15] cby_5__6_/chany_top_in[16] cby_5__6_/chany_top_in[17]
+ cby_5__6_/chany_top_in[18] cby_5__6_/chany_top_in[19] cby_5__6_/chany_top_in[1]
+ cby_5__6_/chany_top_in[2] cby_5__6_/chany_top_in[3] cby_5__6_/chany_top_in[4] cby_5__6_/chany_top_in[5]
+ cby_5__6_/chany_top_in[6] cby_5__6_/chany_top_in[7] cby_5__6_/chany_top_in[8] cby_5__6_/chany_top_in[9]
+ sb_5__6_/chany_top_in[0] sb_5__6_/chany_top_in[10] sb_5__6_/chany_top_in[11] sb_5__6_/chany_top_in[12]
+ sb_5__6_/chany_top_in[13] sb_5__6_/chany_top_in[14] sb_5__6_/chany_top_in[15] sb_5__6_/chany_top_in[16]
+ sb_5__6_/chany_top_in[17] sb_5__6_/chany_top_in[18] sb_5__6_/chany_top_in[19] sb_5__6_/chany_top_in[1]
+ sb_5__6_/chany_top_in[2] sb_5__6_/chany_top_in[3] sb_5__6_/chany_top_in[4] sb_5__6_/chany_top_in[5]
+ sb_5__6_/chany_top_in[6] sb_5__6_/chany_top_in[7] sb_5__6_/chany_top_in[8] sb_5__6_/chany_top_in[9]
+ sb_5__6_/chany_top_out[0] sb_5__6_/chany_top_out[10] sb_5__6_/chany_top_out[11]
+ sb_5__6_/chany_top_out[12] sb_5__6_/chany_top_out[13] sb_5__6_/chany_top_out[14]
+ sb_5__6_/chany_top_out[15] sb_5__6_/chany_top_out[16] sb_5__6_/chany_top_out[17]
+ sb_5__6_/chany_top_out[18] sb_5__6_/chany_top_out[19] sb_5__6_/chany_top_out[1]
+ sb_5__6_/chany_top_out[2] sb_5__6_/chany_top_out[3] sb_5__6_/chany_top_out[4] sb_5__6_/chany_top_out[5]
+ sb_5__6_/chany_top_out[6] sb_5__6_/chany_top_out[7] sb_5__6_/chany_top_out[8] sb_5__6_/chany_top_out[9]
+ sb_5__6_/clk_1_E_out sb_5__6_/clk_1_N_in sb_5__6_/clk_1_W_out sb_5__6_/clk_2_E_out
+ sb_5__6_/clk_2_N_in sb_5__6_/clk_2_N_out sb_5__6_/clk_2_S_out sb_5__6_/clk_2_W_out
+ sb_5__6_/clk_3_E_out sb_5__6_/clk_3_N_in sb_5__6_/clk_3_N_out sb_5__6_/clk_3_S_out
+ sb_5__6_/clk_3_W_out sb_5__6_/left_bottom_grid_pin_34_ sb_5__6_/left_bottom_grid_pin_35_
+ sb_5__6_/left_bottom_grid_pin_36_ sb_5__6_/left_bottom_grid_pin_37_ sb_5__6_/left_bottom_grid_pin_38_
+ sb_5__6_/left_bottom_grid_pin_39_ sb_5__6_/left_bottom_grid_pin_40_ sb_5__6_/left_bottom_grid_pin_41_
+ sb_5__6_/prog_clk_0_N_in sb_5__6_/prog_clk_1_E_out sb_5__6_/prog_clk_1_N_in sb_5__6_/prog_clk_1_W_out
+ sb_5__6_/prog_clk_2_E_out sb_5__6_/prog_clk_2_N_in sb_5__6_/prog_clk_2_N_out sb_5__6_/prog_clk_2_S_out
+ sb_5__6_/prog_clk_2_W_out sb_5__6_/prog_clk_3_E_out sb_5__6_/prog_clk_3_N_in sb_5__6_/prog_clk_3_N_out
+ sb_5__6_/prog_clk_3_S_out sb_5__6_/prog_clk_3_W_out sb_5__6_/right_bottom_grid_pin_34_
+ sb_5__6_/right_bottom_grid_pin_35_ sb_5__6_/right_bottom_grid_pin_36_ sb_5__6_/right_bottom_grid_pin_37_
+ sb_5__6_/right_bottom_grid_pin_38_ sb_5__6_/right_bottom_grid_pin_39_ sb_5__6_/right_bottom_grid_pin_40_
+ sb_5__6_/right_bottom_grid_pin_41_ sb_5__6_/top_left_grid_pin_42_ sb_5__6_/top_left_grid_pin_43_
+ sb_5__6_/top_left_grid_pin_44_ sb_5__6_/top_left_grid_pin_45_ sb_5__6_/top_left_grid_pin_46_
+ sb_5__6_/top_left_grid_pin_47_ sb_5__6_/top_left_grid_pin_48_ sb_5__6_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_2__3_ sb_2__3_/Test_en_N_out sb_2__3_/Test_en_S_in VGND VPWR sb_2__3_/bottom_left_grid_pin_42_
+ sb_2__3_/bottom_left_grid_pin_43_ sb_2__3_/bottom_left_grid_pin_44_ sb_2__3_/bottom_left_grid_pin_45_
+ sb_2__3_/bottom_left_grid_pin_46_ sb_2__3_/bottom_left_grid_pin_47_ sb_2__3_/bottom_left_grid_pin_48_
+ sb_2__3_/bottom_left_grid_pin_49_ sb_2__3_/ccff_head sb_2__3_/ccff_tail sb_2__3_/chanx_left_in[0]
+ sb_2__3_/chanx_left_in[10] sb_2__3_/chanx_left_in[11] sb_2__3_/chanx_left_in[12]
+ sb_2__3_/chanx_left_in[13] sb_2__3_/chanx_left_in[14] sb_2__3_/chanx_left_in[15]
+ sb_2__3_/chanx_left_in[16] sb_2__3_/chanx_left_in[17] sb_2__3_/chanx_left_in[18]
+ sb_2__3_/chanx_left_in[19] sb_2__3_/chanx_left_in[1] sb_2__3_/chanx_left_in[2] sb_2__3_/chanx_left_in[3]
+ sb_2__3_/chanx_left_in[4] sb_2__3_/chanx_left_in[5] sb_2__3_/chanx_left_in[6] sb_2__3_/chanx_left_in[7]
+ sb_2__3_/chanx_left_in[8] sb_2__3_/chanx_left_in[9] sb_2__3_/chanx_left_out[0] sb_2__3_/chanx_left_out[10]
+ sb_2__3_/chanx_left_out[11] sb_2__3_/chanx_left_out[12] sb_2__3_/chanx_left_out[13]
+ sb_2__3_/chanx_left_out[14] sb_2__3_/chanx_left_out[15] sb_2__3_/chanx_left_out[16]
+ sb_2__3_/chanx_left_out[17] sb_2__3_/chanx_left_out[18] sb_2__3_/chanx_left_out[19]
+ sb_2__3_/chanx_left_out[1] sb_2__3_/chanx_left_out[2] sb_2__3_/chanx_left_out[3]
+ sb_2__3_/chanx_left_out[4] sb_2__3_/chanx_left_out[5] sb_2__3_/chanx_left_out[6]
+ sb_2__3_/chanx_left_out[7] sb_2__3_/chanx_left_out[8] sb_2__3_/chanx_left_out[9]
+ sb_2__3_/chanx_right_in[0] sb_2__3_/chanx_right_in[10] sb_2__3_/chanx_right_in[11]
+ sb_2__3_/chanx_right_in[12] sb_2__3_/chanx_right_in[13] sb_2__3_/chanx_right_in[14]
+ sb_2__3_/chanx_right_in[15] sb_2__3_/chanx_right_in[16] sb_2__3_/chanx_right_in[17]
+ sb_2__3_/chanx_right_in[18] sb_2__3_/chanx_right_in[19] sb_2__3_/chanx_right_in[1]
+ sb_2__3_/chanx_right_in[2] sb_2__3_/chanx_right_in[3] sb_2__3_/chanx_right_in[4]
+ sb_2__3_/chanx_right_in[5] sb_2__3_/chanx_right_in[6] sb_2__3_/chanx_right_in[7]
+ sb_2__3_/chanx_right_in[8] sb_2__3_/chanx_right_in[9] cbx_3__3_/chanx_left_in[0]
+ cbx_3__3_/chanx_left_in[10] cbx_3__3_/chanx_left_in[11] cbx_3__3_/chanx_left_in[12]
+ cbx_3__3_/chanx_left_in[13] cbx_3__3_/chanx_left_in[14] cbx_3__3_/chanx_left_in[15]
+ cbx_3__3_/chanx_left_in[16] cbx_3__3_/chanx_left_in[17] cbx_3__3_/chanx_left_in[18]
+ cbx_3__3_/chanx_left_in[19] cbx_3__3_/chanx_left_in[1] cbx_3__3_/chanx_left_in[2]
+ cbx_3__3_/chanx_left_in[3] cbx_3__3_/chanx_left_in[4] cbx_3__3_/chanx_left_in[5]
+ cbx_3__3_/chanx_left_in[6] cbx_3__3_/chanx_left_in[7] cbx_3__3_/chanx_left_in[8]
+ cbx_3__3_/chanx_left_in[9] cby_2__3_/chany_top_out[0] cby_2__3_/chany_top_out[10]
+ cby_2__3_/chany_top_out[11] cby_2__3_/chany_top_out[12] cby_2__3_/chany_top_out[13]
+ cby_2__3_/chany_top_out[14] cby_2__3_/chany_top_out[15] cby_2__3_/chany_top_out[16]
+ cby_2__3_/chany_top_out[17] cby_2__3_/chany_top_out[18] cby_2__3_/chany_top_out[19]
+ cby_2__3_/chany_top_out[1] cby_2__3_/chany_top_out[2] cby_2__3_/chany_top_out[3]
+ cby_2__3_/chany_top_out[4] cby_2__3_/chany_top_out[5] cby_2__3_/chany_top_out[6]
+ cby_2__3_/chany_top_out[7] cby_2__3_/chany_top_out[8] cby_2__3_/chany_top_out[9]
+ cby_2__3_/chany_top_in[0] cby_2__3_/chany_top_in[10] cby_2__3_/chany_top_in[11]
+ cby_2__3_/chany_top_in[12] cby_2__3_/chany_top_in[13] cby_2__3_/chany_top_in[14]
+ cby_2__3_/chany_top_in[15] cby_2__3_/chany_top_in[16] cby_2__3_/chany_top_in[17]
+ cby_2__3_/chany_top_in[18] cby_2__3_/chany_top_in[19] cby_2__3_/chany_top_in[1]
+ cby_2__3_/chany_top_in[2] cby_2__3_/chany_top_in[3] cby_2__3_/chany_top_in[4] cby_2__3_/chany_top_in[5]
+ cby_2__3_/chany_top_in[6] cby_2__3_/chany_top_in[7] cby_2__3_/chany_top_in[8] cby_2__3_/chany_top_in[9]
+ sb_2__3_/chany_top_in[0] sb_2__3_/chany_top_in[10] sb_2__3_/chany_top_in[11] sb_2__3_/chany_top_in[12]
+ sb_2__3_/chany_top_in[13] sb_2__3_/chany_top_in[14] sb_2__3_/chany_top_in[15] sb_2__3_/chany_top_in[16]
+ sb_2__3_/chany_top_in[17] sb_2__3_/chany_top_in[18] sb_2__3_/chany_top_in[19] sb_2__3_/chany_top_in[1]
+ sb_2__3_/chany_top_in[2] sb_2__3_/chany_top_in[3] sb_2__3_/chany_top_in[4] sb_2__3_/chany_top_in[5]
+ sb_2__3_/chany_top_in[6] sb_2__3_/chany_top_in[7] sb_2__3_/chany_top_in[8] sb_2__3_/chany_top_in[9]
+ sb_2__3_/chany_top_out[0] sb_2__3_/chany_top_out[10] sb_2__3_/chany_top_out[11]
+ sb_2__3_/chany_top_out[12] sb_2__3_/chany_top_out[13] sb_2__3_/chany_top_out[14]
+ sb_2__3_/chany_top_out[15] sb_2__3_/chany_top_out[16] sb_2__3_/chany_top_out[17]
+ sb_2__3_/chany_top_out[18] sb_2__3_/chany_top_out[19] sb_2__3_/chany_top_out[1]
+ sb_2__3_/chany_top_out[2] sb_2__3_/chany_top_out[3] sb_2__3_/chany_top_out[4] sb_2__3_/chany_top_out[5]
+ sb_2__3_/chany_top_out[6] sb_2__3_/chany_top_out[7] sb_2__3_/chany_top_out[8] sb_2__3_/chany_top_out[9]
+ sb_2__3_/clk_1_E_out sb_2__3_/clk_1_N_in sb_2__3_/clk_1_W_out sb_2__3_/clk_2_E_out
+ sb_2__3_/clk_2_N_in sb_2__3_/clk_2_N_out sb_2__3_/clk_2_S_out sb_2__3_/clk_2_W_out
+ sb_2__3_/clk_3_E_out sb_2__3_/clk_3_N_in sb_2__3_/clk_3_N_out sb_2__3_/clk_3_S_out
+ sb_2__3_/clk_3_W_out sb_2__3_/left_bottom_grid_pin_34_ sb_2__3_/left_bottom_grid_pin_35_
+ sb_2__3_/left_bottom_grid_pin_36_ sb_2__3_/left_bottom_grid_pin_37_ sb_2__3_/left_bottom_grid_pin_38_
+ sb_2__3_/left_bottom_grid_pin_39_ sb_2__3_/left_bottom_grid_pin_40_ sb_2__3_/left_bottom_grid_pin_41_
+ sb_2__3_/prog_clk_0_N_in sb_2__3_/prog_clk_1_E_out sb_2__3_/prog_clk_1_N_in sb_2__3_/prog_clk_1_W_out
+ sb_2__3_/prog_clk_2_E_out sb_2__3_/prog_clk_2_N_in sb_2__3_/prog_clk_2_N_out sb_2__3_/prog_clk_2_S_out
+ sb_2__3_/prog_clk_2_W_out sb_2__3_/prog_clk_3_E_out sb_2__3_/prog_clk_3_N_in sb_2__3_/prog_clk_3_N_out
+ sb_2__3_/prog_clk_3_S_out sb_2__3_/prog_clk_3_W_out sb_2__3_/right_bottom_grid_pin_34_
+ sb_2__3_/right_bottom_grid_pin_35_ sb_2__3_/right_bottom_grid_pin_36_ sb_2__3_/right_bottom_grid_pin_37_
+ sb_2__3_/right_bottom_grid_pin_38_ sb_2__3_/right_bottom_grid_pin_39_ sb_2__3_/right_bottom_grid_pin_40_
+ sb_2__3_/right_bottom_grid_pin_41_ sb_2__3_/top_left_grid_pin_42_ sb_2__3_/top_left_grid_pin_43_
+ sb_2__3_/top_left_grid_pin_44_ sb_2__3_/top_left_grid_pin_45_ sb_2__3_/top_left_grid_pin_46_
+ sb_2__3_/top_left_grid_pin_47_ sb_2__3_/top_left_grid_pin_48_ sb_2__3_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_8__2_ IO_ISOL_N VGND VPWR cby_8__2_/ccff_head sb_8__1_/ccff_head sb_8__1_/chany_top_out[0]
+ sb_8__1_/chany_top_out[10] sb_8__1_/chany_top_out[11] sb_8__1_/chany_top_out[12]
+ sb_8__1_/chany_top_out[13] sb_8__1_/chany_top_out[14] sb_8__1_/chany_top_out[15]
+ sb_8__1_/chany_top_out[16] sb_8__1_/chany_top_out[17] sb_8__1_/chany_top_out[18]
+ sb_8__1_/chany_top_out[19] sb_8__1_/chany_top_out[1] sb_8__1_/chany_top_out[2] sb_8__1_/chany_top_out[3]
+ sb_8__1_/chany_top_out[4] sb_8__1_/chany_top_out[5] sb_8__1_/chany_top_out[6] sb_8__1_/chany_top_out[7]
+ sb_8__1_/chany_top_out[8] sb_8__1_/chany_top_out[9] sb_8__1_/chany_top_in[0] sb_8__1_/chany_top_in[10]
+ sb_8__1_/chany_top_in[11] sb_8__1_/chany_top_in[12] sb_8__1_/chany_top_in[13] sb_8__1_/chany_top_in[14]
+ sb_8__1_/chany_top_in[15] sb_8__1_/chany_top_in[16] sb_8__1_/chany_top_in[17] sb_8__1_/chany_top_in[18]
+ sb_8__1_/chany_top_in[19] sb_8__1_/chany_top_in[1] sb_8__1_/chany_top_in[2] sb_8__1_/chany_top_in[3]
+ sb_8__1_/chany_top_in[4] sb_8__1_/chany_top_in[5] sb_8__1_/chany_top_in[6] sb_8__1_/chany_top_in[7]
+ sb_8__1_/chany_top_in[8] sb_8__1_/chany_top_in[9] cby_8__2_/chany_top_in[0] cby_8__2_/chany_top_in[10]
+ cby_8__2_/chany_top_in[11] cby_8__2_/chany_top_in[12] cby_8__2_/chany_top_in[13]
+ cby_8__2_/chany_top_in[14] cby_8__2_/chany_top_in[15] cby_8__2_/chany_top_in[16]
+ cby_8__2_/chany_top_in[17] cby_8__2_/chany_top_in[18] cby_8__2_/chany_top_in[19]
+ cby_8__2_/chany_top_in[1] cby_8__2_/chany_top_in[2] cby_8__2_/chany_top_in[3] cby_8__2_/chany_top_in[4]
+ cby_8__2_/chany_top_in[5] cby_8__2_/chany_top_in[6] cby_8__2_/chany_top_in[7] cby_8__2_/chany_top_in[8]
+ cby_8__2_/chany_top_in[9] cby_8__2_/chany_top_out[0] cby_8__2_/chany_top_out[10]
+ cby_8__2_/chany_top_out[11] cby_8__2_/chany_top_out[12] cby_8__2_/chany_top_out[13]
+ cby_8__2_/chany_top_out[14] cby_8__2_/chany_top_out[15] cby_8__2_/chany_top_out[16]
+ cby_8__2_/chany_top_out[17] cby_8__2_/chany_top_out[18] cby_8__2_/chany_top_out[19]
+ cby_8__2_/chany_top_out[1] cby_8__2_/chany_top_out[2] cby_8__2_/chany_top_out[3]
+ cby_8__2_/chany_top_out[4] cby_8__2_/chany_top_out[5] cby_8__2_/chany_top_out[6]
+ cby_8__2_/chany_top_out[7] cby_8__2_/chany_top_out[8] cby_8__2_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
+ cby_8__2_/left_grid_pin_16_ cby_8__2_/left_grid_pin_17_ cby_8__2_/left_grid_pin_18_
+ cby_8__2_/left_grid_pin_19_ cby_8__2_/left_grid_pin_20_ cby_8__2_/left_grid_pin_21_
+ cby_8__2_/left_grid_pin_22_ cby_8__2_/left_grid_pin_23_ cby_8__2_/left_grid_pin_24_
+ cby_8__2_/left_grid_pin_25_ cby_8__2_/left_grid_pin_26_ cby_8__2_/left_grid_pin_27_
+ cby_8__2_/left_grid_pin_28_ cby_8__2_/left_grid_pin_29_ cby_8__2_/left_grid_pin_30_
+ cby_8__2_/left_grid_pin_31_ cby_8__2_/right_grid_pin_0_ sb_8__1_/top_right_grid_pin_1_
+ sb_8__2_/bottom_right_grid_pin_1_ cby_8__2_/prog_clk_0_N_out sb_8__1_/prog_clk_0_N_in
+ cby_8__2_/prog_clk_0_W_in cby_8__2_/right_grid_pin_0_ cby_2__1_
Xcby_1__7_ cby_1__7_/Test_en_W_in cby_1__7_/Test_en_E_out cby_1__7_/Test_en_N_out
+ cby_1__7_/Test_en_W_in cby_1__7_/Test_en_W_in cby_1__7_/Test_en_W_out VGND VPWR
+ cby_1__7_/ccff_head cby_1__7_/ccff_tail sb_1__6_/chany_top_out[0] sb_1__6_/chany_top_out[10]
+ sb_1__6_/chany_top_out[11] sb_1__6_/chany_top_out[12] sb_1__6_/chany_top_out[13]
+ sb_1__6_/chany_top_out[14] sb_1__6_/chany_top_out[15] sb_1__6_/chany_top_out[16]
+ sb_1__6_/chany_top_out[17] sb_1__6_/chany_top_out[18] sb_1__6_/chany_top_out[19]
+ sb_1__6_/chany_top_out[1] sb_1__6_/chany_top_out[2] sb_1__6_/chany_top_out[3] sb_1__6_/chany_top_out[4]
+ sb_1__6_/chany_top_out[5] sb_1__6_/chany_top_out[6] sb_1__6_/chany_top_out[7] sb_1__6_/chany_top_out[8]
+ sb_1__6_/chany_top_out[9] sb_1__6_/chany_top_in[0] sb_1__6_/chany_top_in[10] sb_1__6_/chany_top_in[11]
+ sb_1__6_/chany_top_in[12] sb_1__6_/chany_top_in[13] sb_1__6_/chany_top_in[14] sb_1__6_/chany_top_in[15]
+ sb_1__6_/chany_top_in[16] sb_1__6_/chany_top_in[17] sb_1__6_/chany_top_in[18] sb_1__6_/chany_top_in[19]
+ sb_1__6_/chany_top_in[1] sb_1__6_/chany_top_in[2] sb_1__6_/chany_top_in[3] sb_1__6_/chany_top_in[4]
+ sb_1__6_/chany_top_in[5] sb_1__6_/chany_top_in[6] sb_1__6_/chany_top_in[7] sb_1__6_/chany_top_in[8]
+ sb_1__6_/chany_top_in[9] cby_1__7_/chany_top_in[0] cby_1__7_/chany_top_in[10] cby_1__7_/chany_top_in[11]
+ cby_1__7_/chany_top_in[12] cby_1__7_/chany_top_in[13] cby_1__7_/chany_top_in[14]
+ cby_1__7_/chany_top_in[15] cby_1__7_/chany_top_in[16] cby_1__7_/chany_top_in[17]
+ cby_1__7_/chany_top_in[18] cby_1__7_/chany_top_in[19] cby_1__7_/chany_top_in[1]
+ cby_1__7_/chany_top_in[2] cby_1__7_/chany_top_in[3] cby_1__7_/chany_top_in[4] cby_1__7_/chany_top_in[5]
+ cby_1__7_/chany_top_in[6] cby_1__7_/chany_top_in[7] cby_1__7_/chany_top_in[8] cby_1__7_/chany_top_in[9]
+ cby_1__7_/chany_top_out[0] cby_1__7_/chany_top_out[10] cby_1__7_/chany_top_out[11]
+ cby_1__7_/chany_top_out[12] cby_1__7_/chany_top_out[13] cby_1__7_/chany_top_out[14]
+ cby_1__7_/chany_top_out[15] cby_1__7_/chany_top_out[16] cby_1__7_/chany_top_out[17]
+ cby_1__7_/chany_top_out[18] cby_1__7_/chany_top_out[19] cby_1__7_/chany_top_out[1]
+ cby_1__7_/chany_top_out[2] cby_1__7_/chany_top_out[3] cby_1__7_/chany_top_out[4]
+ cby_1__7_/chany_top_out[5] cby_1__7_/chany_top_out[6] cby_1__7_/chany_top_out[7]
+ cby_1__7_/chany_top_out[8] cby_1__7_/chany_top_out[9] sb_1__7_/clk_1_N_in sb_1__6_/clk_2_N_out
+ cby_1__7_/clk_2_S_out cby_1__7_/clk_3_N_out cby_1__7_/clk_3_S_in cby_1__7_/clk_3_S_out
+ cby_1__7_/left_grid_pin_16_ cby_1__7_/left_grid_pin_17_ cby_1__7_/left_grid_pin_18_
+ cby_1__7_/left_grid_pin_19_ cby_1__7_/left_grid_pin_20_ cby_1__7_/left_grid_pin_21_
+ cby_1__7_/left_grid_pin_22_ cby_1__7_/left_grid_pin_23_ cby_1__7_/left_grid_pin_24_
+ cby_1__7_/left_grid_pin_25_ cby_1__7_/left_grid_pin_26_ cby_1__7_/left_grid_pin_27_
+ cby_1__7_/left_grid_pin_28_ cby_1__7_/left_grid_pin_29_ cby_1__7_/left_grid_pin_30_
+ cby_1__7_/left_grid_pin_31_ cby_1__7_/prog_clk_0_N_out sb_1__6_/prog_clk_0_N_in
+ cby_1__7_/prog_clk_0_W_in sb_1__7_/prog_clk_1_N_in sb_1__6_/prog_clk_2_N_out cby_1__7_/prog_clk_2_S_out
+ cby_1__7_/prog_clk_3_N_out cby_1__7_/prog_clk_3_S_in cby_1__7_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_8__3_ cbx_8__3_/REGIN_FEEDTHROUGH cbx_8__3_/REGOUT_FEEDTHROUGH cbx_8__3_/SC_IN_BOT
+ cbx_8__3_/SC_IN_TOP cbx_8__3_/SC_OUT_BOT cbx_8__3_/SC_OUT_TOP VGND VPWR cbx_8__3_/bottom_grid_pin_0_
+ cbx_8__3_/bottom_grid_pin_10_ cbx_8__3_/bottom_grid_pin_11_ cbx_8__3_/bottom_grid_pin_12_
+ cbx_8__3_/bottom_grid_pin_13_ cbx_8__3_/bottom_grid_pin_14_ cbx_8__3_/bottom_grid_pin_15_
+ cbx_8__3_/bottom_grid_pin_1_ cbx_8__3_/bottom_grid_pin_2_ cbx_8__3_/bottom_grid_pin_3_
+ cbx_8__3_/bottom_grid_pin_4_ cbx_8__3_/bottom_grid_pin_5_ cbx_8__3_/bottom_grid_pin_6_
+ cbx_8__3_/bottom_grid_pin_7_ cbx_8__3_/bottom_grid_pin_8_ cbx_8__3_/bottom_grid_pin_9_
+ sb_8__3_/ccff_tail sb_7__3_/ccff_head cbx_8__3_/chanx_left_in[0] cbx_8__3_/chanx_left_in[10]
+ cbx_8__3_/chanx_left_in[11] cbx_8__3_/chanx_left_in[12] cbx_8__3_/chanx_left_in[13]
+ cbx_8__3_/chanx_left_in[14] cbx_8__3_/chanx_left_in[15] cbx_8__3_/chanx_left_in[16]
+ cbx_8__3_/chanx_left_in[17] cbx_8__3_/chanx_left_in[18] cbx_8__3_/chanx_left_in[19]
+ cbx_8__3_/chanx_left_in[1] cbx_8__3_/chanx_left_in[2] cbx_8__3_/chanx_left_in[3]
+ cbx_8__3_/chanx_left_in[4] cbx_8__3_/chanx_left_in[5] cbx_8__3_/chanx_left_in[6]
+ cbx_8__3_/chanx_left_in[7] cbx_8__3_/chanx_left_in[8] cbx_8__3_/chanx_left_in[9]
+ sb_7__3_/chanx_right_in[0] sb_7__3_/chanx_right_in[10] sb_7__3_/chanx_right_in[11]
+ sb_7__3_/chanx_right_in[12] sb_7__3_/chanx_right_in[13] sb_7__3_/chanx_right_in[14]
+ sb_7__3_/chanx_right_in[15] sb_7__3_/chanx_right_in[16] sb_7__3_/chanx_right_in[17]
+ sb_7__3_/chanx_right_in[18] sb_7__3_/chanx_right_in[19] sb_7__3_/chanx_right_in[1]
+ sb_7__3_/chanx_right_in[2] sb_7__3_/chanx_right_in[3] sb_7__3_/chanx_right_in[4]
+ sb_7__3_/chanx_right_in[5] sb_7__3_/chanx_right_in[6] sb_7__3_/chanx_right_in[7]
+ sb_7__3_/chanx_right_in[8] sb_7__3_/chanx_right_in[9] sb_8__3_/chanx_left_out[0]
+ sb_8__3_/chanx_left_out[10] sb_8__3_/chanx_left_out[11] sb_8__3_/chanx_left_out[12]
+ sb_8__3_/chanx_left_out[13] sb_8__3_/chanx_left_out[14] sb_8__3_/chanx_left_out[15]
+ sb_8__3_/chanx_left_out[16] sb_8__3_/chanx_left_out[17] sb_8__3_/chanx_left_out[18]
+ sb_8__3_/chanx_left_out[19] sb_8__3_/chanx_left_out[1] sb_8__3_/chanx_left_out[2]
+ sb_8__3_/chanx_left_out[3] sb_8__3_/chanx_left_out[4] sb_8__3_/chanx_left_out[5]
+ sb_8__3_/chanx_left_out[6] sb_8__3_/chanx_left_out[7] sb_8__3_/chanx_left_out[8]
+ sb_8__3_/chanx_left_out[9] sb_8__3_/chanx_left_in[0] sb_8__3_/chanx_left_in[10]
+ sb_8__3_/chanx_left_in[11] sb_8__3_/chanx_left_in[12] sb_8__3_/chanx_left_in[13]
+ sb_8__3_/chanx_left_in[14] sb_8__3_/chanx_left_in[15] sb_8__3_/chanx_left_in[16]
+ sb_8__3_/chanx_left_in[17] sb_8__3_/chanx_left_in[18] sb_8__3_/chanx_left_in[19]
+ sb_8__3_/chanx_left_in[1] sb_8__3_/chanx_left_in[2] sb_8__3_/chanx_left_in[3] sb_8__3_/chanx_left_in[4]
+ sb_8__3_/chanx_left_in[5] sb_8__3_/chanx_left_in[6] sb_8__3_/chanx_left_in[7] sb_8__3_/chanx_left_in[8]
+ sb_8__3_/chanx_left_in[9] cbx_8__3_/clk_1_N_out cbx_8__3_/clk_1_S_out sb_7__3_/clk_1_E_out
+ cbx_8__3_/clk_2_E_out cbx_8__3_/clk_2_W_in cbx_8__3_/clk_2_W_out cbx_8__3_/clk_3_E_out
+ cbx_8__3_/clk_3_W_in cbx_8__3_/clk_3_W_out cbx_8__3_/prog_clk_0_N_in cbx_8__3_/prog_clk_0_W_out
+ cbx_8__3_/prog_clk_1_N_out cbx_8__3_/prog_clk_1_S_out sb_7__3_/prog_clk_1_E_out
+ cbx_8__3_/prog_clk_2_E_out cbx_8__3_/prog_clk_2_W_in cbx_8__3_/prog_clk_2_W_out
+ cbx_8__3_/prog_clk_3_E_out cbx_8__3_/prog_clk_3_W_in cbx_8__3_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_7__3_ cbx_7__3_/SC_OUT_BOT cbx_7__2_/SC_IN_TOP grid_clb_7__3_/SC_OUT_TOP
+ cby_6__3_/Test_en_E_out cby_7__3_/Test_en_W_in cby_6__3_/Test_en_E_out grid_clb_7__3_/Test_en_W_out
+ VGND VPWR cbx_7__2_/REGIN_FEEDTHROUGH grid_clb_7__3_/bottom_width_0_height_0__pin_51_
+ cby_6__3_/ccff_tail cby_7__3_/ccff_head cbx_7__3_/clk_1_S_out cbx_7__3_/clk_1_S_out
+ cby_7__3_/prog_clk_0_W_in cbx_7__3_/prog_clk_1_S_out grid_clb_7__3_/prog_clk_0_N_out
+ cbx_7__3_/prog_clk_1_S_out cbx_7__2_/prog_clk_0_N_in grid_clb_7__3_/prog_clk_0_W_out
+ cby_7__3_/left_grid_pin_16_ cby_7__3_/left_grid_pin_17_ cby_7__3_/left_grid_pin_18_
+ cby_7__3_/left_grid_pin_19_ cby_7__3_/left_grid_pin_20_ cby_7__3_/left_grid_pin_21_
+ cby_7__3_/left_grid_pin_22_ cby_7__3_/left_grid_pin_23_ cby_7__3_/left_grid_pin_24_
+ cby_7__3_/left_grid_pin_25_ cby_7__3_/left_grid_pin_26_ cby_7__3_/left_grid_pin_27_
+ cby_7__3_/left_grid_pin_28_ cby_7__3_/left_grid_pin_29_ cby_7__3_/left_grid_pin_30_
+ cby_7__3_/left_grid_pin_31_ sb_7__2_/top_left_grid_pin_42_ sb_7__3_/bottom_left_grid_pin_42_
+ sb_7__2_/top_left_grid_pin_43_ sb_7__3_/bottom_left_grid_pin_43_ sb_7__2_/top_left_grid_pin_44_
+ sb_7__3_/bottom_left_grid_pin_44_ sb_7__2_/top_left_grid_pin_45_ sb_7__3_/bottom_left_grid_pin_45_
+ sb_7__2_/top_left_grid_pin_46_ sb_7__3_/bottom_left_grid_pin_46_ sb_7__2_/top_left_grid_pin_47_
+ sb_7__3_/bottom_left_grid_pin_47_ sb_7__2_/top_left_grid_pin_48_ sb_7__3_/bottom_left_grid_pin_48_
+ sb_7__2_/top_left_grid_pin_49_ sb_7__3_/bottom_left_grid_pin_49_ cbx_7__3_/bottom_grid_pin_0_
+ cbx_7__3_/bottom_grid_pin_10_ cbx_7__3_/bottom_grid_pin_11_ cbx_7__3_/bottom_grid_pin_12_
+ cbx_7__3_/bottom_grid_pin_13_ cbx_7__3_/bottom_grid_pin_14_ cbx_7__3_/bottom_grid_pin_15_
+ cbx_7__3_/bottom_grid_pin_1_ cbx_7__3_/bottom_grid_pin_2_ cbx_7__3_/REGOUT_FEEDTHROUGH
+ grid_clb_7__3_/top_width_0_height_0__pin_33_ sb_7__3_/left_bottom_grid_pin_34_ sb_6__3_/right_bottom_grid_pin_34_
+ sb_7__3_/left_bottom_grid_pin_35_ sb_6__3_/right_bottom_grid_pin_35_ sb_7__3_/left_bottom_grid_pin_36_
+ sb_6__3_/right_bottom_grid_pin_36_ sb_7__3_/left_bottom_grid_pin_37_ sb_6__3_/right_bottom_grid_pin_37_
+ sb_7__3_/left_bottom_grid_pin_38_ sb_6__3_/right_bottom_grid_pin_38_ sb_7__3_/left_bottom_grid_pin_39_
+ sb_6__3_/right_bottom_grid_pin_39_ cbx_7__3_/bottom_grid_pin_3_ sb_7__3_/left_bottom_grid_pin_40_
+ sb_6__3_/right_bottom_grid_pin_40_ sb_7__3_/left_bottom_grid_pin_41_ sb_6__3_/right_bottom_grid_pin_41_
+ cbx_7__3_/bottom_grid_pin_4_ cbx_7__3_/bottom_grid_pin_5_ cbx_7__3_/bottom_grid_pin_6_
+ cbx_7__3_/bottom_grid_pin_7_ cbx_7__3_/bottom_grid_pin_8_ cbx_7__3_/bottom_grid_pin_9_
+ grid_clb
Xcbx_5__0_ IO_ISOL_N cbx_5__0_/SC_IN_BOT cbx_5__0_/SC_IN_TOP sb_5__0_/SC_IN_TOP cbx_5__0_/SC_OUT_TOP
+ VGND VPWR cbx_5__0_/bottom_grid_pin_0_ cbx_5__0_/bottom_grid_pin_10_ cbx_5__0_/bottom_grid_pin_12_
+ cbx_5__0_/bottom_grid_pin_14_ cbx_5__0_/bottom_grid_pin_16_ cbx_5__0_/bottom_grid_pin_2_
+ cbx_5__0_/bottom_grid_pin_4_ cbx_5__0_/bottom_grid_pin_6_ cbx_5__0_/bottom_grid_pin_8_
+ sb_5__0_/ccff_tail sb_4__0_/ccff_head cbx_5__0_/chanx_left_in[0] cbx_5__0_/chanx_left_in[10]
+ cbx_5__0_/chanx_left_in[11] cbx_5__0_/chanx_left_in[12] cbx_5__0_/chanx_left_in[13]
+ cbx_5__0_/chanx_left_in[14] cbx_5__0_/chanx_left_in[15] cbx_5__0_/chanx_left_in[16]
+ cbx_5__0_/chanx_left_in[17] cbx_5__0_/chanx_left_in[18] cbx_5__0_/chanx_left_in[19]
+ cbx_5__0_/chanx_left_in[1] cbx_5__0_/chanx_left_in[2] cbx_5__0_/chanx_left_in[3]
+ cbx_5__0_/chanx_left_in[4] cbx_5__0_/chanx_left_in[5] cbx_5__0_/chanx_left_in[6]
+ cbx_5__0_/chanx_left_in[7] cbx_5__0_/chanx_left_in[8] cbx_5__0_/chanx_left_in[9]
+ sb_4__0_/chanx_right_in[0] sb_4__0_/chanx_right_in[10] sb_4__0_/chanx_right_in[11]
+ sb_4__0_/chanx_right_in[12] sb_4__0_/chanx_right_in[13] sb_4__0_/chanx_right_in[14]
+ sb_4__0_/chanx_right_in[15] sb_4__0_/chanx_right_in[16] sb_4__0_/chanx_right_in[17]
+ sb_4__0_/chanx_right_in[18] sb_4__0_/chanx_right_in[19] sb_4__0_/chanx_right_in[1]
+ sb_4__0_/chanx_right_in[2] sb_4__0_/chanx_right_in[3] sb_4__0_/chanx_right_in[4]
+ sb_4__0_/chanx_right_in[5] sb_4__0_/chanx_right_in[6] sb_4__0_/chanx_right_in[7]
+ sb_4__0_/chanx_right_in[8] sb_4__0_/chanx_right_in[9] sb_5__0_/chanx_left_out[0]
+ sb_5__0_/chanx_left_out[10] sb_5__0_/chanx_left_out[11] sb_5__0_/chanx_left_out[12]
+ sb_5__0_/chanx_left_out[13] sb_5__0_/chanx_left_out[14] sb_5__0_/chanx_left_out[15]
+ sb_5__0_/chanx_left_out[16] sb_5__0_/chanx_left_out[17] sb_5__0_/chanx_left_out[18]
+ sb_5__0_/chanx_left_out[19] sb_5__0_/chanx_left_out[1] sb_5__0_/chanx_left_out[2]
+ sb_5__0_/chanx_left_out[3] sb_5__0_/chanx_left_out[4] sb_5__0_/chanx_left_out[5]
+ sb_5__0_/chanx_left_out[6] sb_5__0_/chanx_left_out[7] sb_5__0_/chanx_left_out[8]
+ sb_5__0_/chanx_left_out[9] sb_5__0_/chanx_left_in[0] sb_5__0_/chanx_left_in[10]
+ sb_5__0_/chanx_left_in[11] sb_5__0_/chanx_left_in[12] sb_5__0_/chanx_left_in[13]
+ sb_5__0_/chanx_left_in[14] sb_5__0_/chanx_left_in[15] sb_5__0_/chanx_left_in[16]
+ sb_5__0_/chanx_left_in[17] sb_5__0_/chanx_left_in[18] sb_5__0_/chanx_left_in[19]
+ sb_5__0_/chanx_left_in[1] sb_5__0_/chanx_left_in[2] sb_5__0_/chanx_left_in[3] sb_5__0_/chanx_left_in[4]
+ sb_5__0_/chanx_left_in[5] sb_5__0_/chanx_left_in[6] sb_5__0_/chanx_left_in[7] sb_5__0_/chanx_left_in[8]
+ sb_5__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51] cbx_5__0_/prog_clk_0_N_in cbx_5__0_/prog_clk_0_W_out
+ cbx_5__0_/bottom_grid_pin_0_ cbx_5__0_/bottom_grid_pin_10_ sb_5__0_/left_bottom_grid_pin_11_
+ sb_4__0_/right_bottom_grid_pin_11_ cbx_5__0_/bottom_grid_pin_12_ sb_5__0_/left_bottom_grid_pin_13_
+ sb_4__0_/right_bottom_grid_pin_13_ cbx_5__0_/bottom_grid_pin_14_ sb_5__0_/left_bottom_grid_pin_15_
+ sb_4__0_/right_bottom_grid_pin_15_ cbx_5__0_/bottom_grid_pin_16_ sb_5__0_/left_bottom_grid_pin_17_
+ sb_4__0_/right_bottom_grid_pin_17_ sb_5__0_/left_bottom_grid_pin_1_ sb_4__0_/right_bottom_grid_pin_1_
+ cbx_5__0_/bottom_grid_pin_2_ sb_5__0_/left_bottom_grid_pin_3_ sb_4__0_/right_bottom_grid_pin_3_
+ cbx_5__0_/bottom_grid_pin_4_ sb_5__0_/left_bottom_grid_pin_5_ sb_4__0_/right_bottom_grid_pin_5_
+ cbx_5__0_/bottom_grid_pin_6_ sb_5__0_/left_bottom_grid_pin_7_ sb_4__0_/right_bottom_grid_pin_7_
+ cbx_5__0_/bottom_grid_pin_8_ sb_5__0_/left_bottom_grid_pin_9_ sb_4__0_/right_bottom_grid_pin_9_
+ cbx_1__0_
Xsb_8__8_ sb_8__8_/SC_IN_BOT sc_tail VGND VPWR sb_8__8_/bottom_left_grid_pin_42_ sb_8__8_/bottom_left_grid_pin_43_
+ sb_8__8_/bottom_left_grid_pin_44_ sb_8__8_/bottom_left_grid_pin_45_ sb_8__8_/bottom_left_grid_pin_46_
+ sb_8__8_/bottom_left_grid_pin_47_ sb_8__8_/bottom_left_grid_pin_48_ sb_8__8_/bottom_left_grid_pin_49_
+ sb_8__8_/bottom_right_grid_pin_1_ ccff_head sb_8__8_/ccff_tail sb_8__8_/chanx_left_in[0]
+ sb_8__8_/chanx_left_in[10] sb_8__8_/chanx_left_in[11] sb_8__8_/chanx_left_in[12]
+ sb_8__8_/chanx_left_in[13] sb_8__8_/chanx_left_in[14] sb_8__8_/chanx_left_in[15]
+ sb_8__8_/chanx_left_in[16] sb_8__8_/chanx_left_in[17] sb_8__8_/chanx_left_in[18]
+ sb_8__8_/chanx_left_in[19] sb_8__8_/chanx_left_in[1] sb_8__8_/chanx_left_in[2] sb_8__8_/chanx_left_in[3]
+ sb_8__8_/chanx_left_in[4] sb_8__8_/chanx_left_in[5] sb_8__8_/chanx_left_in[6] sb_8__8_/chanx_left_in[7]
+ sb_8__8_/chanx_left_in[8] sb_8__8_/chanx_left_in[9] sb_8__8_/chanx_left_out[0] sb_8__8_/chanx_left_out[10]
+ sb_8__8_/chanx_left_out[11] sb_8__8_/chanx_left_out[12] sb_8__8_/chanx_left_out[13]
+ sb_8__8_/chanx_left_out[14] sb_8__8_/chanx_left_out[15] sb_8__8_/chanx_left_out[16]
+ sb_8__8_/chanx_left_out[17] sb_8__8_/chanx_left_out[18] sb_8__8_/chanx_left_out[19]
+ sb_8__8_/chanx_left_out[1] sb_8__8_/chanx_left_out[2] sb_8__8_/chanx_left_out[3]
+ sb_8__8_/chanx_left_out[4] sb_8__8_/chanx_left_out[5] sb_8__8_/chanx_left_out[6]
+ sb_8__8_/chanx_left_out[7] sb_8__8_/chanx_left_out[8] sb_8__8_/chanx_left_out[9]
+ cby_8__8_/chany_top_out[0] cby_8__8_/chany_top_out[10] cby_8__8_/chany_top_out[11]
+ cby_8__8_/chany_top_out[12] cby_8__8_/chany_top_out[13] cby_8__8_/chany_top_out[14]
+ cby_8__8_/chany_top_out[15] cby_8__8_/chany_top_out[16] cby_8__8_/chany_top_out[17]
+ cby_8__8_/chany_top_out[18] cby_8__8_/chany_top_out[19] cby_8__8_/chany_top_out[1]
+ cby_8__8_/chany_top_out[2] cby_8__8_/chany_top_out[3] cby_8__8_/chany_top_out[4]
+ cby_8__8_/chany_top_out[5] cby_8__8_/chany_top_out[6] cby_8__8_/chany_top_out[7]
+ cby_8__8_/chany_top_out[8] cby_8__8_/chany_top_out[9] cby_8__8_/chany_top_in[0]
+ cby_8__8_/chany_top_in[10] cby_8__8_/chany_top_in[11] cby_8__8_/chany_top_in[12]
+ cby_8__8_/chany_top_in[13] cby_8__8_/chany_top_in[14] cby_8__8_/chany_top_in[15]
+ cby_8__8_/chany_top_in[16] cby_8__8_/chany_top_in[17] cby_8__8_/chany_top_in[18]
+ cby_8__8_/chany_top_in[19] cby_8__8_/chany_top_in[1] cby_8__8_/chany_top_in[2] cby_8__8_/chany_top_in[3]
+ cby_8__8_/chany_top_in[4] cby_8__8_/chany_top_in[5] cby_8__8_/chany_top_in[6] cby_8__8_/chany_top_in[7]
+ cby_8__8_/chany_top_in[8] cby_8__8_/chany_top_in[9] sb_8__8_/left_bottom_grid_pin_34_
+ sb_8__8_/left_bottom_grid_pin_35_ sb_8__8_/left_bottom_grid_pin_36_ sb_8__8_/left_bottom_grid_pin_37_
+ sb_8__8_/left_bottom_grid_pin_38_ sb_8__8_/left_bottom_grid_pin_39_ sb_8__8_/left_bottom_grid_pin_40_
+ sb_8__8_/left_bottom_grid_pin_41_ sb_8__8_/left_top_grid_pin_1_ sb_8__8_/prog_clk_0_S_in
+ sb_2__2_
Xcbx_1__8_ IO_ISOL_N cbx_1__8_/SC_IN_BOT sb_0__8_/SC_OUT_BOT cbx_1__8_/SC_OUT_BOT
+ cbx_1__8_/SC_OUT_TOP VGND VPWR cbx_1__8_/bottom_grid_pin_0_ cbx_1__8_/bottom_grid_pin_10_
+ cbx_1__8_/bottom_grid_pin_11_ cbx_1__8_/bottom_grid_pin_12_ cbx_1__8_/bottom_grid_pin_13_
+ cbx_1__8_/bottom_grid_pin_14_ cbx_1__8_/bottom_grid_pin_15_ cbx_1__8_/bottom_grid_pin_1_
+ cbx_1__8_/bottom_grid_pin_2_ cbx_1__8_/bottom_grid_pin_3_ cbx_1__8_/bottom_grid_pin_4_
+ cbx_1__8_/bottom_grid_pin_5_ cbx_1__8_/bottom_grid_pin_6_ cbx_1__8_/bottom_grid_pin_7_
+ cbx_1__8_/bottom_grid_pin_8_ cbx_1__8_/bottom_grid_pin_9_ cbx_1__8_/top_grid_pin_0_
+ sb_1__8_/left_top_grid_pin_1_ sb_0__8_/right_top_grid_pin_1_ sb_1__8_/ccff_tail
+ sb_0__8_/ccff_head cbx_1__8_/chanx_left_in[0] cbx_1__8_/chanx_left_in[10] cbx_1__8_/chanx_left_in[11]
+ cbx_1__8_/chanx_left_in[12] cbx_1__8_/chanx_left_in[13] cbx_1__8_/chanx_left_in[14]
+ cbx_1__8_/chanx_left_in[15] cbx_1__8_/chanx_left_in[16] cbx_1__8_/chanx_left_in[17]
+ cbx_1__8_/chanx_left_in[18] cbx_1__8_/chanx_left_in[19] cbx_1__8_/chanx_left_in[1]
+ cbx_1__8_/chanx_left_in[2] cbx_1__8_/chanx_left_in[3] cbx_1__8_/chanx_left_in[4]
+ cbx_1__8_/chanx_left_in[5] cbx_1__8_/chanx_left_in[6] cbx_1__8_/chanx_left_in[7]
+ cbx_1__8_/chanx_left_in[8] cbx_1__8_/chanx_left_in[9] sb_0__8_/chanx_right_in[0]
+ sb_0__8_/chanx_right_in[10] sb_0__8_/chanx_right_in[11] sb_0__8_/chanx_right_in[12]
+ sb_0__8_/chanx_right_in[13] sb_0__8_/chanx_right_in[14] sb_0__8_/chanx_right_in[15]
+ sb_0__8_/chanx_right_in[16] sb_0__8_/chanx_right_in[17] sb_0__8_/chanx_right_in[18]
+ sb_0__8_/chanx_right_in[19] sb_0__8_/chanx_right_in[1] sb_0__8_/chanx_right_in[2]
+ sb_0__8_/chanx_right_in[3] sb_0__8_/chanx_right_in[4] sb_0__8_/chanx_right_in[5]
+ sb_0__8_/chanx_right_in[6] sb_0__8_/chanx_right_in[7] sb_0__8_/chanx_right_in[8]
+ sb_0__8_/chanx_right_in[9] sb_1__8_/chanx_left_out[0] sb_1__8_/chanx_left_out[10]
+ sb_1__8_/chanx_left_out[11] sb_1__8_/chanx_left_out[12] sb_1__8_/chanx_left_out[13]
+ sb_1__8_/chanx_left_out[14] sb_1__8_/chanx_left_out[15] sb_1__8_/chanx_left_out[16]
+ sb_1__8_/chanx_left_out[17] sb_1__8_/chanx_left_out[18] sb_1__8_/chanx_left_out[19]
+ sb_1__8_/chanx_left_out[1] sb_1__8_/chanx_left_out[2] sb_1__8_/chanx_left_out[3]
+ sb_1__8_/chanx_left_out[4] sb_1__8_/chanx_left_out[5] sb_1__8_/chanx_left_out[6]
+ sb_1__8_/chanx_left_out[7] sb_1__8_/chanx_left_out[8] sb_1__8_/chanx_left_out[9]
+ sb_1__8_/chanx_left_in[0] sb_1__8_/chanx_left_in[10] sb_1__8_/chanx_left_in[11]
+ sb_1__8_/chanx_left_in[12] sb_1__8_/chanx_left_in[13] sb_1__8_/chanx_left_in[14]
+ sb_1__8_/chanx_left_in[15] sb_1__8_/chanx_left_in[16] sb_1__8_/chanx_left_in[17]
+ sb_1__8_/chanx_left_in[18] sb_1__8_/chanx_left_in[19] sb_1__8_/chanx_left_in[1]
+ sb_1__8_/chanx_left_in[2] sb_1__8_/chanx_left_in[3] sb_1__8_/chanx_left_in[4] sb_1__8_/chanx_left_in[5]
+ sb_1__8_/chanx_left_in[6] sb_1__8_/chanx_left_in[7] sb_1__8_/chanx_left_in[8] sb_1__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
+ cbx_1__8_/prog_clk_0_S_in sb_0__8_/prog_clk_0_E_in cbx_1__8_/top_grid_pin_0_ cbx_1__2_
Xsb_5__5_ sb_5__5_/Test_en_N_out sb_5__5_/Test_en_S_in VGND VPWR sb_5__5_/bottom_left_grid_pin_42_
+ sb_5__5_/bottom_left_grid_pin_43_ sb_5__5_/bottom_left_grid_pin_44_ sb_5__5_/bottom_left_grid_pin_45_
+ sb_5__5_/bottom_left_grid_pin_46_ sb_5__5_/bottom_left_grid_pin_47_ sb_5__5_/bottom_left_grid_pin_48_
+ sb_5__5_/bottom_left_grid_pin_49_ sb_5__5_/ccff_head sb_5__5_/ccff_tail sb_5__5_/chanx_left_in[0]
+ sb_5__5_/chanx_left_in[10] sb_5__5_/chanx_left_in[11] sb_5__5_/chanx_left_in[12]
+ sb_5__5_/chanx_left_in[13] sb_5__5_/chanx_left_in[14] sb_5__5_/chanx_left_in[15]
+ sb_5__5_/chanx_left_in[16] sb_5__5_/chanx_left_in[17] sb_5__5_/chanx_left_in[18]
+ sb_5__5_/chanx_left_in[19] sb_5__5_/chanx_left_in[1] sb_5__5_/chanx_left_in[2] sb_5__5_/chanx_left_in[3]
+ sb_5__5_/chanx_left_in[4] sb_5__5_/chanx_left_in[5] sb_5__5_/chanx_left_in[6] sb_5__5_/chanx_left_in[7]
+ sb_5__5_/chanx_left_in[8] sb_5__5_/chanx_left_in[9] sb_5__5_/chanx_left_out[0] sb_5__5_/chanx_left_out[10]
+ sb_5__5_/chanx_left_out[11] sb_5__5_/chanx_left_out[12] sb_5__5_/chanx_left_out[13]
+ sb_5__5_/chanx_left_out[14] sb_5__5_/chanx_left_out[15] sb_5__5_/chanx_left_out[16]
+ sb_5__5_/chanx_left_out[17] sb_5__5_/chanx_left_out[18] sb_5__5_/chanx_left_out[19]
+ sb_5__5_/chanx_left_out[1] sb_5__5_/chanx_left_out[2] sb_5__5_/chanx_left_out[3]
+ sb_5__5_/chanx_left_out[4] sb_5__5_/chanx_left_out[5] sb_5__5_/chanx_left_out[6]
+ sb_5__5_/chanx_left_out[7] sb_5__5_/chanx_left_out[8] sb_5__5_/chanx_left_out[9]
+ sb_5__5_/chanx_right_in[0] sb_5__5_/chanx_right_in[10] sb_5__5_/chanx_right_in[11]
+ sb_5__5_/chanx_right_in[12] sb_5__5_/chanx_right_in[13] sb_5__5_/chanx_right_in[14]
+ sb_5__5_/chanx_right_in[15] sb_5__5_/chanx_right_in[16] sb_5__5_/chanx_right_in[17]
+ sb_5__5_/chanx_right_in[18] sb_5__5_/chanx_right_in[19] sb_5__5_/chanx_right_in[1]
+ sb_5__5_/chanx_right_in[2] sb_5__5_/chanx_right_in[3] sb_5__5_/chanx_right_in[4]
+ sb_5__5_/chanx_right_in[5] sb_5__5_/chanx_right_in[6] sb_5__5_/chanx_right_in[7]
+ sb_5__5_/chanx_right_in[8] sb_5__5_/chanx_right_in[9] cbx_6__5_/chanx_left_in[0]
+ cbx_6__5_/chanx_left_in[10] cbx_6__5_/chanx_left_in[11] cbx_6__5_/chanx_left_in[12]
+ cbx_6__5_/chanx_left_in[13] cbx_6__5_/chanx_left_in[14] cbx_6__5_/chanx_left_in[15]
+ cbx_6__5_/chanx_left_in[16] cbx_6__5_/chanx_left_in[17] cbx_6__5_/chanx_left_in[18]
+ cbx_6__5_/chanx_left_in[19] cbx_6__5_/chanx_left_in[1] cbx_6__5_/chanx_left_in[2]
+ cbx_6__5_/chanx_left_in[3] cbx_6__5_/chanx_left_in[4] cbx_6__5_/chanx_left_in[5]
+ cbx_6__5_/chanx_left_in[6] cbx_6__5_/chanx_left_in[7] cbx_6__5_/chanx_left_in[8]
+ cbx_6__5_/chanx_left_in[9] cby_5__5_/chany_top_out[0] cby_5__5_/chany_top_out[10]
+ cby_5__5_/chany_top_out[11] cby_5__5_/chany_top_out[12] cby_5__5_/chany_top_out[13]
+ cby_5__5_/chany_top_out[14] cby_5__5_/chany_top_out[15] cby_5__5_/chany_top_out[16]
+ cby_5__5_/chany_top_out[17] cby_5__5_/chany_top_out[18] cby_5__5_/chany_top_out[19]
+ cby_5__5_/chany_top_out[1] cby_5__5_/chany_top_out[2] cby_5__5_/chany_top_out[3]
+ cby_5__5_/chany_top_out[4] cby_5__5_/chany_top_out[5] cby_5__5_/chany_top_out[6]
+ cby_5__5_/chany_top_out[7] cby_5__5_/chany_top_out[8] cby_5__5_/chany_top_out[9]
+ cby_5__5_/chany_top_in[0] cby_5__5_/chany_top_in[10] cby_5__5_/chany_top_in[11]
+ cby_5__5_/chany_top_in[12] cby_5__5_/chany_top_in[13] cby_5__5_/chany_top_in[14]
+ cby_5__5_/chany_top_in[15] cby_5__5_/chany_top_in[16] cby_5__5_/chany_top_in[17]
+ cby_5__5_/chany_top_in[18] cby_5__5_/chany_top_in[19] cby_5__5_/chany_top_in[1]
+ cby_5__5_/chany_top_in[2] cby_5__5_/chany_top_in[3] cby_5__5_/chany_top_in[4] cby_5__5_/chany_top_in[5]
+ cby_5__5_/chany_top_in[6] cby_5__5_/chany_top_in[7] cby_5__5_/chany_top_in[8] cby_5__5_/chany_top_in[9]
+ sb_5__5_/chany_top_in[0] sb_5__5_/chany_top_in[10] sb_5__5_/chany_top_in[11] sb_5__5_/chany_top_in[12]
+ sb_5__5_/chany_top_in[13] sb_5__5_/chany_top_in[14] sb_5__5_/chany_top_in[15] sb_5__5_/chany_top_in[16]
+ sb_5__5_/chany_top_in[17] sb_5__5_/chany_top_in[18] sb_5__5_/chany_top_in[19] sb_5__5_/chany_top_in[1]
+ sb_5__5_/chany_top_in[2] sb_5__5_/chany_top_in[3] sb_5__5_/chany_top_in[4] sb_5__5_/chany_top_in[5]
+ sb_5__5_/chany_top_in[6] sb_5__5_/chany_top_in[7] sb_5__5_/chany_top_in[8] sb_5__5_/chany_top_in[9]
+ sb_5__5_/chany_top_out[0] sb_5__5_/chany_top_out[10] sb_5__5_/chany_top_out[11]
+ sb_5__5_/chany_top_out[12] sb_5__5_/chany_top_out[13] sb_5__5_/chany_top_out[14]
+ sb_5__5_/chany_top_out[15] sb_5__5_/chany_top_out[16] sb_5__5_/chany_top_out[17]
+ sb_5__5_/chany_top_out[18] sb_5__5_/chany_top_out[19] sb_5__5_/chany_top_out[1]
+ sb_5__5_/chany_top_out[2] sb_5__5_/chany_top_out[3] sb_5__5_/chany_top_out[4] sb_5__5_/chany_top_out[5]
+ sb_5__5_/chany_top_out[6] sb_5__5_/chany_top_out[7] sb_5__5_/chany_top_out[8] sb_5__5_/chany_top_out[9]
+ sb_5__5_/clk_1_E_out sb_5__5_/clk_1_N_in sb_5__5_/clk_1_W_out sb_5__5_/clk_2_E_out
+ sb_5__5_/clk_2_N_in sb_5__5_/clk_2_N_out sb_5__5_/clk_2_S_out sb_5__5_/clk_2_W_out
+ sb_5__5_/clk_3_E_out sb_5__5_/clk_3_N_in sb_5__5_/clk_3_N_out sb_5__5_/clk_3_S_out
+ sb_5__5_/clk_3_W_out sb_5__5_/left_bottom_grid_pin_34_ sb_5__5_/left_bottom_grid_pin_35_
+ sb_5__5_/left_bottom_grid_pin_36_ sb_5__5_/left_bottom_grid_pin_37_ sb_5__5_/left_bottom_grid_pin_38_
+ sb_5__5_/left_bottom_grid_pin_39_ sb_5__5_/left_bottom_grid_pin_40_ sb_5__5_/left_bottom_grid_pin_41_
+ sb_5__5_/prog_clk_0_N_in sb_5__5_/prog_clk_1_E_out sb_5__5_/prog_clk_1_N_in sb_5__5_/prog_clk_1_W_out
+ sb_5__5_/prog_clk_2_E_out sb_5__5_/prog_clk_2_N_in sb_5__5_/prog_clk_2_N_out sb_5__5_/prog_clk_2_S_out
+ sb_5__5_/prog_clk_2_W_out sb_5__5_/prog_clk_3_E_out sb_5__5_/prog_clk_3_N_in sb_5__5_/prog_clk_3_N_out
+ sb_5__5_/prog_clk_3_S_out sb_5__5_/prog_clk_3_W_out sb_5__5_/right_bottom_grid_pin_34_
+ sb_5__5_/right_bottom_grid_pin_35_ sb_5__5_/right_bottom_grid_pin_36_ sb_5__5_/right_bottom_grid_pin_37_
+ sb_5__5_/right_bottom_grid_pin_38_ sb_5__5_/right_bottom_grid_pin_39_ sb_5__5_/right_bottom_grid_pin_40_
+ sb_5__5_/right_bottom_grid_pin_41_ sb_5__5_/top_left_grid_pin_42_ sb_5__5_/top_left_grid_pin_43_
+ sb_5__5_/top_left_grid_pin_44_ sb_5__5_/top_left_grid_pin_45_ sb_5__5_/top_left_grid_pin_46_
+ sb_5__5_/top_left_grid_pin_47_ sb_5__5_/top_left_grid_pin_48_ sb_5__5_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_8__1_ IO_ISOL_N VGND VPWR cby_8__1_/ccff_head sb_8__0_/ccff_head sb_8__0_/chany_top_out[0]
+ sb_8__0_/chany_top_out[10] sb_8__0_/chany_top_out[11] sb_8__0_/chany_top_out[12]
+ sb_8__0_/chany_top_out[13] sb_8__0_/chany_top_out[14] sb_8__0_/chany_top_out[15]
+ sb_8__0_/chany_top_out[16] sb_8__0_/chany_top_out[17] sb_8__0_/chany_top_out[18]
+ sb_8__0_/chany_top_out[19] sb_8__0_/chany_top_out[1] sb_8__0_/chany_top_out[2] sb_8__0_/chany_top_out[3]
+ sb_8__0_/chany_top_out[4] sb_8__0_/chany_top_out[5] sb_8__0_/chany_top_out[6] sb_8__0_/chany_top_out[7]
+ sb_8__0_/chany_top_out[8] sb_8__0_/chany_top_out[9] sb_8__0_/chany_top_in[0] sb_8__0_/chany_top_in[10]
+ sb_8__0_/chany_top_in[11] sb_8__0_/chany_top_in[12] sb_8__0_/chany_top_in[13] sb_8__0_/chany_top_in[14]
+ sb_8__0_/chany_top_in[15] sb_8__0_/chany_top_in[16] sb_8__0_/chany_top_in[17] sb_8__0_/chany_top_in[18]
+ sb_8__0_/chany_top_in[19] sb_8__0_/chany_top_in[1] sb_8__0_/chany_top_in[2] sb_8__0_/chany_top_in[3]
+ sb_8__0_/chany_top_in[4] sb_8__0_/chany_top_in[5] sb_8__0_/chany_top_in[6] sb_8__0_/chany_top_in[7]
+ sb_8__0_/chany_top_in[8] sb_8__0_/chany_top_in[9] cby_8__1_/chany_top_in[0] cby_8__1_/chany_top_in[10]
+ cby_8__1_/chany_top_in[11] cby_8__1_/chany_top_in[12] cby_8__1_/chany_top_in[13]
+ cby_8__1_/chany_top_in[14] cby_8__1_/chany_top_in[15] cby_8__1_/chany_top_in[16]
+ cby_8__1_/chany_top_in[17] cby_8__1_/chany_top_in[18] cby_8__1_/chany_top_in[19]
+ cby_8__1_/chany_top_in[1] cby_8__1_/chany_top_in[2] cby_8__1_/chany_top_in[3] cby_8__1_/chany_top_in[4]
+ cby_8__1_/chany_top_in[5] cby_8__1_/chany_top_in[6] cby_8__1_/chany_top_in[7] cby_8__1_/chany_top_in[8]
+ cby_8__1_/chany_top_in[9] cby_8__1_/chany_top_out[0] cby_8__1_/chany_top_out[10]
+ cby_8__1_/chany_top_out[11] cby_8__1_/chany_top_out[12] cby_8__1_/chany_top_out[13]
+ cby_8__1_/chany_top_out[14] cby_8__1_/chany_top_out[15] cby_8__1_/chany_top_out[16]
+ cby_8__1_/chany_top_out[17] cby_8__1_/chany_top_out[18] cby_8__1_/chany_top_out[19]
+ cby_8__1_/chany_top_out[1] cby_8__1_/chany_top_out[2] cby_8__1_/chany_top_out[3]
+ cby_8__1_/chany_top_out[4] cby_8__1_/chany_top_out[5] cby_8__1_/chany_top_out[6]
+ cby_8__1_/chany_top_out[7] cby_8__1_/chany_top_out[8] cby_8__1_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
+ cby_8__1_/left_grid_pin_16_ cby_8__1_/left_grid_pin_17_ cby_8__1_/left_grid_pin_18_
+ cby_8__1_/left_grid_pin_19_ cby_8__1_/left_grid_pin_20_ cby_8__1_/left_grid_pin_21_
+ cby_8__1_/left_grid_pin_22_ cby_8__1_/left_grid_pin_23_ cby_8__1_/left_grid_pin_24_
+ cby_8__1_/left_grid_pin_25_ cby_8__1_/left_grid_pin_26_ cby_8__1_/left_grid_pin_27_
+ cby_8__1_/left_grid_pin_28_ cby_8__1_/left_grid_pin_29_ cby_8__1_/left_grid_pin_30_
+ cby_8__1_/left_grid_pin_31_ cby_8__1_/right_grid_pin_0_ sb_8__0_/top_right_grid_pin_1_
+ sb_8__1_/bottom_right_grid_pin_1_ cby_8__1_/prog_clk_0_N_out sb_8__0_/prog_clk_0_N_in
+ cby_8__1_/prog_clk_0_W_in cby_8__1_/right_grid_pin_0_ cby_2__1_
Xsb_2__2_ sb_2__2_/Test_en_N_out sb_2__2_/Test_en_S_in VGND VPWR sb_2__2_/bottom_left_grid_pin_42_
+ sb_2__2_/bottom_left_grid_pin_43_ sb_2__2_/bottom_left_grid_pin_44_ sb_2__2_/bottom_left_grid_pin_45_
+ sb_2__2_/bottom_left_grid_pin_46_ sb_2__2_/bottom_left_grid_pin_47_ sb_2__2_/bottom_left_grid_pin_48_
+ sb_2__2_/bottom_left_grid_pin_49_ sb_2__2_/ccff_head sb_2__2_/ccff_tail sb_2__2_/chanx_left_in[0]
+ sb_2__2_/chanx_left_in[10] sb_2__2_/chanx_left_in[11] sb_2__2_/chanx_left_in[12]
+ sb_2__2_/chanx_left_in[13] sb_2__2_/chanx_left_in[14] sb_2__2_/chanx_left_in[15]
+ sb_2__2_/chanx_left_in[16] sb_2__2_/chanx_left_in[17] sb_2__2_/chanx_left_in[18]
+ sb_2__2_/chanx_left_in[19] sb_2__2_/chanx_left_in[1] sb_2__2_/chanx_left_in[2] sb_2__2_/chanx_left_in[3]
+ sb_2__2_/chanx_left_in[4] sb_2__2_/chanx_left_in[5] sb_2__2_/chanx_left_in[6] sb_2__2_/chanx_left_in[7]
+ sb_2__2_/chanx_left_in[8] sb_2__2_/chanx_left_in[9] sb_2__2_/chanx_left_out[0] sb_2__2_/chanx_left_out[10]
+ sb_2__2_/chanx_left_out[11] sb_2__2_/chanx_left_out[12] sb_2__2_/chanx_left_out[13]
+ sb_2__2_/chanx_left_out[14] sb_2__2_/chanx_left_out[15] sb_2__2_/chanx_left_out[16]
+ sb_2__2_/chanx_left_out[17] sb_2__2_/chanx_left_out[18] sb_2__2_/chanx_left_out[19]
+ sb_2__2_/chanx_left_out[1] sb_2__2_/chanx_left_out[2] sb_2__2_/chanx_left_out[3]
+ sb_2__2_/chanx_left_out[4] sb_2__2_/chanx_left_out[5] sb_2__2_/chanx_left_out[6]
+ sb_2__2_/chanx_left_out[7] sb_2__2_/chanx_left_out[8] sb_2__2_/chanx_left_out[9]
+ sb_2__2_/chanx_right_in[0] sb_2__2_/chanx_right_in[10] sb_2__2_/chanx_right_in[11]
+ sb_2__2_/chanx_right_in[12] sb_2__2_/chanx_right_in[13] sb_2__2_/chanx_right_in[14]
+ sb_2__2_/chanx_right_in[15] sb_2__2_/chanx_right_in[16] sb_2__2_/chanx_right_in[17]
+ sb_2__2_/chanx_right_in[18] sb_2__2_/chanx_right_in[19] sb_2__2_/chanx_right_in[1]
+ sb_2__2_/chanx_right_in[2] sb_2__2_/chanx_right_in[3] sb_2__2_/chanx_right_in[4]
+ sb_2__2_/chanx_right_in[5] sb_2__2_/chanx_right_in[6] sb_2__2_/chanx_right_in[7]
+ sb_2__2_/chanx_right_in[8] sb_2__2_/chanx_right_in[9] cbx_3__2_/chanx_left_in[0]
+ cbx_3__2_/chanx_left_in[10] cbx_3__2_/chanx_left_in[11] cbx_3__2_/chanx_left_in[12]
+ cbx_3__2_/chanx_left_in[13] cbx_3__2_/chanx_left_in[14] cbx_3__2_/chanx_left_in[15]
+ cbx_3__2_/chanx_left_in[16] cbx_3__2_/chanx_left_in[17] cbx_3__2_/chanx_left_in[18]
+ cbx_3__2_/chanx_left_in[19] cbx_3__2_/chanx_left_in[1] cbx_3__2_/chanx_left_in[2]
+ cbx_3__2_/chanx_left_in[3] cbx_3__2_/chanx_left_in[4] cbx_3__2_/chanx_left_in[5]
+ cbx_3__2_/chanx_left_in[6] cbx_3__2_/chanx_left_in[7] cbx_3__2_/chanx_left_in[8]
+ cbx_3__2_/chanx_left_in[9] cby_2__2_/chany_top_out[0] cby_2__2_/chany_top_out[10]
+ cby_2__2_/chany_top_out[11] cby_2__2_/chany_top_out[12] cby_2__2_/chany_top_out[13]
+ cby_2__2_/chany_top_out[14] cby_2__2_/chany_top_out[15] cby_2__2_/chany_top_out[16]
+ cby_2__2_/chany_top_out[17] cby_2__2_/chany_top_out[18] cby_2__2_/chany_top_out[19]
+ cby_2__2_/chany_top_out[1] cby_2__2_/chany_top_out[2] cby_2__2_/chany_top_out[3]
+ cby_2__2_/chany_top_out[4] cby_2__2_/chany_top_out[5] cby_2__2_/chany_top_out[6]
+ cby_2__2_/chany_top_out[7] cby_2__2_/chany_top_out[8] cby_2__2_/chany_top_out[9]
+ cby_2__2_/chany_top_in[0] cby_2__2_/chany_top_in[10] cby_2__2_/chany_top_in[11]
+ cby_2__2_/chany_top_in[12] cby_2__2_/chany_top_in[13] cby_2__2_/chany_top_in[14]
+ cby_2__2_/chany_top_in[15] cby_2__2_/chany_top_in[16] cby_2__2_/chany_top_in[17]
+ cby_2__2_/chany_top_in[18] cby_2__2_/chany_top_in[19] cby_2__2_/chany_top_in[1]
+ cby_2__2_/chany_top_in[2] cby_2__2_/chany_top_in[3] cby_2__2_/chany_top_in[4] cby_2__2_/chany_top_in[5]
+ cby_2__2_/chany_top_in[6] cby_2__2_/chany_top_in[7] cby_2__2_/chany_top_in[8] cby_2__2_/chany_top_in[9]
+ sb_2__2_/chany_top_in[0] sb_2__2_/chany_top_in[10] sb_2__2_/chany_top_in[11] sb_2__2_/chany_top_in[12]
+ sb_2__2_/chany_top_in[13] sb_2__2_/chany_top_in[14] sb_2__2_/chany_top_in[15] sb_2__2_/chany_top_in[16]
+ sb_2__2_/chany_top_in[17] sb_2__2_/chany_top_in[18] sb_2__2_/chany_top_in[19] sb_2__2_/chany_top_in[1]
+ sb_2__2_/chany_top_in[2] sb_2__2_/chany_top_in[3] sb_2__2_/chany_top_in[4] sb_2__2_/chany_top_in[5]
+ sb_2__2_/chany_top_in[6] sb_2__2_/chany_top_in[7] sb_2__2_/chany_top_in[8] sb_2__2_/chany_top_in[9]
+ sb_2__2_/chany_top_out[0] sb_2__2_/chany_top_out[10] sb_2__2_/chany_top_out[11]
+ sb_2__2_/chany_top_out[12] sb_2__2_/chany_top_out[13] sb_2__2_/chany_top_out[14]
+ sb_2__2_/chany_top_out[15] sb_2__2_/chany_top_out[16] sb_2__2_/chany_top_out[17]
+ sb_2__2_/chany_top_out[18] sb_2__2_/chany_top_out[19] sb_2__2_/chany_top_out[1]
+ sb_2__2_/chany_top_out[2] sb_2__2_/chany_top_out[3] sb_2__2_/chany_top_out[4] sb_2__2_/chany_top_out[5]
+ sb_2__2_/chany_top_out[6] sb_2__2_/chany_top_out[7] sb_2__2_/chany_top_out[8] sb_2__2_/chany_top_out[9]
+ sb_2__2_/clk_1_E_out sb_2__2_/clk_1_N_in sb_2__2_/clk_1_W_out sb_2__2_/clk_2_E_out
+ sb_2__2_/clk_2_N_in sb_2__2_/clk_2_N_out sb_2__2_/clk_2_S_out sb_2__2_/clk_2_W_out
+ sb_2__2_/clk_3_E_out sb_2__2_/clk_3_N_in sb_2__2_/clk_3_N_out sb_2__2_/clk_3_S_out
+ sb_2__2_/clk_3_W_out sb_2__2_/left_bottom_grid_pin_34_ sb_2__2_/left_bottom_grid_pin_35_
+ sb_2__2_/left_bottom_grid_pin_36_ sb_2__2_/left_bottom_grid_pin_37_ sb_2__2_/left_bottom_grid_pin_38_
+ sb_2__2_/left_bottom_grid_pin_39_ sb_2__2_/left_bottom_grid_pin_40_ sb_2__2_/left_bottom_grid_pin_41_
+ sb_2__2_/prog_clk_0_N_in sb_2__2_/prog_clk_1_E_out sb_2__2_/prog_clk_1_N_in sb_2__2_/prog_clk_1_W_out
+ sb_2__2_/prog_clk_2_E_out sb_2__2_/prog_clk_2_N_in sb_2__2_/prog_clk_2_N_out sb_2__2_/prog_clk_2_S_out
+ sb_2__2_/prog_clk_2_W_out sb_2__2_/prog_clk_3_E_out sb_2__2_/prog_clk_3_N_in sb_2__2_/prog_clk_3_N_out
+ sb_2__2_/prog_clk_3_S_out sb_2__2_/prog_clk_3_W_out sb_2__2_/right_bottom_grid_pin_34_
+ sb_2__2_/right_bottom_grid_pin_35_ sb_2__2_/right_bottom_grid_pin_36_ sb_2__2_/right_bottom_grid_pin_37_
+ sb_2__2_/right_bottom_grid_pin_38_ sb_2__2_/right_bottom_grid_pin_39_ sb_2__2_/right_bottom_grid_pin_40_
+ sb_2__2_/right_bottom_grid_pin_41_ sb_2__2_/top_left_grid_pin_42_ sb_2__2_/top_left_grid_pin_43_
+ sb_2__2_/top_left_grid_pin_44_ sb_2__2_/top_left_grid_pin_45_ sb_2__2_/top_left_grid_pin_46_
+ sb_2__2_/top_left_grid_pin_47_ sb_2__2_/top_left_grid_pin_48_ sb_2__2_/top_left_grid_pin_49_
+ sb_1__1_
Xcbx_8__2_ cbx_8__2_/REGIN_FEEDTHROUGH cbx_8__2_/REGOUT_FEEDTHROUGH cbx_8__2_/SC_IN_BOT
+ cbx_8__2_/SC_IN_TOP cbx_8__2_/SC_OUT_BOT cbx_8__2_/SC_OUT_TOP VGND VPWR cbx_8__2_/bottom_grid_pin_0_
+ cbx_8__2_/bottom_grid_pin_10_ cbx_8__2_/bottom_grid_pin_11_ cbx_8__2_/bottom_grid_pin_12_
+ cbx_8__2_/bottom_grid_pin_13_ cbx_8__2_/bottom_grid_pin_14_ cbx_8__2_/bottom_grid_pin_15_
+ cbx_8__2_/bottom_grid_pin_1_ cbx_8__2_/bottom_grid_pin_2_ cbx_8__2_/bottom_grid_pin_3_
+ cbx_8__2_/bottom_grid_pin_4_ cbx_8__2_/bottom_grid_pin_5_ cbx_8__2_/bottom_grid_pin_6_
+ cbx_8__2_/bottom_grid_pin_7_ cbx_8__2_/bottom_grid_pin_8_ cbx_8__2_/bottom_grid_pin_9_
+ sb_8__2_/ccff_tail sb_7__2_/ccff_head cbx_8__2_/chanx_left_in[0] cbx_8__2_/chanx_left_in[10]
+ cbx_8__2_/chanx_left_in[11] cbx_8__2_/chanx_left_in[12] cbx_8__2_/chanx_left_in[13]
+ cbx_8__2_/chanx_left_in[14] cbx_8__2_/chanx_left_in[15] cbx_8__2_/chanx_left_in[16]
+ cbx_8__2_/chanx_left_in[17] cbx_8__2_/chanx_left_in[18] cbx_8__2_/chanx_left_in[19]
+ cbx_8__2_/chanx_left_in[1] cbx_8__2_/chanx_left_in[2] cbx_8__2_/chanx_left_in[3]
+ cbx_8__2_/chanx_left_in[4] cbx_8__2_/chanx_left_in[5] cbx_8__2_/chanx_left_in[6]
+ cbx_8__2_/chanx_left_in[7] cbx_8__2_/chanx_left_in[8] cbx_8__2_/chanx_left_in[9]
+ sb_7__2_/chanx_right_in[0] sb_7__2_/chanx_right_in[10] sb_7__2_/chanx_right_in[11]
+ sb_7__2_/chanx_right_in[12] sb_7__2_/chanx_right_in[13] sb_7__2_/chanx_right_in[14]
+ sb_7__2_/chanx_right_in[15] sb_7__2_/chanx_right_in[16] sb_7__2_/chanx_right_in[17]
+ sb_7__2_/chanx_right_in[18] sb_7__2_/chanx_right_in[19] sb_7__2_/chanx_right_in[1]
+ sb_7__2_/chanx_right_in[2] sb_7__2_/chanx_right_in[3] sb_7__2_/chanx_right_in[4]
+ sb_7__2_/chanx_right_in[5] sb_7__2_/chanx_right_in[6] sb_7__2_/chanx_right_in[7]
+ sb_7__2_/chanx_right_in[8] sb_7__2_/chanx_right_in[9] sb_8__2_/chanx_left_out[0]
+ sb_8__2_/chanx_left_out[10] sb_8__2_/chanx_left_out[11] sb_8__2_/chanx_left_out[12]
+ sb_8__2_/chanx_left_out[13] sb_8__2_/chanx_left_out[14] sb_8__2_/chanx_left_out[15]
+ sb_8__2_/chanx_left_out[16] sb_8__2_/chanx_left_out[17] sb_8__2_/chanx_left_out[18]
+ sb_8__2_/chanx_left_out[19] sb_8__2_/chanx_left_out[1] sb_8__2_/chanx_left_out[2]
+ sb_8__2_/chanx_left_out[3] sb_8__2_/chanx_left_out[4] sb_8__2_/chanx_left_out[5]
+ sb_8__2_/chanx_left_out[6] sb_8__2_/chanx_left_out[7] sb_8__2_/chanx_left_out[8]
+ sb_8__2_/chanx_left_out[9] sb_8__2_/chanx_left_in[0] sb_8__2_/chanx_left_in[10]
+ sb_8__2_/chanx_left_in[11] sb_8__2_/chanx_left_in[12] sb_8__2_/chanx_left_in[13]
+ sb_8__2_/chanx_left_in[14] sb_8__2_/chanx_left_in[15] sb_8__2_/chanx_left_in[16]
+ sb_8__2_/chanx_left_in[17] sb_8__2_/chanx_left_in[18] sb_8__2_/chanx_left_in[19]
+ sb_8__2_/chanx_left_in[1] sb_8__2_/chanx_left_in[2] sb_8__2_/chanx_left_in[3] sb_8__2_/chanx_left_in[4]
+ sb_8__2_/chanx_left_in[5] sb_8__2_/chanx_left_in[6] sb_8__2_/chanx_left_in[7] sb_8__2_/chanx_left_in[8]
+ sb_8__2_/chanx_left_in[9] cbx_8__2_/clk_1_N_out cbx_8__2_/clk_1_S_out cbx_8__2_/clk_1_W_in
+ cbx_8__2_/clk_2_E_out cbx_8__2_/clk_2_W_in cbx_8__2_/clk_2_W_out cbx_8__2_/clk_3_E_out
+ cbx_8__2_/clk_3_W_in cbx_8__2_/clk_3_W_out cbx_8__2_/prog_clk_0_N_in cbx_8__2_/prog_clk_0_W_out
+ cbx_8__2_/prog_clk_1_N_out cbx_8__2_/prog_clk_1_S_out cbx_8__2_/prog_clk_1_W_in
+ cbx_8__2_/prog_clk_2_E_out cbx_8__2_/prog_clk_2_W_in cbx_8__2_/prog_clk_2_W_out
+ cbx_8__2_/prog_clk_3_E_out cbx_8__2_/prog_clk_3_W_in cbx_8__2_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_8__7_ VGND VPWR sb_8__7_/bottom_left_grid_pin_42_ sb_8__7_/bottom_left_grid_pin_43_
+ sb_8__7_/bottom_left_grid_pin_44_ sb_8__7_/bottom_left_grid_pin_45_ sb_8__7_/bottom_left_grid_pin_46_
+ sb_8__7_/bottom_left_grid_pin_47_ sb_8__7_/bottom_left_grid_pin_48_ sb_8__7_/bottom_left_grid_pin_49_
+ sb_8__7_/bottom_right_grid_pin_1_ sb_8__7_/ccff_head sb_8__7_/ccff_tail sb_8__7_/chanx_left_in[0]
+ sb_8__7_/chanx_left_in[10] sb_8__7_/chanx_left_in[11] sb_8__7_/chanx_left_in[12]
+ sb_8__7_/chanx_left_in[13] sb_8__7_/chanx_left_in[14] sb_8__7_/chanx_left_in[15]
+ sb_8__7_/chanx_left_in[16] sb_8__7_/chanx_left_in[17] sb_8__7_/chanx_left_in[18]
+ sb_8__7_/chanx_left_in[19] sb_8__7_/chanx_left_in[1] sb_8__7_/chanx_left_in[2] sb_8__7_/chanx_left_in[3]
+ sb_8__7_/chanx_left_in[4] sb_8__7_/chanx_left_in[5] sb_8__7_/chanx_left_in[6] sb_8__7_/chanx_left_in[7]
+ sb_8__7_/chanx_left_in[8] sb_8__7_/chanx_left_in[9] sb_8__7_/chanx_left_out[0] sb_8__7_/chanx_left_out[10]
+ sb_8__7_/chanx_left_out[11] sb_8__7_/chanx_left_out[12] sb_8__7_/chanx_left_out[13]
+ sb_8__7_/chanx_left_out[14] sb_8__7_/chanx_left_out[15] sb_8__7_/chanx_left_out[16]
+ sb_8__7_/chanx_left_out[17] sb_8__7_/chanx_left_out[18] sb_8__7_/chanx_left_out[19]
+ sb_8__7_/chanx_left_out[1] sb_8__7_/chanx_left_out[2] sb_8__7_/chanx_left_out[3]
+ sb_8__7_/chanx_left_out[4] sb_8__7_/chanx_left_out[5] sb_8__7_/chanx_left_out[6]
+ sb_8__7_/chanx_left_out[7] sb_8__7_/chanx_left_out[8] sb_8__7_/chanx_left_out[9]
+ cby_8__7_/chany_top_out[0] cby_8__7_/chany_top_out[10] cby_8__7_/chany_top_out[11]
+ cby_8__7_/chany_top_out[12] cby_8__7_/chany_top_out[13] cby_8__7_/chany_top_out[14]
+ cby_8__7_/chany_top_out[15] cby_8__7_/chany_top_out[16] cby_8__7_/chany_top_out[17]
+ cby_8__7_/chany_top_out[18] cby_8__7_/chany_top_out[19] cby_8__7_/chany_top_out[1]
+ cby_8__7_/chany_top_out[2] cby_8__7_/chany_top_out[3] cby_8__7_/chany_top_out[4]
+ cby_8__7_/chany_top_out[5] cby_8__7_/chany_top_out[6] cby_8__7_/chany_top_out[7]
+ cby_8__7_/chany_top_out[8] cby_8__7_/chany_top_out[9] cby_8__7_/chany_top_in[0]
+ cby_8__7_/chany_top_in[10] cby_8__7_/chany_top_in[11] cby_8__7_/chany_top_in[12]
+ cby_8__7_/chany_top_in[13] cby_8__7_/chany_top_in[14] cby_8__7_/chany_top_in[15]
+ cby_8__7_/chany_top_in[16] cby_8__7_/chany_top_in[17] cby_8__7_/chany_top_in[18]
+ cby_8__7_/chany_top_in[19] cby_8__7_/chany_top_in[1] cby_8__7_/chany_top_in[2] cby_8__7_/chany_top_in[3]
+ cby_8__7_/chany_top_in[4] cby_8__7_/chany_top_in[5] cby_8__7_/chany_top_in[6] cby_8__7_/chany_top_in[7]
+ cby_8__7_/chany_top_in[8] cby_8__7_/chany_top_in[9] sb_8__7_/chany_top_in[0] sb_8__7_/chany_top_in[10]
+ sb_8__7_/chany_top_in[11] sb_8__7_/chany_top_in[12] sb_8__7_/chany_top_in[13] sb_8__7_/chany_top_in[14]
+ sb_8__7_/chany_top_in[15] sb_8__7_/chany_top_in[16] sb_8__7_/chany_top_in[17] sb_8__7_/chany_top_in[18]
+ sb_8__7_/chany_top_in[19] sb_8__7_/chany_top_in[1] sb_8__7_/chany_top_in[2] sb_8__7_/chany_top_in[3]
+ sb_8__7_/chany_top_in[4] sb_8__7_/chany_top_in[5] sb_8__7_/chany_top_in[6] sb_8__7_/chany_top_in[7]
+ sb_8__7_/chany_top_in[8] sb_8__7_/chany_top_in[9] sb_8__7_/chany_top_out[0] sb_8__7_/chany_top_out[10]
+ sb_8__7_/chany_top_out[11] sb_8__7_/chany_top_out[12] sb_8__7_/chany_top_out[13]
+ sb_8__7_/chany_top_out[14] sb_8__7_/chany_top_out[15] sb_8__7_/chany_top_out[16]
+ sb_8__7_/chany_top_out[17] sb_8__7_/chany_top_out[18] sb_8__7_/chany_top_out[19]
+ sb_8__7_/chany_top_out[1] sb_8__7_/chany_top_out[2] sb_8__7_/chany_top_out[3] sb_8__7_/chany_top_out[4]
+ sb_8__7_/chany_top_out[5] sb_8__7_/chany_top_out[6] sb_8__7_/chany_top_out[7] sb_8__7_/chany_top_out[8]
+ sb_8__7_/chany_top_out[9] sb_8__7_/left_bottom_grid_pin_34_ sb_8__7_/left_bottom_grid_pin_35_
+ sb_8__7_/left_bottom_grid_pin_36_ sb_8__7_/left_bottom_grid_pin_37_ sb_8__7_/left_bottom_grid_pin_38_
+ sb_8__7_/left_bottom_grid_pin_39_ sb_8__7_/left_bottom_grid_pin_40_ sb_8__7_/left_bottom_grid_pin_41_
+ sb_8__7_/prog_clk_0_N_in sb_8__7_/top_left_grid_pin_42_ sb_8__7_/top_left_grid_pin_43_
+ sb_8__7_/top_left_grid_pin_44_ sb_8__7_/top_left_grid_pin_45_ sb_8__7_/top_left_grid_pin_46_
+ sb_8__7_/top_left_grid_pin_47_ sb_8__7_/top_left_grid_pin_48_ sb_8__7_/top_left_grid_pin_49_
+ sb_8__7_/top_right_grid_pin_1_ sb_2__1_
Xcby_1__6_ cby_1__6_/Test_en_W_in cby_1__6_/Test_en_E_out cby_1__6_/Test_en_N_out
+ cby_1__6_/Test_en_W_in cby_1__6_/Test_en_W_in cby_1__6_/Test_en_W_out VGND VPWR
+ cby_1__6_/ccff_head cby_1__6_/ccff_tail sb_1__5_/chany_top_out[0] sb_1__5_/chany_top_out[10]
+ sb_1__5_/chany_top_out[11] sb_1__5_/chany_top_out[12] sb_1__5_/chany_top_out[13]
+ sb_1__5_/chany_top_out[14] sb_1__5_/chany_top_out[15] sb_1__5_/chany_top_out[16]
+ sb_1__5_/chany_top_out[17] sb_1__5_/chany_top_out[18] sb_1__5_/chany_top_out[19]
+ sb_1__5_/chany_top_out[1] sb_1__5_/chany_top_out[2] sb_1__5_/chany_top_out[3] sb_1__5_/chany_top_out[4]
+ sb_1__5_/chany_top_out[5] sb_1__5_/chany_top_out[6] sb_1__5_/chany_top_out[7] sb_1__5_/chany_top_out[8]
+ sb_1__5_/chany_top_out[9] sb_1__5_/chany_top_in[0] sb_1__5_/chany_top_in[10] sb_1__5_/chany_top_in[11]
+ sb_1__5_/chany_top_in[12] sb_1__5_/chany_top_in[13] sb_1__5_/chany_top_in[14] sb_1__5_/chany_top_in[15]
+ sb_1__5_/chany_top_in[16] sb_1__5_/chany_top_in[17] sb_1__5_/chany_top_in[18] sb_1__5_/chany_top_in[19]
+ sb_1__5_/chany_top_in[1] sb_1__5_/chany_top_in[2] sb_1__5_/chany_top_in[3] sb_1__5_/chany_top_in[4]
+ sb_1__5_/chany_top_in[5] sb_1__5_/chany_top_in[6] sb_1__5_/chany_top_in[7] sb_1__5_/chany_top_in[8]
+ sb_1__5_/chany_top_in[9] cby_1__6_/chany_top_in[0] cby_1__6_/chany_top_in[10] cby_1__6_/chany_top_in[11]
+ cby_1__6_/chany_top_in[12] cby_1__6_/chany_top_in[13] cby_1__6_/chany_top_in[14]
+ cby_1__6_/chany_top_in[15] cby_1__6_/chany_top_in[16] cby_1__6_/chany_top_in[17]
+ cby_1__6_/chany_top_in[18] cby_1__6_/chany_top_in[19] cby_1__6_/chany_top_in[1]
+ cby_1__6_/chany_top_in[2] cby_1__6_/chany_top_in[3] cby_1__6_/chany_top_in[4] cby_1__6_/chany_top_in[5]
+ cby_1__6_/chany_top_in[6] cby_1__6_/chany_top_in[7] cby_1__6_/chany_top_in[8] cby_1__6_/chany_top_in[9]
+ cby_1__6_/chany_top_out[0] cby_1__6_/chany_top_out[10] cby_1__6_/chany_top_out[11]
+ cby_1__6_/chany_top_out[12] cby_1__6_/chany_top_out[13] cby_1__6_/chany_top_out[14]
+ cby_1__6_/chany_top_out[15] cby_1__6_/chany_top_out[16] cby_1__6_/chany_top_out[17]
+ cby_1__6_/chany_top_out[18] cby_1__6_/chany_top_out[19] cby_1__6_/chany_top_out[1]
+ cby_1__6_/chany_top_out[2] cby_1__6_/chany_top_out[3] cby_1__6_/chany_top_out[4]
+ cby_1__6_/chany_top_out[5] cby_1__6_/chany_top_out[6] cby_1__6_/chany_top_out[7]
+ cby_1__6_/chany_top_out[8] cby_1__6_/chany_top_out[9] cby_1__6_/clk_2_N_out sb_1__6_/clk_2_S_out
+ sb_1__5_/clk_1_N_in cby_1__6_/clk_3_N_out cby_1__6_/clk_3_S_in cby_1__6_/clk_3_S_out
+ cby_1__6_/left_grid_pin_16_ cby_1__6_/left_grid_pin_17_ cby_1__6_/left_grid_pin_18_
+ cby_1__6_/left_grid_pin_19_ cby_1__6_/left_grid_pin_20_ cby_1__6_/left_grid_pin_21_
+ cby_1__6_/left_grid_pin_22_ cby_1__6_/left_grid_pin_23_ cby_1__6_/left_grid_pin_24_
+ cby_1__6_/left_grid_pin_25_ cby_1__6_/left_grid_pin_26_ cby_1__6_/left_grid_pin_27_
+ cby_1__6_/left_grid_pin_28_ cby_1__6_/left_grid_pin_29_ cby_1__6_/left_grid_pin_30_
+ cby_1__6_/left_grid_pin_31_ cby_1__6_/prog_clk_0_N_out sb_1__5_/prog_clk_0_N_in
+ cby_1__6_/prog_clk_0_W_in cby_1__6_/prog_clk_2_N_out sb_1__6_/prog_clk_2_S_out sb_1__5_/prog_clk_1_N_in
+ cby_1__6_/prog_clk_3_N_out cby_1__6_/prog_clk_3_S_in cby_1__6_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_7__2_ cbx_7__2_/SC_OUT_BOT cbx_7__1_/SC_IN_TOP grid_clb_7__2_/SC_OUT_TOP
+ cby_6__2_/Test_en_E_out cby_7__2_/Test_en_W_in cby_6__2_/Test_en_E_out grid_clb_7__2_/Test_en_W_out
+ VGND VPWR cbx_7__1_/REGIN_FEEDTHROUGH grid_clb_7__2_/bottom_width_0_height_0__pin_51_
+ cby_6__2_/ccff_tail cby_7__2_/ccff_head cbx_7__1_/clk_1_N_out cbx_7__1_/clk_1_N_out
+ cby_7__2_/prog_clk_0_W_in cbx_7__1_/prog_clk_1_N_out grid_clb_7__2_/prog_clk_0_N_out
+ cbx_7__1_/prog_clk_1_N_out cbx_7__1_/prog_clk_0_N_in grid_clb_7__2_/prog_clk_0_W_out
+ cby_7__2_/left_grid_pin_16_ cby_7__2_/left_grid_pin_17_ cby_7__2_/left_grid_pin_18_
+ cby_7__2_/left_grid_pin_19_ cby_7__2_/left_grid_pin_20_ cby_7__2_/left_grid_pin_21_
+ cby_7__2_/left_grid_pin_22_ cby_7__2_/left_grid_pin_23_ cby_7__2_/left_grid_pin_24_
+ cby_7__2_/left_grid_pin_25_ cby_7__2_/left_grid_pin_26_ cby_7__2_/left_grid_pin_27_
+ cby_7__2_/left_grid_pin_28_ cby_7__2_/left_grid_pin_29_ cby_7__2_/left_grid_pin_30_
+ cby_7__2_/left_grid_pin_31_ sb_7__1_/top_left_grid_pin_42_ sb_7__2_/bottom_left_grid_pin_42_
+ sb_7__1_/top_left_grid_pin_43_ sb_7__2_/bottom_left_grid_pin_43_ sb_7__1_/top_left_grid_pin_44_
+ sb_7__2_/bottom_left_grid_pin_44_ sb_7__1_/top_left_grid_pin_45_ sb_7__2_/bottom_left_grid_pin_45_
+ sb_7__1_/top_left_grid_pin_46_ sb_7__2_/bottom_left_grid_pin_46_ sb_7__1_/top_left_grid_pin_47_
+ sb_7__2_/bottom_left_grid_pin_47_ sb_7__1_/top_left_grid_pin_48_ sb_7__2_/bottom_left_grid_pin_48_
+ sb_7__1_/top_left_grid_pin_49_ sb_7__2_/bottom_left_grid_pin_49_ cbx_7__2_/bottom_grid_pin_0_
+ cbx_7__2_/bottom_grid_pin_10_ cbx_7__2_/bottom_grid_pin_11_ cbx_7__2_/bottom_grid_pin_12_
+ cbx_7__2_/bottom_grid_pin_13_ cbx_7__2_/bottom_grid_pin_14_ cbx_7__2_/bottom_grid_pin_15_
+ cbx_7__2_/bottom_grid_pin_1_ cbx_7__2_/bottom_grid_pin_2_ cbx_7__2_/REGOUT_FEEDTHROUGH
+ grid_clb_7__2_/top_width_0_height_0__pin_33_ sb_7__2_/left_bottom_grid_pin_34_ sb_6__2_/right_bottom_grid_pin_34_
+ sb_7__2_/left_bottom_grid_pin_35_ sb_6__2_/right_bottom_grid_pin_35_ sb_7__2_/left_bottom_grid_pin_36_
+ sb_6__2_/right_bottom_grid_pin_36_ sb_7__2_/left_bottom_grid_pin_37_ sb_6__2_/right_bottom_grid_pin_37_
+ sb_7__2_/left_bottom_grid_pin_38_ sb_6__2_/right_bottom_grid_pin_38_ sb_7__2_/left_bottom_grid_pin_39_
+ sb_6__2_/right_bottom_grid_pin_39_ cbx_7__2_/bottom_grid_pin_3_ sb_7__2_/left_bottom_grid_pin_40_
+ sb_6__2_/right_bottom_grid_pin_40_ sb_7__2_/left_bottom_grid_pin_41_ sb_6__2_/right_bottom_grid_pin_41_
+ cbx_7__2_/bottom_grid_pin_4_ cbx_7__2_/bottom_grid_pin_5_ cbx_7__2_/bottom_grid_pin_6_
+ cbx_7__2_/bottom_grid_pin_7_ cbx_7__2_/bottom_grid_pin_8_ cbx_7__2_/bottom_grid_pin_9_
+ grid_clb
Xcbx_1__7_ cbx_1__7_/REGIN_FEEDTHROUGH cbx_1__7_/REGOUT_FEEDTHROUGH cbx_1__7_/SC_IN_BOT
+ cbx_1__7_/SC_IN_TOP cbx_1__7_/SC_OUT_BOT cbx_1__7_/SC_OUT_TOP VGND VPWR cbx_1__7_/bottom_grid_pin_0_
+ cbx_1__7_/bottom_grid_pin_10_ cbx_1__7_/bottom_grid_pin_11_ cbx_1__7_/bottom_grid_pin_12_
+ cbx_1__7_/bottom_grid_pin_13_ cbx_1__7_/bottom_grid_pin_14_ cbx_1__7_/bottom_grid_pin_15_
+ cbx_1__7_/bottom_grid_pin_1_ cbx_1__7_/bottom_grid_pin_2_ cbx_1__7_/bottom_grid_pin_3_
+ cbx_1__7_/bottom_grid_pin_4_ cbx_1__7_/bottom_grid_pin_5_ cbx_1__7_/bottom_grid_pin_6_
+ cbx_1__7_/bottom_grid_pin_7_ cbx_1__7_/bottom_grid_pin_8_ cbx_1__7_/bottom_grid_pin_9_
+ sb_1__7_/ccff_tail sb_0__7_/ccff_head cbx_1__7_/chanx_left_in[0] cbx_1__7_/chanx_left_in[10]
+ cbx_1__7_/chanx_left_in[11] cbx_1__7_/chanx_left_in[12] cbx_1__7_/chanx_left_in[13]
+ cbx_1__7_/chanx_left_in[14] cbx_1__7_/chanx_left_in[15] cbx_1__7_/chanx_left_in[16]
+ cbx_1__7_/chanx_left_in[17] cbx_1__7_/chanx_left_in[18] cbx_1__7_/chanx_left_in[19]
+ cbx_1__7_/chanx_left_in[1] cbx_1__7_/chanx_left_in[2] cbx_1__7_/chanx_left_in[3]
+ cbx_1__7_/chanx_left_in[4] cbx_1__7_/chanx_left_in[5] cbx_1__7_/chanx_left_in[6]
+ cbx_1__7_/chanx_left_in[7] cbx_1__7_/chanx_left_in[8] cbx_1__7_/chanx_left_in[9]
+ sb_0__7_/chanx_right_in[0] sb_0__7_/chanx_right_in[10] sb_0__7_/chanx_right_in[11]
+ sb_0__7_/chanx_right_in[12] sb_0__7_/chanx_right_in[13] sb_0__7_/chanx_right_in[14]
+ sb_0__7_/chanx_right_in[15] sb_0__7_/chanx_right_in[16] sb_0__7_/chanx_right_in[17]
+ sb_0__7_/chanx_right_in[18] sb_0__7_/chanx_right_in[19] sb_0__7_/chanx_right_in[1]
+ sb_0__7_/chanx_right_in[2] sb_0__7_/chanx_right_in[3] sb_0__7_/chanx_right_in[4]
+ sb_0__7_/chanx_right_in[5] sb_0__7_/chanx_right_in[6] sb_0__7_/chanx_right_in[7]
+ sb_0__7_/chanx_right_in[8] sb_0__7_/chanx_right_in[9] sb_1__7_/chanx_left_out[0]
+ sb_1__7_/chanx_left_out[10] sb_1__7_/chanx_left_out[11] sb_1__7_/chanx_left_out[12]
+ sb_1__7_/chanx_left_out[13] sb_1__7_/chanx_left_out[14] sb_1__7_/chanx_left_out[15]
+ sb_1__7_/chanx_left_out[16] sb_1__7_/chanx_left_out[17] sb_1__7_/chanx_left_out[18]
+ sb_1__7_/chanx_left_out[19] sb_1__7_/chanx_left_out[1] sb_1__7_/chanx_left_out[2]
+ sb_1__7_/chanx_left_out[3] sb_1__7_/chanx_left_out[4] sb_1__7_/chanx_left_out[5]
+ sb_1__7_/chanx_left_out[6] sb_1__7_/chanx_left_out[7] sb_1__7_/chanx_left_out[8]
+ sb_1__7_/chanx_left_out[9] sb_1__7_/chanx_left_in[0] sb_1__7_/chanx_left_in[10]
+ sb_1__7_/chanx_left_in[11] sb_1__7_/chanx_left_in[12] sb_1__7_/chanx_left_in[13]
+ sb_1__7_/chanx_left_in[14] sb_1__7_/chanx_left_in[15] sb_1__7_/chanx_left_in[16]
+ sb_1__7_/chanx_left_in[17] sb_1__7_/chanx_left_in[18] sb_1__7_/chanx_left_in[19]
+ sb_1__7_/chanx_left_in[1] sb_1__7_/chanx_left_in[2] sb_1__7_/chanx_left_in[3] sb_1__7_/chanx_left_in[4]
+ sb_1__7_/chanx_left_in[5] sb_1__7_/chanx_left_in[6] sb_1__7_/chanx_left_in[7] sb_1__7_/chanx_left_in[8]
+ sb_1__7_/chanx_left_in[9] cbx_1__7_/clk_1_N_out cbx_1__7_/clk_1_S_out sb_1__7_/clk_1_W_out
+ cbx_1__7_/clk_2_E_out cbx_1__7_/clk_2_W_in cbx_1__7_/clk_2_W_out cbx_1__7_/clk_3_E_out
+ cbx_1__7_/clk_3_W_in cbx_1__7_/clk_3_W_out cbx_1__7_/prog_clk_0_N_in sb_0__7_/prog_clk_0_E_in
+ cbx_1__7_/prog_clk_1_N_out cbx_1__7_/prog_clk_1_S_out sb_1__7_/prog_clk_1_W_out
+ cbx_1__7_/prog_clk_2_E_out cbx_1__7_/prog_clk_2_W_in cbx_1__7_/prog_clk_2_W_out
+ cbx_1__7_/prog_clk_3_E_out cbx_1__7_/prog_clk_3_W_in cbx_1__7_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_5__4_ sb_5__4_/Test_en_N_out sb_5__4_/Test_en_S_in VGND VPWR sb_5__4_/bottom_left_grid_pin_42_
+ sb_5__4_/bottom_left_grid_pin_43_ sb_5__4_/bottom_left_grid_pin_44_ sb_5__4_/bottom_left_grid_pin_45_
+ sb_5__4_/bottom_left_grid_pin_46_ sb_5__4_/bottom_left_grid_pin_47_ sb_5__4_/bottom_left_grid_pin_48_
+ sb_5__4_/bottom_left_grid_pin_49_ sb_5__4_/ccff_head sb_5__4_/ccff_tail sb_5__4_/chanx_left_in[0]
+ sb_5__4_/chanx_left_in[10] sb_5__4_/chanx_left_in[11] sb_5__4_/chanx_left_in[12]
+ sb_5__4_/chanx_left_in[13] sb_5__4_/chanx_left_in[14] sb_5__4_/chanx_left_in[15]
+ sb_5__4_/chanx_left_in[16] sb_5__4_/chanx_left_in[17] sb_5__4_/chanx_left_in[18]
+ sb_5__4_/chanx_left_in[19] sb_5__4_/chanx_left_in[1] sb_5__4_/chanx_left_in[2] sb_5__4_/chanx_left_in[3]
+ sb_5__4_/chanx_left_in[4] sb_5__4_/chanx_left_in[5] sb_5__4_/chanx_left_in[6] sb_5__4_/chanx_left_in[7]
+ sb_5__4_/chanx_left_in[8] sb_5__4_/chanx_left_in[9] sb_5__4_/chanx_left_out[0] sb_5__4_/chanx_left_out[10]
+ sb_5__4_/chanx_left_out[11] sb_5__4_/chanx_left_out[12] sb_5__4_/chanx_left_out[13]
+ sb_5__4_/chanx_left_out[14] sb_5__4_/chanx_left_out[15] sb_5__4_/chanx_left_out[16]
+ sb_5__4_/chanx_left_out[17] sb_5__4_/chanx_left_out[18] sb_5__4_/chanx_left_out[19]
+ sb_5__4_/chanx_left_out[1] sb_5__4_/chanx_left_out[2] sb_5__4_/chanx_left_out[3]
+ sb_5__4_/chanx_left_out[4] sb_5__4_/chanx_left_out[5] sb_5__4_/chanx_left_out[6]
+ sb_5__4_/chanx_left_out[7] sb_5__4_/chanx_left_out[8] sb_5__4_/chanx_left_out[9]
+ sb_5__4_/chanx_right_in[0] sb_5__4_/chanx_right_in[10] sb_5__4_/chanx_right_in[11]
+ sb_5__4_/chanx_right_in[12] sb_5__4_/chanx_right_in[13] sb_5__4_/chanx_right_in[14]
+ sb_5__4_/chanx_right_in[15] sb_5__4_/chanx_right_in[16] sb_5__4_/chanx_right_in[17]
+ sb_5__4_/chanx_right_in[18] sb_5__4_/chanx_right_in[19] sb_5__4_/chanx_right_in[1]
+ sb_5__4_/chanx_right_in[2] sb_5__4_/chanx_right_in[3] sb_5__4_/chanx_right_in[4]
+ sb_5__4_/chanx_right_in[5] sb_5__4_/chanx_right_in[6] sb_5__4_/chanx_right_in[7]
+ sb_5__4_/chanx_right_in[8] sb_5__4_/chanx_right_in[9] cbx_6__4_/chanx_left_in[0]
+ cbx_6__4_/chanx_left_in[10] cbx_6__4_/chanx_left_in[11] cbx_6__4_/chanx_left_in[12]
+ cbx_6__4_/chanx_left_in[13] cbx_6__4_/chanx_left_in[14] cbx_6__4_/chanx_left_in[15]
+ cbx_6__4_/chanx_left_in[16] cbx_6__4_/chanx_left_in[17] cbx_6__4_/chanx_left_in[18]
+ cbx_6__4_/chanx_left_in[19] cbx_6__4_/chanx_left_in[1] cbx_6__4_/chanx_left_in[2]
+ cbx_6__4_/chanx_left_in[3] cbx_6__4_/chanx_left_in[4] cbx_6__4_/chanx_left_in[5]
+ cbx_6__4_/chanx_left_in[6] cbx_6__4_/chanx_left_in[7] cbx_6__4_/chanx_left_in[8]
+ cbx_6__4_/chanx_left_in[9] cby_5__4_/chany_top_out[0] cby_5__4_/chany_top_out[10]
+ cby_5__4_/chany_top_out[11] cby_5__4_/chany_top_out[12] cby_5__4_/chany_top_out[13]
+ cby_5__4_/chany_top_out[14] cby_5__4_/chany_top_out[15] cby_5__4_/chany_top_out[16]
+ cby_5__4_/chany_top_out[17] cby_5__4_/chany_top_out[18] cby_5__4_/chany_top_out[19]
+ cby_5__4_/chany_top_out[1] cby_5__4_/chany_top_out[2] cby_5__4_/chany_top_out[3]
+ cby_5__4_/chany_top_out[4] cby_5__4_/chany_top_out[5] cby_5__4_/chany_top_out[6]
+ cby_5__4_/chany_top_out[7] cby_5__4_/chany_top_out[8] cby_5__4_/chany_top_out[9]
+ cby_5__4_/chany_top_in[0] cby_5__4_/chany_top_in[10] cby_5__4_/chany_top_in[11]
+ cby_5__4_/chany_top_in[12] cby_5__4_/chany_top_in[13] cby_5__4_/chany_top_in[14]
+ cby_5__4_/chany_top_in[15] cby_5__4_/chany_top_in[16] cby_5__4_/chany_top_in[17]
+ cby_5__4_/chany_top_in[18] cby_5__4_/chany_top_in[19] cby_5__4_/chany_top_in[1]
+ cby_5__4_/chany_top_in[2] cby_5__4_/chany_top_in[3] cby_5__4_/chany_top_in[4] cby_5__4_/chany_top_in[5]
+ cby_5__4_/chany_top_in[6] cby_5__4_/chany_top_in[7] cby_5__4_/chany_top_in[8] cby_5__4_/chany_top_in[9]
+ sb_5__4_/chany_top_in[0] sb_5__4_/chany_top_in[10] sb_5__4_/chany_top_in[11] sb_5__4_/chany_top_in[12]
+ sb_5__4_/chany_top_in[13] sb_5__4_/chany_top_in[14] sb_5__4_/chany_top_in[15] sb_5__4_/chany_top_in[16]
+ sb_5__4_/chany_top_in[17] sb_5__4_/chany_top_in[18] sb_5__4_/chany_top_in[19] sb_5__4_/chany_top_in[1]
+ sb_5__4_/chany_top_in[2] sb_5__4_/chany_top_in[3] sb_5__4_/chany_top_in[4] sb_5__4_/chany_top_in[5]
+ sb_5__4_/chany_top_in[6] sb_5__4_/chany_top_in[7] sb_5__4_/chany_top_in[8] sb_5__4_/chany_top_in[9]
+ sb_5__4_/chany_top_out[0] sb_5__4_/chany_top_out[10] sb_5__4_/chany_top_out[11]
+ sb_5__4_/chany_top_out[12] sb_5__4_/chany_top_out[13] sb_5__4_/chany_top_out[14]
+ sb_5__4_/chany_top_out[15] sb_5__4_/chany_top_out[16] sb_5__4_/chany_top_out[17]
+ sb_5__4_/chany_top_out[18] sb_5__4_/chany_top_out[19] sb_5__4_/chany_top_out[1]
+ sb_5__4_/chany_top_out[2] sb_5__4_/chany_top_out[3] sb_5__4_/chany_top_out[4] sb_5__4_/chany_top_out[5]
+ sb_5__4_/chany_top_out[6] sb_5__4_/chany_top_out[7] sb_5__4_/chany_top_out[8] sb_5__4_/chany_top_out[9]
+ sb_5__4_/clk_1_E_out sb_5__4_/clk_1_N_in sb_5__4_/clk_1_W_out sb_5__4_/clk_2_E_out
+ sb_5__4_/clk_2_N_in sb_5__4_/clk_2_N_out sb_5__4_/clk_2_S_out sb_5__4_/clk_2_W_out
+ sb_5__4_/clk_3_E_out sb_5__4_/clk_3_N_in sb_5__4_/clk_3_N_out sb_5__4_/clk_3_S_out
+ sb_5__4_/clk_3_W_out sb_5__4_/left_bottom_grid_pin_34_ sb_5__4_/left_bottom_grid_pin_35_
+ sb_5__4_/left_bottom_grid_pin_36_ sb_5__4_/left_bottom_grid_pin_37_ sb_5__4_/left_bottom_grid_pin_38_
+ sb_5__4_/left_bottom_grid_pin_39_ sb_5__4_/left_bottom_grid_pin_40_ sb_5__4_/left_bottom_grid_pin_41_
+ sb_5__4_/prog_clk_0_N_in sb_5__4_/prog_clk_1_E_out sb_5__4_/prog_clk_1_N_in sb_5__4_/prog_clk_1_W_out
+ sb_5__4_/prog_clk_2_E_out sb_5__4_/prog_clk_2_N_in sb_5__4_/prog_clk_2_N_out sb_5__4_/prog_clk_2_S_out
+ sb_5__4_/prog_clk_2_W_out sb_5__4_/prog_clk_3_E_out sb_5__4_/prog_clk_3_N_in sb_5__4_/prog_clk_3_N_out
+ sb_5__4_/prog_clk_3_S_out sb_5__4_/prog_clk_3_W_out sb_5__4_/right_bottom_grid_pin_34_
+ sb_5__4_/right_bottom_grid_pin_35_ sb_5__4_/right_bottom_grid_pin_36_ sb_5__4_/right_bottom_grid_pin_37_
+ sb_5__4_/right_bottom_grid_pin_38_ sb_5__4_/right_bottom_grid_pin_39_ sb_5__4_/right_bottom_grid_pin_40_
+ sb_5__4_/right_bottom_grid_pin_41_ sb_5__4_/top_left_grid_pin_42_ sb_5__4_/top_left_grid_pin_43_
+ sb_5__4_/top_left_grid_pin_44_ sb_5__4_/top_left_grid_pin_45_ sb_5__4_/top_left_grid_pin_46_
+ sb_5__4_/top_left_grid_pin_47_ sb_5__4_/top_left_grid_pin_48_ sb_5__4_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_2__1_ sb_2__1_/Test_en_N_out sb_2__1_/Test_en_S_in VGND VPWR sb_2__1_/bottom_left_grid_pin_42_
+ sb_2__1_/bottom_left_grid_pin_43_ sb_2__1_/bottom_left_grid_pin_44_ sb_2__1_/bottom_left_grid_pin_45_
+ sb_2__1_/bottom_left_grid_pin_46_ sb_2__1_/bottom_left_grid_pin_47_ sb_2__1_/bottom_left_grid_pin_48_
+ sb_2__1_/bottom_left_grid_pin_49_ sb_2__1_/ccff_head sb_2__1_/ccff_tail sb_2__1_/chanx_left_in[0]
+ sb_2__1_/chanx_left_in[10] sb_2__1_/chanx_left_in[11] sb_2__1_/chanx_left_in[12]
+ sb_2__1_/chanx_left_in[13] sb_2__1_/chanx_left_in[14] sb_2__1_/chanx_left_in[15]
+ sb_2__1_/chanx_left_in[16] sb_2__1_/chanx_left_in[17] sb_2__1_/chanx_left_in[18]
+ sb_2__1_/chanx_left_in[19] sb_2__1_/chanx_left_in[1] sb_2__1_/chanx_left_in[2] sb_2__1_/chanx_left_in[3]
+ sb_2__1_/chanx_left_in[4] sb_2__1_/chanx_left_in[5] sb_2__1_/chanx_left_in[6] sb_2__1_/chanx_left_in[7]
+ sb_2__1_/chanx_left_in[8] sb_2__1_/chanx_left_in[9] sb_2__1_/chanx_left_out[0] sb_2__1_/chanx_left_out[10]
+ sb_2__1_/chanx_left_out[11] sb_2__1_/chanx_left_out[12] sb_2__1_/chanx_left_out[13]
+ sb_2__1_/chanx_left_out[14] sb_2__1_/chanx_left_out[15] sb_2__1_/chanx_left_out[16]
+ sb_2__1_/chanx_left_out[17] sb_2__1_/chanx_left_out[18] sb_2__1_/chanx_left_out[19]
+ sb_2__1_/chanx_left_out[1] sb_2__1_/chanx_left_out[2] sb_2__1_/chanx_left_out[3]
+ sb_2__1_/chanx_left_out[4] sb_2__1_/chanx_left_out[5] sb_2__1_/chanx_left_out[6]
+ sb_2__1_/chanx_left_out[7] sb_2__1_/chanx_left_out[8] sb_2__1_/chanx_left_out[9]
+ sb_2__1_/chanx_right_in[0] sb_2__1_/chanx_right_in[10] sb_2__1_/chanx_right_in[11]
+ sb_2__1_/chanx_right_in[12] sb_2__1_/chanx_right_in[13] sb_2__1_/chanx_right_in[14]
+ sb_2__1_/chanx_right_in[15] sb_2__1_/chanx_right_in[16] sb_2__1_/chanx_right_in[17]
+ sb_2__1_/chanx_right_in[18] sb_2__1_/chanx_right_in[19] sb_2__1_/chanx_right_in[1]
+ sb_2__1_/chanx_right_in[2] sb_2__1_/chanx_right_in[3] sb_2__1_/chanx_right_in[4]
+ sb_2__1_/chanx_right_in[5] sb_2__1_/chanx_right_in[6] sb_2__1_/chanx_right_in[7]
+ sb_2__1_/chanx_right_in[8] sb_2__1_/chanx_right_in[9] cbx_3__1_/chanx_left_in[0]
+ cbx_3__1_/chanx_left_in[10] cbx_3__1_/chanx_left_in[11] cbx_3__1_/chanx_left_in[12]
+ cbx_3__1_/chanx_left_in[13] cbx_3__1_/chanx_left_in[14] cbx_3__1_/chanx_left_in[15]
+ cbx_3__1_/chanx_left_in[16] cbx_3__1_/chanx_left_in[17] cbx_3__1_/chanx_left_in[18]
+ cbx_3__1_/chanx_left_in[19] cbx_3__1_/chanx_left_in[1] cbx_3__1_/chanx_left_in[2]
+ cbx_3__1_/chanx_left_in[3] cbx_3__1_/chanx_left_in[4] cbx_3__1_/chanx_left_in[5]
+ cbx_3__1_/chanx_left_in[6] cbx_3__1_/chanx_left_in[7] cbx_3__1_/chanx_left_in[8]
+ cbx_3__1_/chanx_left_in[9] cby_2__1_/chany_top_out[0] cby_2__1_/chany_top_out[10]
+ cby_2__1_/chany_top_out[11] cby_2__1_/chany_top_out[12] cby_2__1_/chany_top_out[13]
+ cby_2__1_/chany_top_out[14] cby_2__1_/chany_top_out[15] cby_2__1_/chany_top_out[16]
+ cby_2__1_/chany_top_out[17] cby_2__1_/chany_top_out[18] cby_2__1_/chany_top_out[19]
+ cby_2__1_/chany_top_out[1] cby_2__1_/chany_top_out[2] cby_2__1_/chany_top_out[3]
+ cby_2__1_/chany_top_out[4] cby_2__1_/chany_top_out[5] cby_2__1_/chany_top_out[6]
+ cby_2__1_/chany_top_out[7] cby_2__1_/chany_top_out[8] cby_2__1_/chany_top_out[9]
+ cby_2__1_/chany_top_in[0] cby_2__1_/chany_top_in[10] cby_2__1_/chany_top_in[11]
+ cby_2__1_/chany_top_in[12] cby_2__1_/chany_top_in[13] cby_2__1_/chany_top_in[14]
+ cby_2__1_/chany_top_in[15] cby_2__1_/chany_top_in[16] cby_2__1_/chany_top_in[17]
+ cby_2__1_/chany_top_in[18] cby_2__1_/chany_top_in[19] cby_2__1_/chany_top_in[1]
+ cby_2__1_/chany_top_in[2] cby_2__1_/chany_top_in[3] cby_2__1_/chany_top_in[4] cby_2__1_/chany_top_in[5]
+ cby_2__1_/chany_top_in[6] cby_2__1_/chany_top_in[7] cby_2__1_/chany_top_in[8] cby_2__1_/chany_top_in[9]
+ sb_2__1_/chany_top_in[0] sb_2__1_/chany_top_in[10] sb_2__1_/chany_top_in[11] sb_2__1_/chany_top_in[12]
+ sb_2__1_/chany_top_in[13] sb_2__1_/chany_top_in[14] sb_2__1_/chany_top_in[15] sb_2__1_/chany_top_in[16]
+ sb_2__1_/chany_top_in[17] sb_2__1_/chany_top_in[18] sb_2__1_/chany_top_in[19] sb_2__1_/chany_top_in[1]
+ sb_2__1_/chany_top_in[2] sb_2__1_/chany_top_in[3] sb_2__1_/chany_top_in[4] sb_2__1_/chany_top_in[5]
+ sb_2__1_/chany_top_in[6] sb_2__1_/chany_top_in[7] sb_2__1_/chany_top_in[8] sb_2__1_/chany_top_in[9]
+ sb_2__1_/chany_top_out[0] sb_2__1_/chany_top_out[10] sb_2__1_/chany_top_out[11]
+ sb_2__1_/chany_top_out[12] sb_2__1_/chany_top_out[13] sb_2__1_/chany_top_out[14]
+ sb_2__1_/chany_top_out[15] sb_2__1_/chany_top_out[16] sb_2__1_/chany_top_out[17]
+ sb_2__1_/chany_top_out[18] sb_2__1_/chany_top_out[19] sb_2__1_/chany_top_out[1]
+ sb_2__1_/chany_top_out[2] sb_2__1_/chany_top_out[3] sb_2__1_/chany_top_out[4] sb_2__1_/chany_top_out[5]
+ sb_2__1_/chany_top_out[6] sb_2__1_/chany_top_out[7] sb_2__1_/chany_top_out[8] sb_2__1_/chany_top_out[9]
+ sb_2__1_/clk_1_E_out sb_2__1_/clk_1_N_in sb_2__1_/clk_1_W_out sb_2__1_/clk_2_E_out
+ sb_2__1_/clk_2_N_in sb_2__1_/clk_2_N_out sb_2__1_/clk_2_S_out sb_2__1_/clk_2_W_out
+ sb_2__1_/clk_3_E_out sb_2__1_/clk_3_N_in sb_2__1_/clk_3_N_out sb_2__1_/clk_3_S_out
+ sb_2__1_/clk_3_W_out sb_2__1_/left_bottom_grid_pin_34_ sb_2__1_/left_bottom_grid_pin_35_
+ sb_2__1_/left_bottom_grid_pin_36_ sb_2__1_/left_bottom_grid_pin_37_ sb_2__1_/left_bottom_grid_pin_38_
+ sb_2__1_/left_bottom_grid_pin_39_ sb_2__1_/left_bottom_grid_pin_40_ sb_2__1_/left_bottom_grid_pin_41_
+ sb_2__1_/prog_clk_0_N_in sb_2__1_/prog_clk_1_E_out sb_2__1_/prog_clk_1_N_in sb_2__1_/prog_clk_1_W_out
+ sb_2__1_/prog_clk_2_E_out sb_2__1_/prog_clk_2_N_in sb_2__1_/prog_clk_2_N_out sb_2__1_/prog_clk_2_S_out
+ sb_2__1_/prog_clk_2_W_out sb_2__1_/prog_clk_3_E_out sb_2__1_/prog_clk_3_N_in sb_2__1_/prog_clk_3_N_out
+ sb_2__1_/prog_clk_3_S_out sb_2__1_/prog_clk_3_W_out sb_2__1_/right_bottom_grid_pin_34_
+ sb_2__1_/right_bottom_grid_pin_35_ sb_2__1_/right_bottom_grid_pin_36_ sb_2__1_/right_bottom_grid_pin_37_
+ sb_2__1_/right_bottom_grid_pin_38_ sb_2__1_/right_bottom_grid_pin_39_ sb_2__1_/right_bottom_grid_pin_40_
+ sb_2__1_/right_bottom_grid_pin_41_ sb_2__1_/top_left_grid_pin_42_ sb_2__1_/top_left_grid_pin_43_
+ sb_2__1_/top_left_grid_pin_44_ sb_2__1_/top_left_grid_pin_45_ sb_2__1_/top_left_grid_pin_46_
+ sb_2__1_/top_left_grid_pin_47_ sb_2__1_/top_left_grid_pin_48_ sb_2__1_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_4__8_ sb_4__7_/Test_en_N_out cby_4__8_/Test_en_E_out cby_4__8_/Test_en_N_out
+ sb_4__7_/Test_en_N_out sb_4__7_/Test_en_N_out cby_4__8_/Test_en_W_out VGND VPWR
+ cby_4__8_/ccff_head cby_4__8_/ccff_tail sb_4__7_/chany_top_out[0] sb_4__7_/chany_top_out[10]
+ sb_4__7_/chany_top_out[11] sb_4__7_/chany_top_out[12] sb_4__7_/chany_top_out[13]
+ sb_4__7_/chany_top_out[14] sb_4__7_/chany_top_out[15] sb_4__7_/chany_top_out[16]
+ sb_4__7_/chany_top_out[17] sb_4__7_/chany_top_out[18] sb_4__7_/chany_top_out[19]
+ sb_4__7_/chany_top_out[1] sb_4__7_/chany_top_out[2] sb_4__7_/chany_top_out[3] sb_4__7_/chany_top_out[4]
+ sb_4__7_/chany_top_out[5] sb_4__7_/chany_top_out[6] sb_4__7_/chany_top_out[7] sb_4__7_/chany_top_out[8]
+ sb_4__7_/chany_top_out[9] sb_4__7_/chany_top_in[0] sb_4__7_/chany_top_in[10] sb_4__7_/chany_top_in[11]
+ sb_4__7_/chany_top_in[12] sb_4__7_/chany_top_in[13] sb_4__7_/chany_top_in[14] sb_4__7_/chany_top_in[15]
+ sb_4__7_/chany_top_in[16] sb_4__7_/chany_top_in[17] sb_4__7_/chany_top_in[18] sb_4__7_/chany_top_in[19]
+ sb_4__7_/chany_top_in[1] sb_4__7_/chany_top_in[2] sb_4__7_/chany_top_in[3] sb_4__7_/chany_top_in[4]
+ sb_4__7_/chany_top_in[5] sb_4__7_/chany_top_in[6] sb_4__7_/chany_top_in[7] sb_4__7_/chany_top_in[8]
+ sb_4__7_/chany_top_in[9] cby_4__8_/chany_top_in[0] cby_4__8_/chany_top_in[10] cby_4__8_/chany_top_in[11]
+ cby_4__8_/chany_top_in[12] cby_4__8_/chany_top_in[13] cby_4__8_/chany_top_in[14]
+ cby_4__8_/chany_top_in[15] cby_4__8_/chany_top_in[16] cby_4__8_/chany_top_in[17]
+ cby_4__8_/chany_top_in[18] cby_4__8_/chany_top_in[19] cby_4__8_/chany_top_in[1]
+ cby_4__8_/chany_top_in[2] cby_4__8_/chany_top_in[3] cby_4__8_/chany_top_in[4] cby_4__8_/chany_top_in[5]
+ cby_4__8_/chany_top_in[6] cby_4__8_/chany_top_in[7] cby_4__8_/chany_top_in[8] cby_4__8_/chany_top_in[9]
+ cby_4__8_/chany_top_out[0] cby_4__8_/chany_top_out[10] cby_4__8_/chany_top_out[11]
+ cby_4__8_/chany_top_out[12] cby_4__8_/chany_top_out[13] cby_4__8_/chany_top_out[14]
+ cby_4__8_/chany_top_out[15] cby_4__8_/chany_top_out[16] cby_4__8_/chany_top_out[17]
+ cby_4__8_/chany_top_out[18] cby_4__8_/chany_top_out[19] cby_4__8_/chany_top_out[1]
+ cby_4__8_/chany_top_out[2] cby_4__8_/chany_top_out[3] cby_4__8_/chany_top_out[4]
+ cby_4__8_/chany_top_out[5] cby_4__8_/chany_top_out[6] cby_4__8_/chany_top_out[7]
+ cby_4__8_/chany_top_out[8] cby_4__8_/chany_top_out[9] cby_4__8_/clk_2_N_out cby_4__8_/clk_2_S_in
+ cby_4__8_/clk_2_S_out cby_4__8_/clk_3_N_out cby_4__8_/clk_3_S_in cby_4__8_/clk_3_S_out
+ cby_4__8_/left_grid_pin_16_ cby_4__8_/left_grid_pin_17_ cby_4__8_/left_grid_pin_18_
+ cby_4__8_/left_grid_pin_19_ cby_4__8_/left_grid_pin_20_ cby_4__8_/left_grid_pin_21_
+ cby_4__8_/left_grid_pin_22_ cby_4__8_/left_grid_pin_23_ cby_4__8_/left_grid_pin_24_
+ cby_4__8_/left_grid_pin_25_ cby_4__8_/left_grid_pin_26_ cby_4__8_/left_grid_pin_27_
+ cby_4__8_/left_grid_pin_28_ cby_4__8_/left_grid_pin_29_ cby_4__8_/left_grid_pin_30_
+ cby_4__8_/left_grid_pin_31_ sb_4__8_/prog_clk_0_S_in sb_4__7_/prog_clk_0_N_in cby_4__8_/prog_clk_0_W_in
+ cby_4__8_/prog_clk_2_N_out cby_4__8_/prog_clk_2_S_in cby_4__8_/prog_clk_2_S_out
+ cby_4__8_/prog_clk_3_N_out cby_4__8_/prog_clk_3_S_in cby_4__8_/prog_clk_3_S_out
+ cby_1__1_
Xcby_1__5_ cby_1__5_/Test_en_W_in cby_1__5_/Test_en_E_out cby_1__5_/Test_en_N_out
+ cby_1__5_/Test_en_W_in cby_1__5_/Test_en_W_in cby_1__5_/Test_en_W_out VGND VPWR
+ cby_1__5_/ccff_head cby_1__5_/ccff_tail sb_1__4_/chany_top_out[0] sb_1__4_/chany_top_out[10]
+ sb_1__4_/chany_top_out[11] sb_1__4_/chany_top_out[12] sb_1__4_/chany_top_out[13]
+ sb_1__4_/chany_top_out[14] sb_1__4_/chany_top_out[15] sb_1__4_/chany_top_out[16]
+ sb_1__4_/chany_top_out[17] sb_1__4_/chany_top_out[18] sb_1__4_/chany_top_out[19]
+ sb_1__4_/chany_top_out[1] sb_1__4_/chany_top_out[2] sb_1__4_/chany_top_out[3] sb_1__4_/chany_top_out[4]
+ sb_1__4_/chany_top_out[5] sb_1__4_/chany_top_out[6] sb_1__4_/chany_top_out[7] sb_1__4_/chany_top_out[8]
+ sb_1__4_/chany_top_out[9] sb_1__4_/chany_top_in[0] sb_1__4_/chany_top_in[10] sb_1__4_/chany_top_in[11]
+ sb_1__4_/chany_top_in[12] sb_1__4_/chany_top_in[13] sb_1__4_/chany_top_in[14] sb_1__4_/chany_top_in[15]
+ sb_1__4_/chany_top_in[16] sb_1__4_/chany_top_in[17] sb_1__4_/chany_top_in[18] sb_1__4_/chany_top_in[19]
+ sb_1__4_/chany_top_in[1] sb_1__4_/chany_top_in[2] sb_1__4_/chany_top_in[3] sb_1__4_/chany_top_in[4]
+ sb_1__4_/chany_top_in[5] sb_1__4_/chany_top_in[6] sb_1__4_/chany_top_in[7] sb_1__4_/chany_top_in[8]
+ sb_1__4_/chany_top_in[9] cby_1__5_/chany_top_in[0] cby_1__5_/chany_top_in[10] cby_1__5_/chany_top_in[11]
+ cby_1__5_/chany_top_in[12] cby_1__5_/chany_top_in[13] cby_1__5_/chany_top_in[14]
+ cby_1__5_/chany_top_in[15] cby_1__5_/chany_top_in[16] cby_1__5_/chany_top_in[17]
+ cby_1__5_/chany_top_in[18] cby_1__5_/chany_top_in[19] cby_1__5_/chany_top_in[1]
+ cby_1__5_/chany_top_in[2] cby_1__5_/chany_top_in[3] cby_1__5_/chany_top_in[4] cby_1__5_/chany_top_in[5]
+ cby_1__5_/chany_top_in[6] cby_1__5_/chany_top_in[7] cby_1__5_/chany_top_in[8] cby_1__5_/chany_top_in[9]
+ cby_1__5_/chany_top_out[0] cby_1__5_/chany_top_out[10] cby_1__5_/chany_top_out[11]
+ cby_1__5_/chany_top_out[12] cby_1__5_/chany_top_out[13] cby_1__5_/chany_top_out[14]
+ cby_1__5_/chany_top_out[15] cby_1__5_/chany_top_out[16] cby_1__5_/chany_top_out[17]
+ cby_1__5_/chany_top_out[18] cby_1__5_/chany_top_out[19] cby_1__5_/chany_top_out[1]
+ cby_1__5_/chany_top_out[2] cby_1__5_/chany_top_out[3] cby_1__5_/chany_top_out[4]
+ cby_1__5_/chany_top_out[5] cby_1__5_/chany_top_out[6] cby_1__5_/chany_top_out[7]
+ cby_1__5_/chany_top_out[8] cby_1__5_/chany_top_out[9] cby_1__5_/clk_2_N_out cby_1__5_/clk_2_S_in
+ cby_1__5_/clk_2_S_out cby_1__5_/clk_3_N_out cby_1__5_/clk_3_S_in cby_1__5_/clk_3_S_out
+ cby_1__5_/left_grid_pin_16_ cby_1__5_/left_grid_pin_17_ cby_1__5_/left_grid_pin_18_
+ cby_1__5_/left_grid_pin_19_ cby_1__5_/left_grid_pin_20_ cby_1__5_/left_grid_pin_21_
+ cby_1__5_/left_grid_pin_22_ cby_1__5_/left_grid_pin_23_ cby_1__5_/left_grid_pin_24_
+ cby_1__5_/left_grid_pin_25_ cby_1__5_/left_grid_pin_26_ cby_1__5_/left_grid_pin_27_
+ cby_1__5_/left_grid_pin_28_ cby_1__5_/left_grid_pin_29_ cby_1__5_/left_grid_pin_30_
+ cby_1__5_/left_grid_pin_31_ cby_1__5_/prog_clk_0_N_out sb_1__4_/prog_clk_0_N_in
+ cby_1__5_/prog_clk_0_W_in cby_1__5_/prog_clk_2_N_out cby_1__5_/prog_clk_2_S_in cby_1__5_/prog_clk_2_S_out
+ cby_1__5_/prog_clk_3_N_out cby_1__5_/prog_clk_3_S_in cby_1__5_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_8__1_ cbx_8__1_/REGIN_FEEDTHROUGH cbx_8__1_/REGOUT_FEEDTHROUGH cbx_8__1_/SC_IN_BOT
+ cbx_8__1_/SC_IN_TOP cbx_8__1_/SC_OUT_BOT cbx_8__1_/SC_OUT_TOP VGND VPWR cbx_8__1_/bottom_grid_pin_0_
+ cbx_8__1_/bottom_grid_pin_10_ cbx_8__1_/bottom_grid_pin_11_ cbx_8__1_/bottom_grid_pin_12_
+ cbx_8__1_/bottom_grid_pin_13_ cbx_8__1_/bottom_grid_pin_14_ cbx_8__1_/bottom_grid_pin_15_
+ cbx_8__1_/bottom_grid_pin_1_ cbx_8__1_/bottom_grid_pin_2_ cbx_8__1_/bottom_grid_pin_3_
+ cbx_8__1_/bottom_grid_pin_4_ cbx_8__1_/bottom_grid_pin_5_ cbx_8__1_/bottom_grid_pin_6_
+ cbx_8__1_/bottom_grid_pin_7_ cbx_8__1_/bottom_grid_pin_8_ cbx_8__1_/bottom_grid_pin_9_
+ sb_8__1_/ccff_tail sb_7__1_/ccff_head cbx_8__1_/chanx_left_in[0] cbx_8__1_/chanx_left_in[10]
+ cbx_8__1_/chanx_left_in[11] cbx_8__1_/chanx_left_in[12] cbx_8__1_/chanx_left_in[13]
+ cbx_8__1_/chanx_left_in[14] cbx_8__1_/chanx_left_in[15] cbx_8__1_/chanx_left_in[16]
+ cbx_8__1_/chanx_left_in[17] cbx_8__1_/chanx_left_in[18] cbx_8__1_/chanx_left_in[19]
+ cbx_8__1_/chanx_left_in[1] cbx_8__1_/chanx_left_in[2] cbx_8__1_/chanx_left_in[3]
+ cbx_8__1_/chanx_left_in[4] cbx_8__1_/chanx_left_in[5] cbx_8__1_/chanx_left_in[6]
+ cbx_8__1_/chanx_left_in[7] cbx_8__1_/chanx_left_in[8] cbx_8__1_/chanx_left_in[9]
+ sb_7__1_/chanx_right_in[0] sb_7__1_/chanx_right_in[10] sb_7__1_/chanx_right_in[11]
+ sb_7__1_/chanx_right_in[12] sb_7__1_/chanx_right_in[13] sb_7__1_/chanx_right_in[14]
+ sb_7__1_/chanx_right_in[15] sb_7__1_/chanx_right_in[16] sb_7__1_/chanx_right_in[17]
+ sb_7__1_/chanx_right_in[18] sb_7__1_/chanx_right_in[19] sb_7__1_/chanx_right_in[1]
+ sb_7__1_/chanx_right_in[2] sb_7__1_/chanx_right_in[3] sb_7__1_/chanx_right_in[4]
+ sb_7__1_/chanx_right_in[5] sb_7__1_/chanx_right_in[6] sb_7__1_/chanx_right_in[7]
+ sb_7__1_/chanx_right_in[8] sb_7__1_/chanx_right_in[9] sb_8__1_/chanx_left_out[0]
+ sb_8__1_/chanx_left_out[10] sb_8__1_/chanx_left_out[11] sb_8__1_/chanx_left_out[12]
+ sb_8__1_/chanx_left_out[13] sb_8__1_/chanx_left_out[14] sb_8__1_/chanx_left_out[15]
+ sb_8__1_/chanx_left_out[16] sb_8__1_/chanx_left_out[17] sb_8__1_/chanx_left_out[18]
+ sb_8__1_/chanx_left_out[19] sb_8__1_/chanx_left_out[1] sb_8__1_/chanx_left_out[2]
+ sb_8__1_/chanx_left_out[3] sb_8__1_/chanx_left_out[4] sb_8__1_/chanx_left_out[5]
+ sb_8__1_/chanx_left_out[6] sb_8__1_/chanx_left_out[7] sb_8__1_/chanx_left_out[8]
+ sb_8__1_/chanx_left_out[9] sb_8__1_/chanx_left_in[0] sb_8__1_/chanx_left_in[10]
+ sb_8__1_/chanx_left_in[11] sb_8__1_/chanx_left_in[12] sb_8__1_/chanx_left_in[13]
+ sb_8__1_/chanx_left_in[14] sb_8__1_/chanx_left_in[15] sb_8__1_/chanx_left_in[16]
+ sb_8__1_/chanx_left_in[17] sb_8__1_/chanx_left_in[18] sb_8__1_/chanx_left_in[19]
+ sb_8__1_/chanx_left_in[1] sb_8__1_/chanx_left_in[2] sb_8__1_/chanx_left_in[3] sb_8__1_/chanx_left_in[4]
+ sb_8__1_/chanx_left_in[5] sb_8__1_/chanx_left_in[6] sb_8__1_/chanx_left_in[7] sb_8__1_/chanx_left_in[8]
+ sb_8__1_/chanx_left_in[9] cbx_8__1_/clk_1_N_out cbx_8__1_/clk_1_S_out sb_7__1_/clk_1_E_out
+ cbx_8__1_/clk_2_E_out cbx_8__1_/clk_2_W_in cbx_8__1_/clk_2_W_out cbx_8__1_/clk_3_E_out
+ cbx_8__1_/clk_3_W_in cbx_8__1_/clk_3_W_out cbx_8__1_/prog_clk_0_N_in cbx_8__1_/prog_clk_0_W_out
+ cbx_8__1_/prog_clk_1_N_out cbx_8__1_/prog_clk_1_S_out sb_7__1_/prog_clk_1_E_out
+ cbx_8__1_/prog_clk_2_E_out cbx_8__1_/prog_clk_2_W_in cbx_8__1_/prog_clk_2_W_out
+ cbx_8__1_/prog_clk_3_E_out cbx_8__1_/prog_clk_3_W_in cbx_8__1_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_8__6_ VGND VPWR sb_8__6_/bottom_left_grid_pin_42_ sb_8__6_/bottom_left_grid_pin_43_
+ sb_8__6_/bottom_left_grid_pin_44_ sb_8__6_/bottom_left_grid_pin_45_ sb_8__6_/bottom_left_grid_pin_46_
+ sb_8__6_/bottom_left_grid_pin_47_ sb_8__6_/bottom_left_grid_pin_48_ sb_8__6_/bottom_left_grid_pin_49_
+ sb_8__6_/bottom_right_grid_pin_1_ sb_8__6_/ccff_head sb_8__6_/ccff_tail sb_8__6_/chanx_left_in[0]
+ sb_8__6_/chanx_left_in[10] sb_8__6_/chanx_left_in[11] sb_8__6_/chanx_left_in[12]
+ sb_8__6_/chanx_left_in[13] sb_8__6_/chanx_left_in[14] sb_8__6_/chanx_left_in[15]
+ sb_8__6_/chanx_left_in[16] sb_8__6_/chanx_left_in[17] sb_8__6_/chanx_left_in[18]
+ sb_8__6_/chanx_left_in[19] sb_8__6_/chanx_left_in[1] sb_8__6_/chanx_left_in[2] sb_8__6_/chanx_left_in[3]
+ sb_8__6_/chanx_left_in[4] sb_8__6_/chanx_left_in[5] sb_8__6_/chanx_left_in[6] sb_8__6_/chanx_left_in[7]
+ sb_8__6_/chanx_left_in[8] sb_8__6_/chanx_left_in[9] sb_8__6_/chanx_left_out[0] sb_8__6_/chanx_left_out[10]
+ sb_8__6_/chanx_left_out[11] sb_8__6_/chanx_left_out[12] sb_8__6_/chanx_left_out[13]
+ sb_8__6_/chanx_left_out[14] sb_8__6_/chanx_left_out[15] sb_8__6_/chanx_left_out[16]
+ sb_8__6_/chanx_left_out[17] sb_8__6_/chanx_left_out[18] sb_8__6_/chanx_left_out[19]
+ sb_8__6_/chanx_left_out[1] sb_8__6_/chanx_left_out[2] sb_8__6_/chanx_left_out[3]
+ sb_8__6_/chanx_left_out[4] sb_8__6_/chanx_left_out[5] sb_8__6_/chanx_left_out[6]
+ sb_8__6_/chanx_left_out[7] sb_8__6_/chanx_left_out[8] sb_8__6_/chanx_left_out[9]
+ cby_8__6_/chany_top_out[0] cby_8__6_/chany_top_out[10] cby_8__6_/chany_top_out[11]
+ cby_8__6_/chany_top_out[12] cby_8__6_/chany_top_out[13] cby_8__6_/chany_top_out[14]
+ cby_8__6_/chany_top_out[15] cby_8__6_/chany_top_out[16] cby_8__6_/chany_top_out[17]
+ cby_8__6_/chany_top_out[18] cby_8__6_/chany_top_out[19] cby_8__6_/chany_top_out[1]
+ cby_8__6_/chany_top_out[2] cby_8__6_/chany_top_out[3] cby_8__6_/chany_top_out[4]
+ cby_8__6_/chany_top_out[5] cby_8__6_/chany_top_out[6] cby_8__6_/chany_top_out[7]
+ cby_8__6_/chany_top_out[8] cby_8__6_/chany_top_out[9] cby_8__6_/chany_top_in[0]
+ cby_8__6_/chany_top_in[10] cby_8__6_/chany_top_in[11] cby_8__6_/chany_top_in[12]
+ cby_8__6_/chany_top_in[13] cby_8__6_/chany_top_in[14] cby_8__6_/chany_top_in[15]
+ cby_8__6_/chany_top_in[16] cby_8__6_/chany_top_in[17] cby_8__6_/chany_top_in[18]
+ cby_8__6_/chany_top_in[19] cby_8__6_/chany_top_in[1] cby_8__6_/chany_top_in[2] cby_8__6_/chany_top_in[3]
+ cby_8__6_/chany_top_in[4] cby_8__6_/chany_top_in[5] cby_8__6_/chany_top_in[6] cby_8__6_/chany_top_in[7]
+ cby_8__6_/chany_top_in[8] cby_8__6_/chany_top_in[9] sb_8__6_/chany_top_in[0] sb_8__6_/chany_top_in[10]
+ sb_8__6_/chany_top_in[11] sb_8__6_/chany_top_in[12] sb_8__6_/chany_top_in[13] sb_8__6_/chany_top_in[14]
+ sb_8__6_/chany_top_in[15] sb_8__6_/chany_top_in[16] sb_8__6_/chany_top_in[17] sb_8__6_/chany_top_in[18]
+ sb_8__6_/chany_top_in[19] sb_8__6_/chany_top_in[1] sb_8__6_/chany_top_in[2] sb_8__6_/chany_top_in[3]
+ sb_8__6_/chany_top_in[4] sb_8__6_/chany_top_in[5] sb_8__6_/chany_top_in[6] sb_8__6_/chany_top_in[7]
+ sb_8__6_/chany_top_in[8] sb_8__6_/chany_top_in[9] sb_8__6_/chany_top_out[0] sb_8__6_/chany_top_out[10]
+ sb_8__6_/chany_top_out[11] sb_8__6_/chany_top_out[12] sb_8__6_/chany_top_out[13]
+ sb_8__6_/chany_top_out[14] sb_8__6_/chany_top_out[15] sb_8__6_/chany_top_out[16]
+ sb_8__6_/chany_top_out[17] sb_8__6_/chany_top_out[18] sb_8__6_/chany_top_out[19]
+ sb_8__6_/chany_top_out[1] sb_8__6_/chany_top_out[2] sb_8__6_/chany_top_out[3] sb_8__6_/chany_top_out[4]
+ sb_8__6_/chany_top_out[5] sb_8__6_/chany_top_out[6] sb_8__6_/chany_top_out[7] sb_8__6_/chany_top_out[8]
+ sb_8__6_/chany_top_out[9] sb_8__6_/left_bottom_grid_pin_34_ sb_8__6_/left_bottom_grid_pin_35_
+ sb_8__6_/left_bottom_grid_pin_36_ sb_8__6_/left_bottom_grid_pin_37_ sb_8__6_/left_bottom_grid_pin_38_
+ sb_8__6_/left_bottom_grid_pin_39_ sb_8__6_/left_bottom_grid_pin_40_ sb_8__6_/left_bottom_grid_pin_41_
+ sb_8__6_/prog_clk_0_N_in sb_8__6_/top_left_grid_pin_42_ sb_8__6_/top_left_grid_pin_43_
+ sb_8__6_/top_left_grid_pin_44_ sb_8__6_/top_left_grid_pin_45_ sb_8__6_/top_left_grid_pin_46_
+ sb_8__6_/top_left_grid_pin_47_ sb_8__6_/top_left_grid_pin_48_ sb_8__6_/top_left_grid_pin_49_
+ sb_8__6_/top_right_grid_pin_1_ sb_2__1_
Xcbx_1__6_ cbx_1__6_/REGIN_FEEDTHROUGH cbx_1__6_/REGOUT_FEEDTHROUGH cbx_1__6_/SC_IN_BOT
+ cbx_1__6_/SC_IN_TOP cbx_1__6_/SC_OUT_BOT cbx_1__6_/SC_OUT_TOP VGND VPWR cbx_1__6_/bottom_grid_pin_0_
+ cbx_1__6_/bottom_grid_pin_10_ cbx_1__6_/bottom_grid_pin_11_ cbx_1__6_/bottom_grid_pin_12_
+ cbx_1__6_/bottom_grid_pin_13_ cbx_1__6_/bottom_grid_pin_14_ cbx_1__6_/bottom_grid_pin_15_
+ cbx_1__6_/bottom_grid_pin_1_ cbx_1__6_/bottom_grid_pin_2_ cbx_1__6_/bottom_grid_pin_3_
+ cbx_1__6_/bottom_grid_pin_4_ cbx_1__6_/bottom_grid_pin_5_ cbx_1__6_/bottom_grid_pin_6_
+ cbx_1__6_/bottom_grid_pin_7_ cbx_1__6_/bottom_grid_pin_8_ cbx_1__6_/bottom_grid_pin_9_
+ sb_1__6_/ccff_tail sb_0__6_/ccff_head cbx_1__6_/chanx_left_in[0] cbx_1__6_/chanx_left_in[10]
+ cbx_1__6_/chanx_left_in[11] cbx_1__6_/chanx_left_in[12] cbx_1__6_/chanx_left_in[13]
+ cbx_1__6_/chanx_left_in[14] cbx_1__6_/chanx_left_in[15] cbx_1__6_/chanx_left_in[16]
+ cbx_1__6_/chanx_left_in[17] cbx_1__6_/chanx_left_in[18] cbx_1__6_/chanx_left_in[19]
+ cbx_1__6_/chanx_left_in[1] cbx_1__6_/chanx_left_in[2] cbx_1__6_/chanx_left_in[3]
+ cbx_1__6_/chanx_left_in[4] cbx_1__6_/chanx_left_in[5] cbx_1__6_/chanx_left_in[6]
+ cbx_1__6_/chanx_left_in[7] cbx_1__6_/chanx_left_in[8] cbx_1__6_/chanx_left_in[9]
+ sb_0__6_/chanx_right_in[0] sb_0__6_/chanx_right_in[10] sb_0__6_/chanx_right_in[11]
+ sb_0__6_/chanx_right_in[12] sb_0__6_/chanx_right_in[13] sb_0__6_/chanx_right_in[14]
+ sb_0__6_/chanx_right_in[15] sb_0__6_/chanx_right_in[16] sb_0__6_/chanx_right_in[17]
+ sb_0__6_/chanx_right_in[18] sb_0__6_/chanx_right_in[19] sb_0__6_/chanx_right_in[1]
+ sb_0__6_/chanx_right_in[2] sb_0__6_/chanx_right_in[3] sb_0__6_/chanx_right_in[4]
+ sb_0__6_/chanx_right_in[5] sb_0__6_/chanx_right_in[6] sb_0__6_/chanx_right_in[7]
+ sb_0__6_/chanx_right_in[8] sb_0__6_/chanx_right_in[9] sb_1__6_/chanx_left_out[0]
+ sb_1__6_/chanx_left_out[10] sb_1__6_/chanx_left_out[11] sb_1__6_/chanx_left_out[12]
+ sb_1__6_/chanx_left_out[13] sb_1__6_/chanx_left_out[14] sb_1__6_/chanx_left_out[15]
+ sb_1__6_/chanx_left_out[16] sb_1__6_/chanx_left_out[17] sb_1__6_/chanx_left_out[18]
+ sb_1__6_/chanx_left_out[19] sb_1__6_/chanx_left_out[1] sb_1__6_/chanx_left_out[2]
+ sb_1__6_/chanx_left_out[3] sb_1__6_/chanx_left_out[4] sb_1__6_/chanx_left_out[5]
+ sb_1__6_/chanx_left_out[6] sb_1__6_/chanx_left_out[7] sb_1__6_/chanx_left_out[8]
+ sb_1__6_/chanx_left_out[9] sb_1__6_/chanx_left_in[0] sb_1__6_/chanx_left_in[10]
+ sb_1__6_/chanx_left_in[11] sb_1__6_/chanx_left_in[12] sb_1__6_/chanx_left_in[13]
+ sb_1__6_/chanx_left_in[14] sb_1__6_/chanx_left_in[15] sb_1__6_/chanx_left_in[16]
+ sb_1__6_/chanx_left_in[17] sb_1__6_/chanx_left_in[18] sb_1__6_/chanx_left_in[19]
+ sb_1__6_/chanx_left_in[1] sb_1__6_/chanx_left_in[2] sb_1__6_/chanx_left_in[3] sb_1__6_/chanx_left_in[4]
+ sb_1__6_/chanx_left_in[5] sb_1__6_/chanx_left_in[6] sb_1__6_/chanx_left_in[7] sb_1__6_/chanx_left_in[8]
+ sb_1__6_/chanx_left_in[9] cbx_1__6_/clk_1_N_out cbx_1__6_/clk_1_S_out cbx_1__6_/clk_1_W_in
+ cbx_1__6_/clk_2_E_out cbx_1__6_/clk_2_W_in cbx_1__6_/clk_2_W_out cbx_1__6_/clk_3_E_out
+ cbx_1__6_/clk_3_W_in cbx_1__6_/clk_3_W_out cbx_1__6_/prog_clk_0_N_in sb_0__6_/prog_clk_0_E_in
+ cbx_1__6_/prog_clk_1_N_out cbx_1__6_/prog_clk_1_S_out cbx_1__6_/prog_clk_1_W_in
+ cbx_1__6_/prog_clk_2_E_out cbx_1__6_/prog_clk_2_W_in cbx_1__6_/prog_clk_2_W_out
+ cbx_1__6_/prog_clk_3_E_out cbx_1__6_/prog_clk_3_W_in cbx_1__6_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_5__3_ sb_5__3_/Test_en_N_out sb_5__3_/Test_en_S_in VGND VPWR sb_5__3_/bottom_left_grid_pin_42_
+ sb_5__3_/bottom_left_grid_pin_43_ sb_5__3_/bottom_left_grid_pin_44_ sb_5__3_/bottom_left_grid_pin_45_
+ sb_5__3_/bottom_left_grid_pin_46_ sb_5__3_/bottom_left_grid_pin_47_ sb_5__3_/bottom_left_grid_pin_48_
+ sb_5__3_/bottom_left_grid_pin_49_ sb_5__3_/ccff_head sb_5__3_/ccff_tail sb_5__3_/chanx_left_in[0]
+ sb_5__3_/chanx_left_in[10] sb_5__3_/chanx_left_in[11] sb_5__3_/chanx_left_in[12]
+ sb_5__3_/chanx_left_in[13] sb_5__3_/chanx_left_in[14] sb_5__3_/chanx_left_in[15]
+ sb_5__3_/chanx_left_in[16] sb_5__3_/chanx_left_in[17] sb_5__3_/chanx_left_in[18]
+ sb_5__3_/chanx_left_in[19] sb_5__3_/chanx_left_in[1] sb_5__3_/chanx_left_in[2] sb_5__3_/chanx_left_in[3]
+ sb_5__3_/chanx_left_in[4] sb_5__3_/chanx_left_in[5] sb_5__3_/chanx_left_in[6] sb_5__3_/chanx_left_in[7]
+ sb_5__3_/chanx_left_in[8] sb_5__3_/chanx_left_in[9] sb_5__3_/chanx_left_out[0] sb_5__3_/chanx_left_out[10]
+ sb_5__3_/chanx_left_out[11] sb_5__3_/chanx_left_out[12] sb_5__3_/chanx_left_out[13]
+ sb_5__3_/chanx_left_out[14] sb_5__3_/chanx_left_out[15] sb_5__3_/chanx_left_out[16]
+ sb_5__3_/chanx_left_out[17] sb_5__3_/chanx_left_out[18] sb_5__3_/chanx_left_out[19]
+ sb_5__3_/chanx_left_out[1] sb_5__3_/chanx_left_out[2] sb_5__3_/chanx_left_out[3]
+ sb_5__3_/chanx_left_out[4] sb_5__3_/chanx_left_out[5] sb_5__3_/chanx_left_out[6]
+ sb_5__3_/chanx_left_out[7] sb_5__3_/chanx_left_out[8] sb_5__3_/chanx_left_out[9]
+ sb_5__3_/chanx_right_in[0] sb_5__3_/chanx_right_in[10] sb_5__3_/chanx_right_in[11]
+ sb_5__3_/chanx_right_in[12] sb_5__3_/chanx_right_in[13] sb_5__3_/chanx_right_in[14]
+ sb_5__3_/chanx_right_in[15] sb_5__3_/chanx_right_in[16] sb_5__3_/chanx_right_in[17]
+ sb_5__3_/chanx_right_in[18] sb_5__3_/chanx_right_in[19] sb_5__3_/chanx_right_in[1]
+ sb_5__3_/chanx_right_in[2] sb_5__3_/chanx_right_in[3] sb_5__3_/chanx_right_in[4]
+ sb_5__3_/chanx_right_in[5] sb_5__3_/chanx_right_in[6] sb_5__3_/chanx_right_in[7]
+ sb_5__3_/chanx_right_in[8] sb_5__3_/chanx_right_in[9] cbx_6__3_/chanx_left_in[0]
+ cbx_6__3_/chanx_left_in[10] cbx_6__3_/chanx_left_in[11] cbx_6__3_/chanx_left_in[12]
+ cbx_6__3_/chanx_left_in[13] cbx_6__3_/chanx_left_in[14] cbx_6__3_/chanx_left_in[15]
+ cbx_6__3_/chanx_left_in[16] cbx_6__3_/chanx_left_in[17] cbx_6__3_/chanx_left_in[18]
+ cbx_6__3_/chanx_left_in[19] cbx_6__3_/chanx_left_in[1] cbx_6__3_/chanx_left_in[2]
+ cbx_6__3_/chanx_left_in[3] cbx_6__3_/chanx_left_in[4] cbx_6__3_/chanx_left_in[5]
+ cbx_6__3_/chanx_left_in[6] cbx_6__3_/chanx_left_in[7] cbx_6__3_/chanx_left_in[8]
+ cbx_6__3_/chanx_left_in[9] cby_5__3_/chany_top_out[0] cby_5__3_/chany_top_out[10]
+ cby_5__3_/chany_top_out[11] cby_5__3_/chany_top_out[12] cby_5__3_/chany_top_out[13]
+ cby_5__3_/chany_top_out[14] cby_5__3_/chany_top_out[15] cby_5__3_/chany_top_out[16]
+ cby_5__3_/chany_top_out[17] cby_5__3_/chany_top_out[18] cby_5__3_/chany_top_out[19]
+ cby_5__3_/chany_top_out[1] cby_5__3_/chany_top_out[2] cby_5__3_/chany_top_out[3]
+ cby_5__3_/chany_top_out[4] cby_5__3_/chany_top_out[5] cby_5__3_/chany_top_out[6]
+ cby_5__3_/chany_top_out[7] cby_5__3_/chany_top_out[8] cby_5__3_/chany_top_out[9]
+ cby_5__3_/chany_top_in[0] cby_5__3_/chany_top_in[10] cby_5__3_/chany_top_in[11]
+ cby_5__3_/chany_top_in[12] cby_5__3_/chany_top_in[13] cby_5__3_/chany_top_in[14]
+ cby_5__3_/chany_top_in[15] cby_5__3_/chany_top_in[16] cby_5__3_/chany_top_in[17]
+ cby_5__3_/chany_top_in[18] cby_5__3_/chany_top_in[19] cby_5__3_/chany_top_in[1]
+ cby_5__3_/chany_top_in[2] cby_5__3_/chany_top_in[3] cby_5__3_/chany_top_in[4] cby_5__3_/chany_top_in[5]
+ cby_5__3_/chany_top_in[6] cby_5__3_/chany_top_in[7] cby_5__3_/chany_top_in[8] cby_5__3_/chany_top_in[9]
+ sb_5__3_/chany_top_in[0] sb_5__3_/chany_top_in[10] sb_5__3_/chany_top_in[11] sb_5__3_/chany_top_in[12]
+ sb_5__3_/chany_top_in[13] sb_5__3_/chany_top_in[14] sb_5__3_/chany_top_in[15] sb_5__3_/chany_top_in[16]
+ sb_5__3_/chany_top_in[17] sb_5__3_/chany_top_in[18] sb_5__3_/chany_top_in[19] sb_5__3_/chany_top_in[1]
+ sb_5__3_/chany_top_in[2] sb_5__3_/chany_top_in[3] sb_5__3_/chany_top_in[4] sb_5__3_/chany_top_in[5]
+ sb_5__3_/chany_top_in[6] sb_5__3_/chany_top_in[7] sb_5__3_/chany_top_in[8] sb_5__3_/chany_top_in[9]
+ sb_5__3_/chany_top_out[0] sb_5__3_/chany_top_out[10] sb_5__3_/chany_top_out[11]
+ sb_5__3_/chany_top_out[12] sb_5__3_/chany_top_out[13] sb_5__3_/chany_top_out[14]
+ sb_5__3_/chany_top_out[15] sb_5__3_/chany_top_out[16] sb_5__3_/chany_top_out[17]
+ sb_5__3_/chany_top_out[18] sb_5__3_/chany_top_out[19] sb_5__3_/chany_top_out[1]
+ sb_5__3_/chany_top_out[2] sb_5__3_/chany_top_out[3] sb_5__3_/chany_top_out[4] sb_5__3_/chany_top_out[5]
+ sb_5__3_/chany_top_out[6] sb_5__3_/chany_top_out[7] sb_5__3_/chany_top_out[8] sb_5__3_/chany_top_out[9]
+ sb_5__3_/clk_1_E_out sb_5__3_/clk_1_N_in sb_5__3_/clk_1_W_out sb_5__3_/clk_2_E_out
+ sb_5__3_/clk_2_N_in sb_5__3_/clk_2_N_out sb_5__3_/clk_2_S_out sb_5__3_/clk_2_W_out
+ sb_5__3_/clk_3_E_out sb_5__3_/clk_3_N_in sb_5__3_/clk_3_N_out sb_5__3_/clk_3_S_out
+ sb_5__3_/clk_3_W_out sb_5__3_/left_bottom_grid_pin_34_ sb_5__3_/left_bottom_grid_pin_35_
+ sb_5__3_/left_bottom_grid_pin_36_ sb_5__3_/left_bottom_grid_pin_37_ sb_5__3_/left_bottom_grid_pin_38_
+ sb_5__3_/left_bottom_grid_pin_39_ sb_5__3_/left_bottom_grid_pin_40_ sb_5__3_/left_bottom_grid_pin_41_
+ sb_5__3_/prog_clk_0_N_in sb_5__3_/prog_clk_1_E_out sb_5__3_/prog_clk_1_N_in sb_5__3_/prog_clk_1_W_out
+ sb_5__3_/prog_clk_2_E_out sb_5__3_/prog_clk_2_N_in sb_5__3_/prog_clk_2_N_out sb_5__3_/prog_clk_2_S_out
+ sb_5__3_/prog_clk_2_W_out sb_5__3_/prog_clk_3_E_out sb_5__3_/prog_clk_3_N_in sb_5__3_/prog_clk_3_N_out
+ sb_5__3_/prog_clk_3_S_out sb_5__3_/prog_clk_3_W_out sb_5__3_/right_bottom_grid_pin_34_
+ sb_5__3_/right_bottom_grid_pin_35_ sb_5__3_/right_bottom_grid_pin_36_ sb_5__3_/right_bottom_grid_pin_37_
+ sb_5__3_/right_bottom_grid_pin_38_ sb_5__3_/right_bottom_grid_pin_39_ sb_5__3_/right_bottom_grid_pin_40_
+ sb_5__3_/right_bottom_grid_pin_41_ sb_5__3_/top_left_grid_pin_42_ sb_5__3_/top_left_grid_pin_43_
+ sb_5__3_/top_left_grid_pin_44_ sb_5__3_/top_left_grid_pin_45_ sb_5__3_/top_left_grid_pin_46_
+ sb_5__3_/top_left_grid_pin_47_ sb_5__3_/top_left_grid_pin_48_ sb_5__3_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_7__1_ cbx_7__1_/SC_OUT_BOT cbx_7__0_/SC_IN_TOP grid_clb_7__1_/SC_OUT_TOP
+ cby_6__1_/Test_en_E_out cby_7__1_/Test_en_W_in cby_6__1_/Test_en_E_out grid_clb_7__1_/Test_en_W_out
+ VGND VPWR grid_clb_7__1_/bottom_width_0_height_0__pin_50_ grid_clb_7__1_/bottom_width_0_height_0__pin_51_
+ cby_6__1_/ccff_tail cby_7__1_/ccff_head cbx_7__1_/clk_1_S_out cbx_7__1_/clk_1_S_out
+ cby_7__1_/prog_clk_0_W_in cbx_7__1_/prog_clk_1_S_out grid_clb_7__1_/prog_clk_0_N_out
+ cbx_7__1_/prog_clk_1_S_out cbx_7__0_/prog_clk_0_N_in grid_clb_7__1_/prog_clk_0_W_out
+ cby_7__1_/left_grid_pin_16_ cby_7__1_/left_grid_pin_17_ cby_7__1_/left_grid_pin_18_
+ cby_7__1_/left_grid_pin_19_ cby_7__1_/left_grid_pin_20_ cby_7__1_/left_grid_pin_21_
+ cby_7__1_/left_grid_pin_22_ cby_7__1_/left_grid_pin_23_ cby_7__1_/left_grid_pin_24_
+ cby_7__1_/left_grid_pin_25_ cby_7__1_/left_grid_pin_26_ cby_7__1_/left_grid_pin_27_
+ cby_7__1_/left_grid_pin_28_ cby_7__1_/left_grid_pin_29_ cby_7__1_/left_grid_pin_30_
+ cby_7__1_/left_grid_pin_31_ sb_7__0_/top_left_grid_pin_42_ sb_7__1_/bottom_left_grid_pin_42_
+ sb_7__0_/top_left_grid_pin_43_ sb_7__1_/bottom_left_grid_pin_43_ sb_7__0_/top_left_grid_pin_44_
+ sb_7__1_/bottom_left_grid_pin_44_ sb_7__0_/top_left_grid_pin_45_ sb_7__1_/bottom_left_grid_pin_45_
+ sb_7__0_/top_left_grid_pin_46_ sb_7__1_/bottom_left_grid_pin_46_ sb_7__0_/top_left_grid_pin_47_
+ sb_7__1_/bottom_left_grid_pin_47_ sb_7__0_/top_left_grid_pin_48_ sb_7__1_/bottom_left_grid_pin_48_
+ sb_7__0_/top_left_grid_pin_49_ sb_7__1_/bottom_left_grid_pin_49_ cbx_7__1_/bottom_grid_pin_0_
+ cbx_7__1_/bottom_grid_pin_10_ cbx_7__1_/bottom_grid_pin_11_ cbx_7__1_/bottom_grid_pin_12_
+ cbx_7__1_/bottom_grid_pin_13_ cbx_7__1_/bottom_grid_pin_14_ cbx_7__1_/bottom_grid_pin_15_
+ cbx_7__1_/bottom_grid_pin_1_ cbx_7__1_/bottom_grid_pin_2_ cbx_7__1_/REGOUT_FEEDTHROUGH
+ grid_clb_7__1_/top_width_0_height_0__pin_33_ sb_7__1_/left_bottom_grid_pin_34_ sb_6__1_/right_bottom_grid_pin_34_
+ sb_7__1_/left_bottom_grid_pin_35_ sb_6__1_/right_bottom_grid_pin_35_ sb_7__1_/left_bottom_grid_pin_36_
+ sb_6__1_/right_bottom_grid_pin_36_ sb_7__1_/left_bottom_grid_pin_37_ sb_6__1_/right_bottom_grid_pin_37_
+ sb_7__1_/left_bottom_grid_pin_38_ sb_6__1_/right_bottom_grid_pin_38_ sb_7__1_/left_bottom_grid_pin_39_
+ sb_6__1_/right_bottom_grid_pin_39_ cbx_7__1_/bottom_grid_pin_3_ sb_7__1_/left_bottom_grid_pin_40_
+ sb_6__1_/right_bottom_grid_pin_40_ sb_7__1_/left_bottom_grid_pin_41_ sb_6__1_/right_bottom_grid_pin_41_
+ cbx_7__1_/bottom_grid_pin_4_ cbx_7__1_/bottom_grid_pin_5_ cbx_7__1_/bottom_grid_pin_6_
+ cbx_7__1_/bottom_grid_pin_7_ cbx_7__1_/bottom_grid_pin_8_ cbx_7__1_/bottom_grid_pin_9_
+ grid_clb
Xsb_2__0_ sb_2__0_/SC_IN_TOP sb_2__0_/SC_OUT_TOP sb_2__0_/Test_en_N_out sb_2__0_/Test_en_S_in
+ VGND VPWR sb_2__0_/ccff_head sb_2__0_/ccff_tail sb_2__0_/chanx_left_in[0] sb_2__0_/chanx_left_in[10]
+ sb_2__0_/chanx_left_in[11] sb_2__0_/chanx_left_in[12] sb_2__0_/chanx_left_in[13]
+ sb_2__0_/chanx_left_in[14] sb_2__0_/chanx_left_in[15] sb_2__0_/chanx_left_in[16]
+ sb_2__0_/chanx_left_in[17] sb_2__0_/chanx_left_in[18] sb_2__0_/chanx_left_in[19]
+ sb_2__0_/chanx_left_in[1] sb_2__0_/chanx_left_in[2] sb_2__0_/chanx_left_in[3] sb_2__0_/chanx_left_in[4]
+ sb_2__0_/chanx_left_in[5] sb_2__0_/chanx_left_in[6] sb_2__0_/chanx_left_in[7] sb_2__0_/chanx_left_in[8]
+ sb_2__0_/chanx_left_in[9] sb_2__0_/chanx_left_out[0] sb_2__0_/chanx_left_out[10]
+ sb_2__0_/chanx_left_out[11] sb_2__0_/chanx_left_out[12] sb_2__0_/chanx_left_out[13]
+ sb_2__0_/chanx_left_out[14] sb_2__0_/chanx_left_out[15] sb_2__0_/chanx_left_out[16]
+ sb_2__0_/chanx_left_out[17] sb_2__0_/chanx_left_out[18] sb_2__0_/chanx_left_out[19]
+ sb_2__0_/chanx_left_out[1] sb_2__0_/chanx_left_out[2] sb_2__0_/chanx_left_out[3]
+ sb_2__0_/chanx_left_out[4] sb_2__0_/chanx_left_out[5] sb_2__0_/chanx_left_out[6]
+ sb_2__0_/chanx_left_out[7] sb_2__0_/chanx_left_out[8] sb_2__0_/chanx_left_out[9]
+ sb_2__0_/chanx_right_in[0] sb_2__0_/chanx_right_in[10] sb_2__0_/chanx_right_in[11]
+ sb_2__0_/chanx_right_in[12] sb_2__0_/chanx_right_in[13] sb_2__0_/chanx_right_in[14]
+ sb_2__0_/chanx_right_in[15] sb_2__0_/chanx_right_in[16] sb_2__0_/chanx_right_in[17]
+ sb_2__0_/chanx_right_in[18] sb_2__0_/chanx_right_in[19] sb_2__0_/chanx_right_in[1]
+ sb_2__0_/chanx_right_in[2] sb_2__0_/chanx_right_in[3] sb_2__0_/chanx_right_in[4]
+ sb_2__0_/chanx_right_in[5] sb_2__0_/chanx_right_in[6] sb_2__0_/chanx_right_in[7]
+ sb_2__0_/chanx_right_in[8] sb_2__0_/chanx_right_in[9] cbx_3__0_/chanx_left_in[0]
+ cbx_3__0_/chanx_left_in[10] cbx_3__0_/chanx_left_in[11] cbx_3__0_/chanx_left_in[12]
+ cbx_3__0_/chanx_left_in[13] cbx_3__0_/chanx_left_in[14] cbx_3__0_/chanx_left_in[15]
+ cbx_3__0_/chanx_left_in[16] cbx_3__0_/chanx_left_in[17] cbx_3__0_/chanx_left_in[18]
+ cbx_3__0_/chanx_left_in[19] cbx_3__0_/chanx_left_in[1] cbx_3__0_/chanx_left_in[2]
+ cbx_3__0_/chanx_left_in[3] cbx_3__0_/chanx_left_in[4] cbx_3__0_/chanx_left_in[5]
+ cbx_3__0_/chanx_left_in[6] cbx_3__0_/chanx_left_in[7] cbx_3__0_/chanx_left_in[8]
+ cbx_3__0_/chanx_left_in[9] sb_2__0_/chany_top_in[0] sb_2__0_/chany_top_in[10] sb_2__0_/chany_top_in[11]
+ sb_2__0_/chany_top_in[12] sb_2__0_/chany_top_in[13] sb_2__0_/chany_top_in[14] sb_2__0_/chany_top_in[15]
+ sb_2__0_/chany_top_in[16] sb_2__0_/chany_top_in[17] sb_2__0_/chany_top_in[18] sb_2__0_/chany_top_in[19]
+ sb_2__0_/chany_top_in[1] sb_2__0_/chany_top_in[2] sb_2__0_/chany_top_in[3] sb_2__0_/chany_top_in[4]
+ sb_2__0_/chany_top_in[5] sb_2__0_/chany_top_in[6] sb_2__0_/chany_top_in[7] sb_2__0_/chany_top_in[8]
+ sb_2__0_/chany_top_in[9] sb_2__0_/chany_top_out[0] sb_2__0_/chany_top_out[10] sb_2__0_/chany_top_out[11]
+ sb_2__0_/chany_top_out[12] sb_2__0_/chany_top_out[13] sb_2__0_/chany_top_out[14]
+ sb_2__0_/chany_top_out[15] sb_2__0_/chany_top_out[16] sb_2__0_/chany_top_out[17]
+ sb_2__0_/chany_top_out[18] sb_2__0_/chany_top_out[19] sb_2__0_/chany_top_out[1]
+ sb_2__0_/chany_top_out[2] sb_2__0_/chany_top_out[3] sb_2__0_/chany_top_out[4] sb_2__0_/chany_top_out[5]
+ sb_2__0_/chany_top_out[6] sb_2__0_/chany_top_out[7] sb_2__0_/chany_top_out[8] sb_2__0_/chany_top_out[9]
+ sb_2__0_/clk_3_N_out sb_2__0_/clk_3_S_in sb_2__0_/left_bottom_grid_pin_11_ sb_2__0_/left_bottom_grid_pin_13_
+ sb_2__0_/left_bottom_grid_pin_15_ sb_2__0_/left_bottom_grid_pin_17_ sb_2__0_/left_bottom_grid_pin_1_
+ sb_2__0_/left_bottom_grid_pin_3_ sb_2__0_/left_bottom_grid_pin_5_ sb_2__0_/left_bottom_grid_pin_7_
+ sb_2__0_/left_bottom_grid_pin_9_ sb_2__0_/prog_clk_0_N_in sb_2__0_/prog_clk_3_N_out
+ sb_2__0_/prog_clk_3_S_in sb_2__0_/right_bottom_grid_pin_11_ sb_2__0_/right_bottom_grid_pin_13_
+ sb_2__0_/right_bottom_grid_pin_15_ sb_2__0_/right_bottom_grid_pin_17_ sb_2__0_/right_bottom_grid_pin_1_
+ sb_2__0_/right_bottom_grid_pin_3_ sb_2__0_/right_bottom_grid_pin_5_ sb_2__0_/right_bottom_grid_pin_7_
+ sb_2__0_/right_bottom_grid_pin_9_ sb_2__0_/top_left_grid_pin_42_ sb_2__0_/top_left_grid_pin_43_
+ sb_2__0_/top_left_grid_pin_44_ sb_2__0_/top_left_grid_pin_45_ sb_2__0_/top_left_grid_pin_46_
+ sb_2__0_/top_left_grid_pin_47_ sb_2__0_/top_left_grid_pin_48_ sb_2__0_/top_left_grid_pin_49_
+ sb_1__0_
Xcby_4__7_ sb_4__6_/Test_en_N_out cby_4__7_/Test_en_E_out sb_4__7_/Test_en_S_in sb_4__6_/Test_en_N_out
+ sb_4__6_/Test_en_N_out cby_4__7_/Test_en_W_out VGND VPWR cby_4__7_/ccff_head cby_4__7_/ccff_tail
+ sb_4__6_/chany_top_out[0] sb_4__6_/chany_top_out[10] sb_4__6_/chany_top_out[11]
+ sb_4__6_/chany_top_out[12] sb_4__6_/chany_top_out[13] sb_4__6_/chany_top_out[14]
+ sb_4__6_/chany_top_out[15] sb_4__6_/chany_top_out[16] sb_4__6_/chany_top_out[17]
+ sb_4__6_/chany_top_out[18] sb_4__6_/chany_top_out[19] sb_4__6_/chany_top_out[1]
+ sb_4__6_/chany_top_out[2] sb_4__6_/chany_top_out[3] sb_4__6_/chany_top_out[4] sb_4__6_/chany_top_out[5]
+ sb_4__6_/chany_top_out[6] sb_4__6_/chany_top_out[7] sb_4__6_/chany_top_out[8] sb_4__6_/chany_top_out[9]
+ sb_4__6_/chany_top_in[0] sb_4__6_/chany_top_in[10] sb_4__6_/chany_top_in[11] sb_4__6_/chany_top_in[12]
+ sb_4__6_/chany_top_in[13] sb_4__6_/chany_top_in[14] sb_4__6_/chany_top_in[15] sb_4__6_/chany_top_in[16]
+ sb_4__6_/chany_top_in[17] sb_4__6_/chany_top_in[18] sb_4__6_/chany_top_in[19] sb_4__6_/chany_top_in[1]
+ sb_4__6_/chany_top_in[2] sb_4__6_/chany_top_in[3] sb_4__6_/chany_top_in[4] sb_4__6_/chany_top_in[5]
+ sb_4__6_/chany_top_in[6] sb_4__6_/chany_top_in[7] sb_4__6_/chany_top_in[8] sb_4__6_/chany_top_in[9]
+ cby_4__7_/chany_top_in[0] cby_4__7_/chany_top_in[10] cby_4__7_/chany_top_in[11]
+ cby_4__7_/chany_top_in[12] cby_4__7_/chany_top_in[13] cby_4__7_/chany_top_in[14]
+ cby_4__7_/chany_top_in[15] cby_4__7_/chany_top_in[16] cby_4__7_/chany_top_in[17]
+ cby_4__7_/chany_top_in[18] cby_4__7_/chany_top_in[19] cby_4__7_/chany_top_in[1]
+ cby_4__7_/chany_top_in[2] cby_4__7_/chany_top_in[3] cby_4__7_/chany_top_in[4] cby_4__7_/chany_top_in[5]
+ cby_4__7_/chany_top_in[6] cby_4__7_/chany_top_in[7] cby_4__7_/chany_top_in[8] cby_4__7_/chany_top_in[9]
+ cby_4__7_/chany_top_out[0] cby_4__7_/chany_top_out[10] cby_4__7_/chany_top_out[11]
+ cby_4__7_/chany_top_out[12] cby_4__7_/chany_top_out[13] cby_4__7_/chany_top_out[14]
+ cby_4__7_/chany_top_out[15] cby_4__7_/chany_top_out[16] cby_4__7_/chany_top_out[17]
+ cby_4__7_/chany_top_out[18] cby_4__7_/chany_top_out[19] cby_4__7_/chany_top_out[1]
+ cby_4__7_/chany_top_out[2] cby_4__7_/chany_top_out[3] cby_4__7_/chany_top_out[4]
+ cby_4__7_/chany_top_out[5] cby_4__7_/chany_top_out[6] cby_4__7_/chany_top_out[7]
+ cby_4__7_/chany_top_out[8] cby_4__7_/chany_top_out[9] cby_4__7_/clk_2_N_out cby_4__7_/clk_2_S_in
+ cby_4__7_/clk_2_S_out cby_4__7_/clk_3_N_out cby_4__7_/clk_3_S_in cby_4__7_/clk_3_S_out
+ cby_4__7_/left_grid_pin_16_ cby_4__7_/left_grid_pin_17_ cby_4__7_/left_grid_pin_18_
+ cby_4__7_/left_grid_pin_19_ cby_4__7_/left_grid_pin_20_ cby_4__7_/left_grid_pin_21_
+ cby_4__7_/left_grid_pin_22_ cby_4__7_/left_grid_pin_23_ cby_4__7_/left_grid_pin_24_
+ cby_4__7_/left_grid_pin_25_ cby_4__7_/left_grid_pin_26_ cby_4__7_/left_grid_pin_27_
+ cby_4__7_/left_grid_pin_28_ cby_4__7_/left_grid_pin_29_ cby_4__7_/left_grid_pin_30_
+ cby_4__7_/left_grid_pin_31_ cby_4__7_/prog_clk_0_N_out sb_4__6_/prog_clk_0_N_in
+ cby_4__7_/prog_clk_0_W_in cby_4__7_/prog_clk_2_N_out cby_4__7_/prog_clk_2_S_in cby_4__7_/prog_clk_2_S_out
+ cby_4__7_/prog_clk_3_N_out cby_4__7_/prog_clk_3_S_in cby_4__7_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_4__8_ IO_ISOL_N cbx_4__8_/SC_IN_BOT cbx_4__8_/SC_IN_TOP cbx_4__8_/SC_OUT_BOT
+ sb_4__8_/SC_IN_BOT VGND VPWR cbx_4__8_/bottom_grid_pin_0_ cbx_4__8_/bottom_grid_pin_10_
+ cbx_4__8_/bottom_grid_pin_11_ cbx_4__8_/bottom_grid_pin_12_ cbx_4__8_/bottom_grid_pin_13_
+ cbx_4__8_/bottom_grid_pin_14_ cbx_4__8_/bottom_grid_pin_15_ cbx_4__8_/bottom_grid_pin_1_
+ cbx_4__8_/bottom_grid_pin_2_ cbx_4__8_/bottom_grid_pin_3_ cbx_4__8_/bottom_grid_pin_4_
+ cbx_4__8_/bottom_grid_pin_5_ cbx_4__8_/bottom_grid_pin_6_ cbx_4__8_/bottom_grid_pin_7_
+ cbx_4__8_/bottom_grid_pin_8_ cbx_4__8_/bottom_grid_pin_9_ cbx_4__8_/top_grid_pin_0_
+ sb_4__8_/left_top_grid_pin_1_ sb_3__8_/right_top_grid_pin_1_ sb_4__8_/ccff_tail
+ sb_3__8_/ccff_head cbx_4__8_/chanx_left_in[0] cbx_4__8_/chanx_left_in[10] cbx_4__8_/chanx_left_in[11]
+ cbx_4__8_/chanx_left_in[12] cbx_4__8_/chanx_left_in[13] cbx_4__8_/chanx_left_in[14]
+ cbx_4__8_/chanx_left_in[15] cbx_4__8_/chanx_left_in[16] cbx_4__8_/chanx_left_in[17]
+ cbx_4__8_/chanx_left_in[18] cbx_4__8_/chanx_left_in[19] cbx_4__8_/chanx_left_in[1]
+ cbx_4__8_/chanx_left_in[2] cbx_4__8_/chanx_left_in[3] cbx_4__8_/chanx_left_in[4]
+ cbx_4__8_/chanx_left_in[5] cbx_4__8_/chanx_left_in[6] cbx_4__8_/chanx_left_in[7]
+ cbx_4__8_/chanx_left_in[8] cbx_4__8_/chanx_left_in[9] sb_3__8_/chanx_right_in[0]
+ sb_3__8_/chanx_right_in[10] sb_3__8_/chanx_right_in[11] sb_3__8_/chanx_right_in[12]
+ sb_3__8_/chanx_right_in[13] sb_3__8_/chanx_right_in[14] sb_3__8_/chanx_right_in[15]
+ sb_3__8_/chanx_right_in[16] sb_3__8_/chanx_right_in[17] sb_3__8_/chanx_right_in[18]
+ sb_3__8_/chanx_right_in[19] sb_3__8_/chanx_right_in[1] sb_3__8_/chanx_right_in[2]
+ sb_3__8_/chanx_right_in[3] sb_3__8_/chanx_right_in[4] sb_3__8_/chanx_right_in[5]
+ sb_3__8_/chanx_right_in[6] sb_3__8_/chanx_right_in[7] sb_3__8_/chanx_right_in[8]
+ sb_3__8_/chanx_right_in[9] sb_4__8_/chanx_left_out[0] sb_4__8_/chanx_left_out[10]
+ sb_4__8_/chanx_left_out[11] sb_4__8_/chanx_left_out[12] sb_4__8_/chanx_left_out[13]
+ sb_4__8_/chanx_left_out[14] sb_4__8_/chanx_left_out[15] sb_4__8_/chanx_left_out[16]
+ sb_4__8_/chanx_left_out[17] sb_4__8_/chanx_left_out[18] sb_4__8_/chanx_left_out[19]
+ sb_4__8_/chanx_left_out[1] sb_4__8_/chanx_left_out[2] sb_4__8_/chanx_left_out[3]
+ sb_4__8_/chanx_left_out[4] sb_4__8_/chanx_left_out[5] sb_4__8_/chanx_left_out[6]
+ sb_4__8_/chanx_left_out[7] sb_4__8_/chanx_left_out[8] sb_4__8_/chanx_left_out[9]
+ sb_4__8_/chanx_left_in[0] sb_4__8_/chanx_left_in[10] sb_4__8_/chanx_left_in[11]
+ sb_4__8_/chanx_left_in[12] sb_4__8_/chanx_left_in[13] sb_4__8_/chanx_left_in[14]
+ sb_4__8_/chanx_left_in[15] sb_4__8_/chanx_left_in[16] sb_4__8_/chanx_left_in[17]
+ sb_4__8_/chanx_left_in[18] sb_4__8_/chanx_left_in[19] sb_4__8_/chanx_left_in[1]
+ sb_4__8_/chanx_left_in[2] sb_4__8_/chanx_left_in[3] sb_4__8_/chanx_left_in[4] sb_4__8_/chanx_left_in[5]
+ sb_4__8_/chanx_left_in[6] sb_4__8_/chanx_left_in[7] sb_4__8_/chanx_left_in[8] sb_4__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
+ cbx_4__8_/prog_clk_0_S_in cbx_4__8_/prog_clk_0_W_out cbx_4__8_/top_grid_pin_0_ cbx_1__2_
Xsb_8__5_ VGND VPWR sb_8__5_/bottom_left_grid_pin_42_ sb_8__5_/bottom_left_grid_pin_43_
+ sb_8__5_/bottom_left_grid_pin_44_ sb_8__5_/bottom_left_grid_pin_45_ sb_8__5_/bottom_left_grid_pin_46_
+ sb_8__5_/bottom_left_grid_pin_47_ sb_8__5_/bottom_left_grid_pin_48_ sb_8__5_/bottom_left_grid_pin_49_
+ sb_8__5_/bottom_right_grid_pin_1_ sb_8__5_/ccff_head sb_8__5_/ccff_tail sb_8__5_/chanx_left_in[0]
+ sb_8__5_/chanx_left_in[10] sb_8__5_/chanx_left_in[11] sb_8__5_/chanx_left_in[12]
+ sb_8__5_/chanx_left_in[13] sb_8__5_/chanx_left_in[14] sb_8__5_/chanx_left_in[15]
+ sb_8__5_/chanx_left_in[16] sb_8__5_/chanx_left_in[17] sb_8__5_/chanx_left_in[18]
+ sb_8__5_/chanx_left_in[19] sb_8__5_/chanx_left_in[1] sb_8__5_/chanx_left_in[2] sb_8__5_/chanx_left_in[3]
+ sb_8__5_/chanx_left_in[4] sb_8__5_/chanx_left_in[5] sb_8__5_/chanx_left_in[6] sb_8__5_/chanx_left_in[7]
+ sb_8__5_/chanx_left_in[8] sb_8__5_/chanx_left_in[9] sb_8__5_/chanx_left_out[0] sb_8__5_/chanx_left_out[10]
+ sb_8__5_/chanx_left_out[11] sb_8__5_/chanx_left_out[12] sb_8__5_/chanx_left_out[13]
+ sb_8__5_/chanx_left_out[14] sb_8__5_/chanx_left_out[15] sb_8__5_/chanx_left_out[16]
+ sb_8__5_/chanx_left_out[17] sb_8__5_/chanx_left_out[18] sb_8__5_/chanx_left_out[19]
+ sb_8__5_/chanx_left_out[1] sb_8__5_/chanx_left_out[2] sb_8__5_/chanx_left_out[3]
+ sb_8__5_/chanx_left_out[4] sb_8__5_/chanx_left_out[5] sb_8__5_/chanx_left_out[6]
+ sb_8__5_/chanx_left_out[7] sb_8__5_/chanx_left_out[8] sb_8__5_/chanx_left_out[9]
+ cby_8__5_/chany_top_out[0] cby_8__5_/chany_top_out[10] cby_8__5_/chany_top_out[11]
+ cby_8__5_/chany_top_out[12] cby_8__5_/chany_top_out[13] cby_8__5_/chany_top_out[14]
+ cby_8__5_/chany_top_out[15] cby_8__5_/chany_top_out[16] cby_8__5_/chany_top_out[17]
+ cby_8__5_/chany_top_out[18] cby_8__5_/chany_top_out[19] cby_8__5_/chany_top_out[1]
+ cby_8__5_/chany_top_out[2] cby_8__5_/chany_top_out[3] cby_8__5_/chany_top_out[4]
+ cby_8__5_/chany_top_out[5] cby_8__5_/chany_top_out[6] cby_8__5_/chany_top_out[7]
+ cby_8__5_/chany_top_out[8] cby_8__5_/chany_top_out[9] cby_8__5_/chany_top_in[0]
+ cby_8__5_/chany_top_in[10] cby_8__5_/chany_top_in[11] cby_8__5_/chany_top_in[12]
+ cby_8__5_/chany_top_in[13] cby_8__5_/chany_top_in[14] cby_8__5_/chany_top_in[15]
+ cby_8__5_/chany_top_in[16] cby_8__5_/chany_top_in[17] cby_8__5_/chany_top_in[18]
+ cby_8__5_/chany_top_in[19] cby_8__5_/chany_top_in[1] cby_8__5_/chany_top_in[2] cby_8__5_/chany_top_in[3]
+ cby_8__5_/chany_top_in[4] cby_8__5_/chany_top_in[5] cby_8__5_/chany_top_in[6] cby_8__5_/chany_top_in[7]
+ cby_8__5_/chany_top_in[8] cby_8__5_/chany_top_in[9] sb_8__5_/chany_top_in[0] sb_8__5_/chany_top_in[10]
+ sb_8__5_/chany_top_in[11] sb_8__5_/chany_top_in[12] sb_8__5_/chany_top_in[13] sb_8__5_/chany_top_in[14]
+ sb_8__5_/chany_top_in[15] sb_8__5_/chany_top_in[16] sb_8__5_/chany_top_in[17] sb_8__5_/chany_top_in[18]
+ sb_8__5_/chany_top_in[19] sb_8__5_/chany_top_in[1] sb_8__5_/chany_top_in[2] sb_8__5_/chany_top_in[3]
+ sb_8__5_/chany_top_in[4] sb_8__5_/chany_top_in[5] sb_8__5_/chany_top_in[6] sb_8__5_/chany_top_in[7]
+ sb_8__5_/chany_top_in[8] sb_8__5_/chany_top_in[9] sb_8__5_/chany_top_out[0] sb_8__5_/chany_top_out[10]
+ sb_8__5_/chany_top_out[11] sb_8__5_/chany_top_out[12] sb_8__5_/chany_top_out[13]
+ sb_8__5_/chany_top_out[14] sb_8__5_/chany_top_out[15] sb_8__5_/chany_top_out[16]
+ sb_8__5_/chany_top_out[17] sb_8__5_/chany_top_out[18] sb_8__5_/chany_top_out[19]
+ sb_8__5_/chany_top_out[1] sb_8__5_/chany_top_out[2] sb_8__5_/chany_top_out[3] sb_8__5_/chany_top_out[4]
+ sb_8__5_/chany_top_out[5] sb_8__5_/chany_top_out[6] sb_8__5_/chany_top_out[7] sb_8__5_/chany_top_out[8]
+ sb_8__5_/chany_top_out[9] sb_8__5_/left_bottom_grid_pin_34_ sb_8__5_/left_bottom_grid_pin_35_
+ sb_8__5_/left_bottom_grid_pin_36_ sb_8__5_/left_bottom_grid_pin_37_ sb_8__5_/left_bottom_grid_pin_38_
+ sb_8__5_/left_bottom_grid_pin_39_ sb_8__5_/left_bottom_grid_pin_40_ sb_8__5_/left_bottom_grid_pin_41_
+ sb_8__5_/prog_clk_0_N_in sb_8__5_/top_left_grid_pin_42_ sb_8__5_/top_left_grid_pin_43_
+ sb_8__5_/top_left_grid_pin_44_ sb_8__5_/top_left_grid_pin_45_ sb_8__5_/top_left_grid_pin_46_
+ sb_8__5_/top_left_grid_pin_47_ sb_8__5_/top_left_grid_pin_48_ sb_8__5_/top_left_grid_pin_49_
+ sb_8__5_/top_right_grid_pin_1_ sb_2__1_
Xcby_1__4_ cby_1__4_/Test_en_W_in cby_1__4_/Test_en_E_out cby_1__4_/Test_en_N_out
+ cby_1__4_/Test_en_W_in cby_1__4_/Test_en_W_in cby_1__4_/Test_en_W_out VGND VPWR
+ cby_1__4_/ccff_head cby_1__4_/ccff_tail sb_1__3_/chany_top_out[0] sb_1__3_/chany_top_out[10]
+ sb_1__3_/chany_top_out[11] sb_1__3_/chany_top_out[12] sb_1__3_/chany_top_out[13]
+ sb_1__3_/chany_top_out[14] sb_1__3_/chany_top_out[15] sb_1__3_/chany_top_out[16]
+ sb_1__3_/chany_top_out[17] sb_1__3_/chany_top_out[18] sb_1__3_/chany_top_out[19]
+ sb_1__3_/chany_top_out[1] sb_1__3_/chany_top_out[2] sb_1__3_/chany_top_out[3] sb_1__3_/chany_top_out[4]
+ sb_1__3_/chany_top_out[5] sb_1__3_/chany_top_out[6] sb_1__3_/chany_top_out[7] sb_1__3_/chany_top_out[8]
+ sb_1__3_/chany_top_out[9] sb_1__3_/chany_top_in[0] sb_1__3_/chany_top_in[10] sb_1__3_/chany_top_in[11]
+ sb_1__3_/chany_top_in[12] sb_1__3_/chany_top_in[13] sb_1__3_/chany_top_in[14] sb_1__3_/chany_top_in[15]
+ sb_1__3_/chany_top_in[16] sb_1__3_/chany_top_in[17] sb_1__3_/chany_top_in[18] sb_1__3_/chany_top_in[19]
+ sb_1__3_/chany_top_in[1] sb_1__3_/chany_top_in[2] sb_1__3_/chany_top_in[3] sb_1__3_/chany_top_in[4]
+ sb_1__3_/chany_top_in[5] sb_1__3_/chany_top_in[6] sb_1__3_/chany_top_in[7] sb_1__3_/chany_top_in[8]
+ sb_1__3_/chany_top_in[9] cby_1__4_/chany_top_in[0] cby_1__4_/chany_top_in[10] cby_1__4_/chany_top_in[11]
+ cby_1__4_/chany_top_in[12] cby_1__4_/chany_top_in[13] cby_1__4_/chany_top_in[14]
+ cby_1__4_/chany_top_in[15] cby_1__4_/chany_top_in[16] cby_1__4_/chany_top_in[17]
+ cby_1__4_/chany_top_in[18] cby_1__4_/chany_top_in[19] cby_1__4_/chany_top_in[1]
+ cby_1__4_/chany_top_in[2] cby_1__4_/chany_top_in[3] cby_1__4_/chany_top_in[4] cby_1__4_/chany_top_in[5]
+ cby_1__4_/chany_top_in[6] cby_1__4_/chany_top_in[7] cby_1__4_/chany_top_in[8] cby_1__4_/chany_top_in[9]
+ cby_1__4_/chany_top_out[0] cby_1__4_/chany_top_out[10] cby_1__4_/chany_top_out[11]
+ cby_1__4_/chany_top_out[12] cby_1__4_/chany_top_out[13] cby_1__4_/chany_top_out[14]
+ cby_1__4_/chany_top_out[15] cby_1__4_/chany_top_out[16] cby_1__4_/chany_top_out[17]
+ cby_1__4_/chany_top_out[18] cby_1__4_/chany_top_out[19] cby_1__4_/chany_top_out[1]
+ cby_1__4_/chany_top_out[2] cby_1__4_/chany_top_out[3] cby_1__4_/chany_top_out[4]
+ cby_1__4_/chany_top_out[5] cby_1__4_/chany_top_out[6] cby_1__4_/chany_top_out[7]
+ cby_1__4_/chany_top_out[8] cby_1__4_/chany_top_out[9] cby_1__4_/clk_2_N_out cby_1__4_/clk_2_S_in
+ cby_1__4_/clk_2_S_out cby_1__4_/clk_3_N_out cby_1__4_/clk_3_S_in cby_1__4_/clk_3_S_out
+ cby_1__4_/left_grid_pin_16_ cby_1__4_/left_grid_pin_17_ cby_1__4_/left_grid_pin_18_
+ cby_1__4_/left_grid_pin_19_ cby_1__4_/left_grid_pin_20_ cby_1__4_/left_grid_pin_21_
+ cby_1__4_/left_grid_pin_22_ cby_1__4_/left_grid_pin_23_ cby_1__4_/left_grid_pin_24_
+ cby_1__4_/left_grid_pin_25_ cby_1__4_/left_grid_pin_26_ cby_1__4_/left_grid_pin_27_
+ cby_1__4_/left_grid_pin_28_ cby_1__4_/left_grid_pin_29_ cby_1__4_/left_grid_pin_30_
+ cby_1__4_/left_grid_pin_31_ cby_1__4_/prog_clk_0_N_out sb_1__3_/prog_clk_0_N_in
+ cby_1__4_/prog_clk_0_W_in cby_1__4_/prog_clk_2_N_out cby_1__4_/prog_clk_2_S_in cby_1__4_/prog_clk_2_S_out
+ cby_1__4_/prog_clk_3_N_out cby_1__4_/prog_clk_3_S_in cby_1__4_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_8__0_ IO_ISOL_N sb_7__0_/SC_OUT_TOP cbx_8__0_/SC_IN_TOP cbx_8__0_/SC_OUT_BOT
+ cbx_8__0_/SC_OUT_TOP VGND VPWR cbx_8__0_/bottom_grid_pin_0_ cbx_8__0_/bottom_grid_pin_10_
+ cbx_8__0_/bottom_grid_pin_12_ cbx_8__0_/bottom_grid_pin_14_ cbx_8__0_/bottom_grid_pin_16_
+ cbx_8__0_/bottom_grid_pin_2_ cbx_8__0_/bottom_grid_pin_4_ cbx_8__0_/bottom_grid_pin_6_
+ cbx_8__0_/bottom_grid_pin_8_ sb_8__0_/ccff_tail sb_7__0_/ccff_head cbx_8__0_/chanx_left_in[0]
+ cbx_8__0_/chanx_left_in[10] cbx_8__0_/chanx_left_in[11] cbx_8__0_/chanx_left_in[12]
+ cbx_8__0_/chanx_left_in[13] cbx_8__0_/chanx_left_in[14] cbx_8__0_/chanx_left_in[15]
+ cbx_8__0_/chanx_left_in[16] cbx_8__0_/chanx_left_in[17] cbx_8__0_/chanx_left_in[18]
+ cbx_8__0_/chanx_left_in[19] cbx_8__0_/chanx_left_in[1] cbx_8__0_/chanx_left_in[2]
+ cbx_8__0_/chanx_left_in[3] cbx_8__0_/chanx_left_in[4] cbx_8__0_/chanx_left_in[5]
+ cbx_8__0_/chanx_left_in[6] cbx_8__0_/chanx_left_in[7] cbx_8__0_/chanx_left_in[8]
+ cbx_8__0_/chanx_left_in[9] sb_7__0_/chanx_right_in[0] sb_7__0_/chanx_right_in[10]
+ sb_7__0_/chanx_right_in[11] sb_7__0_/chanx_right_in[12] sb_7__0_/chanx_right_in[13]
+ sb_7__0_/chanx_right_in[14] sb_7__0_/chanx_right_in[15] sb_7__0_/chanx_right_in[16]
+ sb_7__0_/chanx_right_in[17] sb_7__0_/chanx_right_in[18] sb_7__0_/chanx_right_in[19]
+ sb_7__0_/chanx_right_in[1] sb_7__0_/chanx_right_in[2] sb_7__0_/chanx_right_in[3]
+ sb_7__0_/chanx_right_in[4] sb_7__0_/chanx_right_in[5] sb_7__0_/chanx_right_in[6]
+ sb_7__0_/chanx_right_in[7] sb_7__0_/chanx_right_in[8] sb_7__0_/chanx_right_in[9]
+ sb_8__0_/chanx_left_out[0] sb_8__0_/chanx_left_out[10] sb_8__0_/chanx_left_out[11]
+ sb_8__0_/chanx_left_out[12] sb_8__0_/chanx_left_out[13] sb_8__0_/chanx_left_out[14]
+ sb_8__0_/chanx_left_out[15] sb_8__0_/chanx_left_out[16] sb_8__0_/chanx_left_out[17]
+ sb_8__0_/chanx_left_out[18] sb_8__0_/chanx_left_out[19] sb_8__0_/chanx_left_out[1]
+ sb_8__0_/chanx_left_out[2] sb_8__0_/chanx_left_out[3] sb_8__0_/chanx_left_out[4]
+ sb_8__0_/chanx_left_out[5] sb_8__0_/chanx_left_out[6] sb_8__0_/chanx_left_out[7]
+ sb_8__0_/chanx_left_out[8] sb_8__0_/chanx_left_out[9] sb_8__0_/chanx_left_in[0]
+ sb_8__0_/chanx_left_in[10] sb_8__0_/chanx_left_in[11] sb_8__0_/chanx_left_in[12]
+ sb_8__0_/chanx_left_in[13] sb_8__0_/chanx_left_in[14] sb_8__0_/chanx_left_in[15]
+ sb_8__0_/chanx_left_in[16] sb_8__0_/chanx_left_in[17] sb_8__0_/chanx_left_in[18]
+ sb_8__0_/chanx_left_in[19] sb_8__0_/chanx_left_in[1] sb_8__0_/chanx_left_in[2] sb_8__0_/chanx_left_in[3]
+ sb_8__0_/chanx_left_in[4] sb_8__0_/chanx_left_in[5] sb_8__0_/chanx_left_in[6] sb_8__0_/chanx_left_in[7]
+ sb_8__0_/chanx_left_in[8] sb_8__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24] cbx_8__0_/prog_clk_0_N_in
+ cbx_8__0_/prog_clk_0_W_out cbx_8__0_/bottom_grid_pin_0_ cbx_8__0_/bottom_grid_pin_10_
+ sb_8__0_/left_bottom_grid_pin_11_ sb_7__0_/right_bottom_grid_pin_11_ cbx_8__0_/bottom_grid_pin_12_
+ sb_8__0_/left_bottom_grid_pin_13_ sb_7__0_/right_bottom_grid_pin_13_ cbx_8__0_/bottom_grid_pin_14_
+ sb_8__0_/left_bottom_grid_pin_15_ sb_7__0_/right_bottom_grid_pin_15_ cbx_8__0_/bottom_grid_pin_16_
+ sb_8__0_/left_bottom_grid_pin_17_ sb_7__0_/right_bottom_grid_pin_17_ sb_8__0_/left_bottom_grid_pin_1_
+ sb_7__0_/right_bottom_grid_pin_1_ cbx_8__0_/bottom_grid_pin_2_ sb_8__0_/left_bottom_grid_pin_3_
+ sb_7__0_/right_bottom_grid_pin_3_ cbx_8__0_/bottom_grid_pin_4_ sb_8__0_/left_bottom_grid_pin_5_
+ sb_7__0_/right_bottom_grid_pin_5_ cbx_8__0_/bottom_grid_pin_6_ sb_8__0_/left_bottom_grid_pin_7_
+ sb_7__0_/right_bottom_grid_pin_7_ cbx_8__0_/bottom_grid_pin_8_ sb_8__0_/left_bottom_grid_pin_9_
+ sb_7__0_/right_bottom_grid_pin_9_ cbx_1__0_
Xgrid_clb_3__8_ cbx_3__8_/SC_OUT_BOT cbx_3__7_/SC_IN_TOP grid_clb_3__8_/SC_OUT_TOP
+ cby_3__8_/Test_en_W_out grid_clb_3__8_/Test_en_E_out cby_3__8_/Test_en_W_out cby_2__8_/Test_en_W_in
+ VGND VPWR cbx_3__7_/REGIN_FEEDTHROUGH grid_clb_3__8_/bottom_width_0_height_0__pin_51_
+ cby_2__8_/ccff_tail cby_3__8_/ccff_head cbx_3__7_/clk_1_N_out cbx_3__7_/clk_1_N_out
+ cby_3__8_/prog_clk_0_W_in cbx_3__7_/prog_clk_1_N_out cbx_3__8_/prog_clk_0_S_in cbx_3__7_/prog_clk_1_N_out
+ cbx_3__7_/prog_clk_0_N_in grid_clb_3__8_/prog_clk_0_W_out cby_3__8_/left_grid_pin_16_
+ cby_3__8_/left_grid_pin_17_ cby_3__8_/left_grid_pin_18_ cby_3__8_/left_grid_pin_19_
+ cby_3__8_/left_grid_pin_20_ cby_3__8_/left_grid_pin_21_ cby_3__8_/left_grid_pin_22_
+ cby_3__8_/left_grid_pin_23_ cby_3__8_/left_grid_pin_24_ cby_3__8_/left_grid_pin_25_
+ cby_3__8_/left_grid_pin_26_ cby_3__8_/left_grid_pin_27_ cby_3__8_/left_grid_pin_28_
+ cby_3__8_/left_grid_pin_29_ cby_3__8_/left_grid_pin_30_ cby_3__8_/left_grid_pin_31_
+ sb_3__7_/top_left_grid_pin_42_ sb_3__8_/bottom_left_grid_pin_42_ sb_3__7_/top_left_grid_pin_43_
+ sb_3__8_/bottom_left_grid_pin_43_ sb_3__7_/top_left_grid_pin_44_ sb_3__8_/bottom_left_grid_pin_44_
+ sb_3__7_/top_left_grid_pin_45_ sb_3__8_/bottom_left_grid_pin_45_ sb_3__7_/top_left_grid_pin_46_
+ sb_3__8_/bottom_left_grid_pin_46_ sb_3__7_/top_left_grid_pin_47_ sb_3__8_/bottom_left_grid_pin_47_
+ sb_3__7_/top_left_grid_pin_48_ sb_3__8_/bottom_left_grid_pin_48_ sb_3__7_/top_left_grid_pin_49_
+ sb_3__8_/bottom_left_grid_pin_49_ cbx_3__8_/bottom_grid_pin_0_ cbx_3__8_/bottom_grid_pin_10_
+ cbx_3__8_/bottom_grid_pin_11_ cbx_3__8_/bottom_grid_pin_12_ cbx_3__8_/bottom_grid_pin_13_
+ cbx_3__8_/bottom_grid_pin_14_ cbx_3__8_/bottom_grid_pin_15_ cbx_3__8_/bottom_grid_pin_1_
+ cbx_3__8_/bottom_grid_pin_2_ tie_array/x[2] grid_clb_3__8_/top_width_0_height_0__pin_33_
+ sb_3__8_/left_bottom_grid_pin_34_ sb_2__8_/right_bottom_grid_pin_34_ sb_3__8_/left_bottom_grid_pin_35_
+ sb_2__8_/right_bottom_grid_pin_35_ sb_3__8_/left_bottom_grid_pin_36_ sb_2__8_/right_bottom_grid_pin_36_
+ sb_3__8_/left_bottom_grid_pin_37_ sb_2__8_/right_bottom_grid_pin_37_ sb_3__8_/left_bottom_grid_pin_38_
+ sb_2__8_/right_bottom_grid_pin_38_ sb_3__8_/left_bottom_grid_pin_39_ sb_2__8_/right_bottom_grid_pin_39_
+ cbx_3__8_/bottom_grid_pin_3_ sb_3__8_/left_bottom_grid_pin_40_ sb_2__8_/right_bottom_grid_pin_40_
+ sb_3__8_/left_bottom_grid_pin_41_ sb_2__8_/right_bottom_grid_pin_41_ cbx_3__8_/bottom_grid_pin_4_
+ cbx_3__8_/bottom_grid_pin_5_ cbx_3__8_/bottom_grid_pin_6_ cbx_3__8_/bottom_grid_pin_7_
+ cbx_3__8_/bottom_grid_pin_8_ cbx_3__8_/bottom_grid_pin_9_ grid_clb
Xcbx_1__5_ cbx_1__5_/REGIN_FEEDTHROUGH cbx_1__5_/REGOUT_FEEDTHROUGH cbx_1__5_/SC_IN_BOT
+ cbx_1__5_/SC_IN_TOP cbx_1__5_/SC_OUT_BOT cbx_1__5_/SC_OUT_TOP VGND VPWR cbx_1__5_/bottom_grid_pin_0_
+ cbx_1__5_/bottom_grid_pin_10_ cbx_1__5_/bottom_grid_pin_11_ cbx_1__5_/bottom_grid_pin_12_
+ cbx_1__5_/bottom_grid_pin_13_ cbx_1__5_/bottom_grid_pin_14_ cbx_1__5_/bottom_grid_pin_15_
+ cbx_1__5_/bottom_grid_pin_1_ cbx_1__5_/bottom_grid_pin_2_ cbx_1__5_/bottom_grid_pin_3_
+ cbx_1__5_/bottom_grid_pin_4_ cbx_1__5_/bottom_grid_pin_5_ cbx_1__5_/bottom_grid_pin_6_
+ cbx_1__5_/bottom_grid_pin_7_ cbx_1__5_/bottom_grid_pin_8_ cbx_1__5_/bottom_grid_pin_9_
+ sb_1__5_/ccff_tail sb_0__5_/ccff_head cbx_1__5_/chanx_left_in[0] cbx_1__5_/chanx_left_in[10]
+ cbx_1__5_/chanx_left_in[11] cbx_1__5_/chanx_left_in[12] cbx_1__5_/chanx_left_in[13]
+ cbx_1__5_/chanx_left_in[14] cbx_1__5_/chanx_left_in[15] cbx_1__5_/chanx_left_in[16]
+ cbx_1__5_/chanx_left_in[17] cbx_1__5_/chanx_left_in[18] cbx_1__5_/chanx_left_in[19]
+ cbx_1__5_/chanx_left_in[1] cbx_1__5_/chanx_left_in[2] cbx_1__5_/chanx_left_in[3]
+ cbx_1__5_/chanx_left_in[4] cbx_1__5_/chanx_left_in[5] cbx_1__5_/chanx_left_in[6]
+ cbx_1__5_/chanx_left_in[7] cbx_1__5_/chanx_left_in[8] cbx_1__5_/chanx_left_in[9]
+ sb_0__5_/chanx_right_in[0] sb_0__5_/chanx_right_in[10] sb_0__5_/chanx_right_in[11]
+ sb_0__5_/chanx_right_in[12] sb_0__5_/chanx_right_in[13] sb_0__5_/chanx_right_in[14]
+ sb_0__5_/chanx_right_in[15] sb_0__5_/chanx_right_in[16] sb_0__5_/chanx_right_in[17]
+ sb_0__5_/chanx_right_in[18] sb_0__5_/chanx_right_in[19] sb_0__5_/chanx_right_in[1]
+ sb_0__5_/chanx_right_in[2] sb_0__5_/chanx_right_in[3] sb_0__5_/chanx_right_in[4]
+ sb_0__5_/chanx_right_in[5] sb_0__5_/chanx_right_in[6] sb_0__5_/chanx_right_in[7]
+ sb_0__5_/chanx_right_in[8] sb_0__5_/chanx_right_in[9] sb_1__5_/chanx_left_out[0]
+ sb_1__5_/chanx_left_out[10] sb_1__5_/chanx_left_out[11] sb_1__5_/chanx_left_out[12]
+ sb_1__5_/chanx_left_out[13] sb_1__5_/chanx_left_out[14] sb_1__5_/chanx_left_out[15]
+ sb_1__5_/chanx_left_out[16] sb_1__5_/chanx_left_out[17] sb_1__5_/chanx_left_out[18]
+ sb_1__5_/chanx_left_out[19] sb_1__5_/chanx_left_out[1] sb_1__5_/chanx_left_out[2]
+ sb_1__5_/chanx_left_out[3] sb_1__5_/chanx_left_out[4] sb_1__5_/chanx_left_out[5]
+ sb_1__5_/chanx_left_out[6] sb_1__5_/chanx_left_out[7] sb_1__5_/chanx_left_out[8]
+ sb_1__5_/chanx_left_out[9] sb_1__5_/chanx_left_in[0] sb_1__5_/chanx_left_in[10]
+ sb_1__5_/chanx_left_in[11] sb_1__5_/chanx_left_in[12] sb_1__5_/chanx_left_in[13]
+ sb_1__5_/chanx_left_in[14] sb_1__5_/chanx_left_in[15] sb_1__5_/chanx_left_in[16]
+ sb_1__5_/chanx_left_in[17] sb_1__5_/chanx_left_in[18] sb_1__5_/chanx_left_in[19]
+ sb_1__5_/chanx_left_in[1] sb_1__5_/chanx_left_in[2] sb_1__5_/chanx_left_in[3] sb_1__5_/chanx_left_in[4]
+ sb_1__5_/chanx_left_in[5] sb_1__5_/chanx_left_in[6] sb_1__5_/chanx_left_in[7] sb_1__5_/chanx_left_in[8]
+ sb_1__5_/chanx_left_in[9] cbx_1__5_/clk_1_N_out cbx_1__5_/clk_1_S_out sb_1__5_/clk_1_W_out
+ cbx_1__5_/clk_2_E_out cbx_1__5_/clk_2_W_in cbx_1__5_/clk_2_W_out cbx_1__5_/clk_3_E_out
+ cbx_1__5_/clk_3_W_in cbx_1__5_/clk_3_W_out cbx_1__5_/prog_clk_0_N_in sb_0__5_/prog_clk_0_E_in
+ cbx_1__5_/prog_clk_1_N_out cbx_1__5_/prog_clk_1_S_out sb_1__5_/prog_clk_1_W_out
+ cbx_1__5_/prog_clk_2_E_out cbx_1__5_/prog_clk_2_W_in cbx_1__5_/prog_clk_2_W_out
+ cbx_1__5_/prog_clk_3_E_out cbx_1__5_/prog_clk_3_W_in cbx_1__5_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_5__2_ sb_5__2_/Test_en_N_out sb_5__2_/Test_en_S_in VGND VPWR sb_5__2_/bottom_left_grid_pin_42_
+ sb_5__2_/bottom_left_grid_pin_43_ sb_5__2_/bottom_left_grid_pin_44_ sb_5__2_/bottom_left_grid_pin_45_
+ sb_5__2_/bottom_left_grid_pin_46_ sb_5__2_/bottom_left_grid_pin_47_ sb_5__2_/bottom_left_grid_pin_48_
+ sb_5__2_/bottom_left_grid_pin_49_ sb_5__2_/ccff_head sb_5__2_/ccff_tail sb_5__2_/chanx_left_in[0]
+ sb_5__2_/chanx_left_in[10] sb_5__2_/chanx_left_in[11] sb_5__2_/chanx_left_in[12]
+ sb_5__2_/chanx_left_in[13] sb_5__2_/chanx_left_in[14] sb_5__2_/chanx_left_in[15]
+ sb_5__2_/chanx_left_in[16] sb_5__2_/chanx_left_in[17] sb_5__2_/chanx_left_in[18]
+ sb_5__2_/chanx_left_in[19] sb_5__2_/chanx_left_in[1] sb_5__2_/chanx_left_in[2] sb_5__2_/chanx_left_in[3]
+ sb_5__2_/chanx_left_in[4] sb_5__2_/chanx_left_in[5] sb_5__2_/chanx_left_in[6] sb_5__2_/chanx_left_in[7]
+ sb_5__2_/chanx_left_in[8] sb_5__2_/chanx_left_in[9] sb_5__2_/chanx_left_out[0] sb_5__2_/chanx_left_out[10]
+ sb_5__2_/chanx_left_out[11] sb_5__2_/chanx_left_out[12] sb_5__2_/chanx_left_out[13]
+ sb_5__2_/chanx_left_out[14] sb_5__2_/chanx_left_out[15] sb_5__2_/chanx_left_out[16]
+ sb_5__2_/chanx_left_out[17] sb_5__2_/chanx_left_out[18] sb_5__2_/chanx_left_out[19]
+ sb_5__2_/chanx_left_out[1] sb_5__2_/chanx_left_out[2] sb_5__2_/chanx_left_out[3]
+ sb_5__2_/chanx_left_out[4] sb_5__2_/chanx_left_out[5] sb_5__2_/chanx_left_out[6]
+ sb_5__2_/chanx_left_out[7] sb_5__2_/chanx_left_out[8] sb_5__2_/chanx_left_out[9]
+ sb_5__2_/chanx_right_in[0] sb_5__2_/chanx_right_in[10] sb_5__2_/chanx_right_in[11]
+ sb_5__2_/chanx_right_in[12] sb_5__2_/chanx_right_in[13] sb_5__2_/chanx_right_in[14]
+ sb_5__2_/chanx_right_in[15] sb_5__2_/chanx_right_in[16] sb_5__2_/chanx_right_in[17]
+ sb_5__2_/chanx_right_in[18] sb_5__2_/chanx_right_in[19] sb_5__2_/chanx_right_in[1]
+ sb_5__2_/chanx_right_in[2] sb_5__2_/chanx_right_in[3] sb_5__2_/chanx_right_in[4]
+ sb_5__2_/chanx_right_in[5] sb_5__2_/chanx_right_in[6] sb_5__2_/chanx_right_in[7]
+ sb_5__2_/chanx_right_in[8] sb_5__2_/chanx_right_in[9] cbx_6__2_/chanx_left_in[0]
+ cbx_6__2_/chanx_left_in[10] cbx_6__2_/chanx_left_in[11] cbx_6__2_/chanx_left_in[12]
+ cbx_6__2_/chanx_left_in[13] cbx_6__2_/chanx_left_in[14] cbx_6__2_/chanx_left_in[15]
+ cbx_6__2_/chanx_left_in[16] cbx_6__2_/chanx_left_in[17] cbx_6__2_/chanx_left_in[18]
+ cbx_6__2_/chanx_left_in[19] cbx_6__2_/chanx_left_in[1] cbx_6__2_/chanx_left_in[2]
+ cbx_6__2_/chanx_left_in[3] cbx_6__2_/chanx_left_in[4] cbx_6__2_/chanx_left_in[5]
+ cbx_6__2_/chanx_left_in[6] cbx_6__2_/chanx_left_in[7] cbx_6__2_/chanx_left_in[8]
+ cbx_6__2_/chanx_left_in[9] cby_5__2_/chany_top_out[0] cby_5__2_/chany_top_out[10]
+ cby_5__2_/chany_top_out[11] cby_5__2_/chany_top_out[12] cby_5__2_/chany_top_out[13]
+ cby_5__2_/chany_top_out[14] cby_5__2_/chany_top_out[15] cby_5__2_/chany_top_out[16]
+ cby_5__2_/chany_top_out[17] cby_5__2_/chany_top_out[18] cby_5__2_/chany_top_out[19]
+ cby_5__2_/chany_top_out[1] cby_5__2_/chany_top_out[2] cby_5__2_/chany_top_out[3]
+ cby_5__2_/chany_top_out[4] cby_5__2_/chany_top_out[5] cby_5__2_/chany_top_out[6]
+ cby_5__2_/chany_top_out[7] cby_5__2_/chany_top_out[8] cby_5__2_/chany_top_out[9]
+ cby_5__2_/chany_top_in[0] cby_5__2_/chany_top_in[10] cby_5__2_/chany_top_in[11]
+ cby_5__2_/chany_top_in[12] cby_5__2_/chany_top_in[13] cby_5__2_/chany_top_in[14]
+ cby_5__2_/chany_top_in[15] cby_5__2_/chany_top_in[16] cby_5__2_/chany_top_in[17]
+ cby_5__2_/chany_top_in[18] cby_5__2_/chany_top_in[19] cby_5__2_/chany_top_in[1]
+ cby_5__2_/chany_top_in[2] cby_5__2_/chany_top_in[3] cby_5__2_/chany_top_in[4] cby_5__2_/chany_top_in[5]
+ cby_5__2_/chany_top_in[6] cby_5__2_/chany_top_in[7] cby_5__2_/chany_top_in[8] cby_5__2_/chany_top_in[9]
+ sb_5__2_/chany_top_in[0] sb_5__2_/chany_top_in[10] sb_5__2_/chany_top_in[11] sb_5__2_/chany_top_in[12]
+ sb_5__2_/chany_top_in[13] sb_5__2_/chany_top_in[14] sb_5__2_/chany_top_in[15] sb_5__2_/chany_top_in[16]
+ sb_5__2_/chany_top_in[17] sb_5__2_/chany_top_in[18] sb_5__2_/chany_top_in[19] sb_5__2_/chany_top_in[1]
+ sb_5__2_/chany_top_in[2] sb_5__2_/chany_top_in[3] sb_5__2_/chany_top_in[4] sb_5__2_/chany_top_in[5]
+ sb_5__2_/chany_top_in[6] sb_5__2_/chany_top_in[7] sb_5__2_/chany_top_in[8] sb_5__2_/chany_top_in[9]
+ sb_5__2_/chany_top_out[0] sb_5__2_/chany_top_out[10] sb_5__2_/chany_top_out[11]
+ sb_5__2_/chany_top_out[12] sb_5__2_/chany_top_out[13] sb_5__2_/chany_top_out[14]
+ sb_5__2_/chany_top_out[15] sb_5__2_/chany_top_out[16] sb_5__2_/chany_top_out[17]
+ sb_5__2_/chany_top_out[18] sb_5__2_/chany_top_out[19] sb_5__2_/chany_top_out[1]
+ sb_5__2_/chany_top_out[2] sb_5__2_/chany_top_out[3] sb_5__2_/chany_top_out[4] sb_5__2_/chany_top_out[5]
+ sb_5__2_/chany_top_out[6] sb_5__2_/chany_top_out[7] sb_5__2_/chany_top_out[8] sb_5__2_/chany_top_out[9]
+ sb_5__2_/clk_1_E_out sb_5__2_/clk_1_N_in sb_5__2_/clk_1_W_out sb_5__2_/clk_2_E_out
+ sb_5__2_/clk_2_N_in sb_5__2_/clk_2_N_out sb_5__2_/clk_2_S_out sb_5__2_/clk_2_W_out
+ sb_5__2_/clk_3_E_out sb_5__2_/clk_3_N_in sb_5__2_/clk_3_N_out sb_5__2_/clk_3_S_out
+ sb_5__2_/clk_3_W_out sb_5__2_/left_bottom_grid_pin_34_ sb_5__2_/left_bottom_grid_pin_35_
+ sb_5__2_/left_bottom_grid_pin_36_ sb_5__2_/left_bottom_grid_pin_37_ sb_5__2_/left_bottom_grid_pin_38_
+ sb_5__2_/left_bottom_grid_pin_39_ sb_5__2_/left_bottom_grid_pin_40_ sb_5__2_/left_bottom_grid_pin_41_
+ sb_5__2_/prog_clk_0_N_in sb_5__2_/prog_clk_1_E_out sb_5__2_/prog_clk_1_N_in sb_5__2_/prog_clk_1_W_out
+ sb_5__2_/prog_clk_2_E_out sb_5__2_/prog_clk_2_N_in sb_5__2_/prog_clk_2_N_out sb_5__2_/prog_clk_2_S_out
+ sb_5__2_/prog_clk_2_W_out sb_5__2_/prog_clk_3_E_out sb_5__2_/prog_clk_3_N_in sb_5__2_/prog_clk_3_N_out
+ sb_5__2_/prog_clk_3_S_out sb_5__2_/prog_clk_3_W_out sb_5__2_/right_bottom_grid_pin_34_
+ sb_5__2_/right_bottom_grid_pin_35_ sb_5__2_/right_bottom_grid_pin_36_ sb_5__2_/right_bottom_grid_pin_37_
+ sb_5__2_/right_bottom_grid_pin_38_ sb_5__2_/right_bottom_grid_pin_39_ sb_5__2_/right_bottom_grid_pin_40_
+ sb_5__2_/right_bottom_grid_pin_41_ sb_5__2_/top_left_grid_pin_42_ sb_5__2_/top_left_grid_pin_43_
+ sb_5__2_/top_left_grid_pin_44_ sb_5__2_/top_left_grid_pin_45_ sb_5__2_/top_left_grid_pin_46_
+ sb_5__2_/top_left_grid_pin_47_ sb_5__2_/top_left_grid_pin_48_ sb_5__2_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_4__6_ sb_4__5_/Test_en_N_out cby_4__6_/Test_en_E_out sb_4__6_/Test_en_S_in sb_4__5_/Test_en_N_out
+ sb_4__5_/Test_en_N_out cby_4__6_/Test_en_W_out VGND VPWR cby_4__6_/ccff_head cby_4__6_/ccff_tail
+ sb_4__5_/chany_top_out[0] sb_4__5_/chany_top_out[10] sb_4__5_/chany_top_out[11]
+ sb_4__5_/chany_top_out[12] sb_4__5_/chany_top_out[13] sb_4__5_/chany_top_out[14]
+ sb_4__5_/chany_top_out[15] sb_4__5_/chany_top_out[16] sb_4__5_/chany_top_out[17]
+ sb_4__5_/chany_top_out[18] sb_4__5_/chany_top_out[19] sb_4__5_/chany_top_out[1]
+ sb_4__5_/chany_top_out[2] sb_4__5_/chany_top_out[3] sb_4__5_/chany_top_out[4] sb_4__5_/chany_top_out[5]
+ sb_4__5_/chany_top_out[6] sb_4__5_/chany_top_out[7] sb_4__5_/chany_top_out[8] sb_4__5_/chany_top_out[9]
+ sb_4__5_/chany_top_in[0] sb_4__5_/chany_top_in[10] sb_4__5_/chany_top_in[11] sb_4__5_/chany_top_in[12]
+ sb_4__5_/chany_top_in[13] sb_4__5_/chany_top_in[14] sb_4__5_/chany_top_in[15] sb_4__5_/chany_top_in[16]
+ sb_4__5_/chany_top_in[17] sb_4__5_/chany_top_in[18] sb_4__5_/chany_top_in[19] sb_4__5_/chany_top_in[1]
+ sb_4__5_/chany_top_in[2] sb_4__5_/chany_top_in[3] sb_4__5_/chany_top_in[4] sb_4__5_/chany_top_in[5]
+ sb_4__5_/chany_top_in[6] sb_4__5_/chany_top_in[7] sb_4__5_/chany_top_in[8] sb_4__5_/chany_top_in[9]
+ cby_4__6_/chany_top_in[0] cby_4__6_/chany_top_in[10] cby_4__6_/chany_top_in[11]
+ cby_4__6_/chany_top_in[12] cby_4__6_/chany_top_in[13] cby_4__6_/chany_top_in[14]
+ cby_4__6_/chany_top_in[15] cby_4__6_/chany_top_in[16] cby_4__6_/chany_top_in[17]
+ cby_4__6_/chany_top_in[18] cby_4__6_/chany_top_in[19] cby_4__6_/chany_top_in[1]
+ cby_4__6_/chany_top_in[2] cby_4__6_/chany_top_in[3] cby_4__6_/chany_top_in[4] cby_4__6_/chany_top_in[5]
+ cby_4__6_/chany_top_in[6] cby_4__6_/chany_top_in[7] cby_4__6_/chany_top_in[8] cby_4__6_/chany_top_in[9]
+ cby_4__6_/chany_top_out[0] cby_4__6_/chany_top_out[10] cby_4__6_/chany_top_out[11]
+ cby_4__6_/chany_top_out[12] cby_4__6_/chany_top_out[13] cby_4__6_/chany_top_out[14]
+ cby_4__6_/chany_top_out[15] cby_4__6_/chany_top_out[16] cby_4__6_/chany_top_out[17]
+ cby_4__6_/chany_top_out[18] cby_4__6_/chany_top_out[19] cby_4__6_/chany_top_out[1]
+ cby_4__6_/chany_top_out[2] cby_4__6_/chany_top_out[3] cby_4__6_/chany_top_out[4]
+ cby_4__6_/chany_top_out[5] cby_4__6_/chany_top_out[6] cby_4__6_/chany_top_out[7]
+ cby_4__6_/chany_top_out[8] cby_4__6_/chany_top_out[9] cby_4__6_/clk_2_N_out cby_4__6_/clk_2_S_in
+ cby_4__6_/clk_2_S_out cby_4__6_/clk_3_N_out cby_4__6_/clk_3_S_in cby_4__6_/clk_3_S_out
+ cby_4__6_/left_grid_pin_16_ cby_4__6_/left_grid_pin_17_ cby_4__6_/left_grid_pin_18_
+ cby_4__6_/left_grid_pin_19_ cby_4__6_/left_grid_pin_20_ cby_4__6_/left_grid_pin_21_
+ cby_4__6_/left_grid_pin_22_ cby_4__6_/left_grid_pin_23_ cby_4__6_/left_grid_pin_24_
+ cby_4__6_/left_grid_pin_25_ cby_4__6_/left_grid_pin_26_ cby_4__6_/left_grid_pin_27_
+ cby_4__6_/left_grid_pin_28_ cby_4__6_/left_grid_pin_29_ cby_4__6_/left_grid_pin_30_
+ cby_4__6_/left_grid_pin_31_ cby_4__6_/prog_clk_0_N_out sb_4__5_/prog_clk_0_N_in
+ cby_4__6_/prog_clk_0_W_in cby_4__6_/prog_clk_2_N_out cby_4__6_/prog_clk_2_S_in cby_4__6_/prog_clk_2_S_out
+ cby_4__6_/prog_clk_3_N_out cby_4__6_/prog_clk_3_S_in cby_4__6_/prog_clk_3_S_out
+ cby_1__1_
Xcby_1__3_ cby_1__3_/Test_en_W_in cby_1__3_/Test_en_E_out cby_1__3_/Test_en_N_out
+ cby_1__3_/Test_en_W_in cby_1__3_/Test_en_W_in cby_1__3_/Test_en_W_out VGND VPWR
+ cby_1__3_/ccff_head cby_1__3_/ccff_tail sb_1__2_/chany_top_out[0] sb_1__2_/chany_top_out[10]
+ sb_1__2_/chany_top_out[11] sb_1__2_/chany_top_out[12] sb_1__2_/chany_top_out[13]
+ sb_1__2_/chany_top_out[14] sb_1__2_/chany_top_out[15] sb_1__2_/chany_top_out[16]
+ sb_1__2_/chany_top_out[17] sb_1__2_/chany_top_out[18] sb_1__2_/chany_top_out[19]
+ sb_1__2_/chany_top_out[1] sb_1__2_/chany_top_out[2] sb_1__2_/chany_top_out[3] sb_1__2_/chany_top_out[4]
+ sb_1__2_/chany_top_out[5] sb_1__2_/chany_top_out[6] sb_1__2_/chany_top_out[7] sb_1__2_/chany_top_out[8]
+ sb_1__2_/chany_top_out[9] sb_1__2_/chany_top_in[0] sb_1__2_/chany_top_in[10] sb_1__2_/chany_top_in[11]
+ sb_1__2_/chany_top_in[12] sb_1__2_/chany_top_in[13] sb_1__2_/chany_top_in[14] sb_1__2_/chany_top_in[15]
+ sb_1__2_/chany_top_in[16] sb_1__2_/chany_top_in[17] sb_1__2_/chany_top_in[18] sb_1__2_/chany_top_in[19]
+ sb_1__2_/chany_top_in[1] sb_1__2_/chany_top_in[2] sb_1__2_/chany_top_in[3] sb_1__2_/chany_top_in[4]
+ sb_1__2_/chany_top_in[5] sb_1__2_/chany_top_in[6] sb_1__2_/chany_top_in[7] sb_1__2_/chany_top_in[8]
+ sb_1__2_/chany_top_in[9] cby_1__3_/chany_top_in[0] cby_1__3_/chany_top_in[10] cby_1__3_/chany_top_in[11]
+ cby_1__3_/chany_top_in[12] cby_1__3_/chany_top_in[13] cby_1__3_/chany_top_in[14]
+ cby_1__3_/chany_top_in[15] cby_1__3_/chany_top_in[16] cby_1__3_/chany_top_in[17]
+ cby_1__3_/chany_top_in[18] cby_1__3_/chany_top_in[19] cby_1__3_/chany_top_in[1]
+ cby_1__3_/chany_top_in[2] cby_1__3_/chany_top_in[3] cby_1__3_/chany_top_in[4] cby_1__3_/chany_top_in[5]
+ cby_1__3_/chany_top_in[6] cby_1__3_/chany_top_in[7] cby_1__3_/chany_top_in[8] cby_1__3_/chany_top_in[9]
+ cby_1__3_/chany_top_out[0] cby_1__3_/chany_top_out[10] cby_1__3_/chany_top_out[11]
+ cby_1__3_/chany_top_out[12] cby_1__3_/chany_top_out[13] cby_1__3_/chany_top_out[14]
+ cby_1__3_/chany_top_out[15] cby_1__3_/chany_top_out[16] cby_1__3_/chany_top_out[17]
+ cby_1__3_/chany_top_out[18] cby_1__3_/chany_top_out[19] cby_1__3_/chany_top_out[1]
+ cby_1__3_/chany_top_out[2] cby_1__3_/chany_top_out[3] cby_1__3_/chany_top_out[4]
+ cby_1__3_/chany_top_out[5] cby_1__3_/chany_top_out[6] cby_1__3_/chany_top_out[7]
+ cby_1__3_/chany_top_out[8] cby_1__3_/chany_top_out[9] sb_1__3_/clk_1_N_in sb_1__2_/clk_2_N_out
+ cby_1__3_/clk_2_S_out cby_1__3_/clk_3_N_out cby_1__3_/clk_3_S_in cby_1__3_/clk_3_S_out
+ cby_1__3_/left_grid_pin_16_ cby_1__3_/left_grid_pin_17_ cby_1__3_/left_grid_pin_18_
+ cby_1__3_/left_grid_pin_19_ cby_1__3_/left_grid_pin_20_ cby_1__3_/left_grid_pin_21_
+ cby_1__3_/left_grid_pin_22_ cby_1__3_/left_grid_pin_23_ cby_1__3_/left_grid_pin_24_
+ cby_1__3_/left_grid_pin_25_ cby_1__3_/left_grid_pin_26_ cby_1__3_/left_grid_pin_27_
+ cby_1__3_/left_grid_pin_28_ cby_1__3_/left_grid_pin_29_ cby_1__3_/left_grid_pin_30_
+ cby_1__3_/left_grid_pin_31_ cby_1__3_/prog_clk_0_N_out sb_1__2_/prog_clk_0_N_in
+ cby_1__3_/prog_clk_0_W_in sb_1__3_/prog_clk_1_N_in sb_1__2_/prog_clk_2_N_out cby_1__3_/prog_clk_2_S_out
+ cby_1__3_/prog_clk_3_N_out cby_1__3_/prog_clk_3_S_in cby_1__3_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_4__7_ cbx_4__7_/REGIN_FEEDTHROUGH cbx_4__7_/REGOUT_FEEDTHROUGH cbx_4__7_/SC_IN_BOT
+ cbx_4__7_/SC_IN_TOP cbx_4__7_/SC_OUT_BOT cbx_4__7_/SC_OUT_TOP VGND VPWR cbx_4__7_/bottom_grid_pin_0_
+ cbx_4__7_/bottom_grid_pin_10_ cbx_4__7_/bottom_grid_pin_11_ cbx_4__7_/bottom_grid_pin_12_
+ cbx_4__7_/bottom_grid_pin_13_ cbx_4__7_/bottom_grid_pin_14_ cbx_4__7_/bottom_grid_pin_15_
+ cbx_4__7_/bottom_grid_pin_1_ cbx_4__7_/bottom_grid_pin_2_ cbx_4__7_/bottom_grid_pin_3_
+ cbx_4__7_/bottom_grid_pin_4_ cbx_4__7_/bottom_grid_pin_5_ cbx_4__7_/bottom_grid_pin_6_
+ cbx_4__7_/bottom_grid_pin_7_ cbx_4__7_/bottom_grid_pin_8_ cbx_4__7_/bottom_grid_pin_9_
+ sb_4__7_/ccff_tail sb_3__7_/ccff_head cbx_4__7_/chanx_left_in[0] cbx_4__7_/chanx_left_in[10]
+ cbx_4__7_/chanx_left_in[11] cbx_4__7_/chanx_left_in[12] cbx_4__7_/chanx_left_in[13]
+ cbx_4__7_/chanx_left_in[14] cbx_4__7_/chanx_left_in[15] cbx_4__7_/chanx_left_in[16]
+ cbx_4__7_/chanx_left_in[17] cbx_4__7_/chanx_left_in[18] cbx_4__7_/chanx_left_in[19]
+ cbx_4__7_/chanx_left_in[1] cbx_4__7_/chanx_left_in[2] cbx_4__7_/chanx_left_in[3]
+ cbx_4__7_/chanx_left_in[4] cbx_4__7_/chanx_left_in[5] cbx_4__7_/chanx_left_in[6]
+ cbx_4__7_/chanx_left_in[7] cbx_4__7_/chanx_left_in[8] cbx_4__7_/chanx_left_in[9]
+ sb_3__7_/chanx_right_in[0] sb_3__7_/chanx_right_in[10] sb_3__7_/chanx_right_in[11]
+ sb_3__7_/chanx_right_in[12] sb_3__7_/chanx_right_in[13] sb_3__7_/chanx_right_in[14]
+ sb_3__7_/chanx_right_in[15] sb_3__7_/chanx_right_in[16] sb_3__7_/chanx_right_in[17]
+ sb_3__7_/chanx_right_in[18] sb_3__7_/chanx_right_in[19] sb_3__7_/chanx_right_in[1]
+ sb_3__7_/chanx_right_in[2] sb_3__7_/chanx_right_in[3] sb_3__7_/chanx_right_in[4]
+ sb_3__7_/chanx_right_in[5] sb_3__7_/chanx_right_in[6] sb_3__7_/chanx_right_in[7]
+ sb_3__7_/chanx_right_in[8] sb_3__7_/chanx_right_in[9] sb_4__7_/chanx_left_out[0]
+ sb_4__7_/chanx_left_out[10] sb_4__7_/chanx_left_out[11] sb_4__7_/chanx_left_out[12]
+ sb_4__7_/chanx_left_out[13] sb_4__7_/chanx_left_out[14] sb_4__7_/chanx_left_out[15]
+ sb_4__7_/chanx_left_out[16] sb_4__7_/chanx_left_out[17] sb_4__7_/chanx_left_out[18]
+ sb_4__7_/chanx_left_out[19] sb_4__7_/chanx_left_out[1] sb_4__7_/chanx_left_out[2]
+ sb_4__7_/chanx_left_out[3] sb_4__7_/chanx_left_out[4] sb_4__7_/chanx_left_out[5]
+ sb_4__7_/chanx_left_out[6] sb_4__7_/chanx_left_out[7] sb_4__7_/chanx_left_out[8]
+ sb_4__7_/chanx_left_out[9] sb_4__7_/chanx_left_in[0] sb_4__7_/chanx_left_in[10]
+ sb_4__7_/chanx_left_in[11] sb_4__7_/chanx_left_in[12] sb_4__7_/chanx_left_in[13]
+ sb_4__7_/chanx_left_in[14] sb_4__7_/chanx_left_in[15] sb_4__7_/chanx_left_in[16]
+ sb_4__7_/chanx_left_in[17] sb_4__7_/chanx_left_in[18] sb_4__7_/chanx_left_in[19]
+ sb_4__7_/chanx_left_in[1] sb_4__7_/chanx_left_in[2] sb_4__7_/chanx_left_in[3] sb_4__7_/chanx_left_in[4]
+ sb_4__7_/chanx_left_in[5] sb_4__7_/chanx_left_in[6] sb_4__7_/chanx_left_in[7] sb_4__7_/chanx_left_in[8]
+ sb_4__7_/chanx_left_in[9] cbx_4__7_/clk_1_N_out cbx_4__7_/clk_1_S_out sb_3__7_/clk_1_E_out
+ cbx_4__7_/clk_2_E_out cbx_4__7_/clk_2_W_in cbx_4__7_/clk_2_W_out cbx_4__7_/clk_3_E_out
+ cbx_4__7_/clk_3_W_in cbx_4__7_/clk_3_W_out cbx_4__7_/prog_clk_0_N_in cbx_4__7_/prog_clk_0_W_out
+ cbx_4__7_/prog_clk_1_N_out cbx_4__7_/prog_clk_1_S_out sb_3__7_/prog_clk_1_E_out
+ cbx_4__7_/prog_clk_2_E_out cbx_4__7_/prog_clk_2_W_in cbx_4__7_/prog_clk_2_W_out
+ cbx_4__7_/prog_clk_3_E_out cbx_4__7_/prog_clk_3_W_in cbx_4__7_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_3__7_ cbx_3__7_/SC_OUT_BOT cbx_3__6_/SC_IN_TOP grid_clb_3__7_/SC_OUT_TOP
+ cby_3__7_/Test_en_W_out grid_clb_3__7_/Test_en_E_out cby_3__7_/Test_en_W_out cby_2__7_/Test_en_W_in
+ VGND VPWR cbx_3__6_/REGIN_FEEDTHROUGH grid_clb_3__7_/bottom_width_0_height_0__pin_51_
+ cby_2__7_/ccff_tail cby_3__7_/ccff_head cbx_3__7_/clk_1_S_out cbx_3__7_/clk_1_S_out
+ cby_3__7_/prog_clk_0_W_in cbx_3__7_/prog_clk_1_S_out grid_clb_3__7_/prog_clk_0_N_out
+ cbx_3__7_/prog_clk_1_S_out cbx_3__6_/prog_clk_0_N_in grid_clb_3__7_/prog_clk_0_W_out
+ cby_3__7_/left_grid_pin_16_ cby_3__7_/left_grid_pin_17_ cby_3__7_/left_grid_pin_18_
+ cby_3__7_/left_grid_pin_19_ cby_3__7_/left_grid_pin_20_ cby_3__7_/left_grid_pin_21_
+ cby_3__7_/left_grid_pin_22_ cby_3__7_/left_grid_pin_23_ cby_3__7_/left_grid_pin_24_
+ cby_3__7_/left_grid_pin_25_ cby_3__7_/left_grid_pin_26_ cby_3__7_/left_grid_pin_27_
+ cby_3__7_/left_grid_pin_28_ cby_3__7_/left_grid_pin_29_ cby_3__7_/left_grid_pin_30_
+ cby_3__7_/left_grid_pin_31_ sb_3__6_/top_left_grid_pin_42_ sb_3__7_/bottom_left_grid_pin_42_
+ sb_3__6_/top_left_grid_pin_43_ sb_3__7_/bottom_left_grid_pin_43_ sb_3__6_/top_left_grid_pin_44_
+ sb_3__7_/bottom_left_grid_pin_44_ sb_3__6_/top_left_grid_pin_45_ sb_3__7_/bottom_left_grid_pin_45_
+ sb_3__6_/top_left_grid_pin_46_ sb_3__7_/bottom_left_grid_pin_46_ sb_3__6_/top_left_grid_pin_47_
+ sb_3__7_/bottom_left_grid_pin_47_ sb_3__6_/top_left_grid_pin_48_ sb_3__7_/bottom_left_grid_pin_48_
+ sb_3__6_/top_left_grid_pin_49_ sb_3__7_/bottom_left_grid_pin_49_ cbx_3__7_/bottom_grid_pin_0_
+ cbx_3__7_/bottom_grid_pin_10_ cbx_3__7_/bottom_grid_pin_11_ cbx_3__7_/bottom_grid_pin_12_
+ cbx_3__7_/bottom_grid_pin_13_ cbx_3__7_/bottom_grid_pin_14_ cbx_3__7_/bottom_grid_pin_15_
+ cbx_3__7_/bottom_grid_pin_1_ cbx_3__7_/bottom_grid_pin_2_ cbx_3__7_/REGOUT_FEEDTHROUGH
+ grid_clb_3__7_/top_width_0_height_0__pin_33_ sb_3__7_/left_bottom_grid_pin_34_ sb_2__7_/right_bottom_grid_pin_34_
+ sb_3__7_/left_bottom_grid_pin_35_ sb_2__7_/right_bottom_grid_pin_35_ sb_3__7_/left_bottom_grid_pin_36_
+ sb_2__7_/right_bottom_grid_pin_36_ sb_3__7_/left_bottom_grid_pin_37_ sb_2__7_/right_bottom_grid_pin_37_
+ sb_3__7_/left_bottom_grid_pin_38_ sb_2__7_/right_bottom_grid_pin_38_ sb_3__7_/left_bottom_grid_pin_39_
+ sb_2__7_/right_bottom_grid_pin_39_ cbx_3__7_/bottom_grid_pin_3_ sb_3__7_/left_bottom_grid_pin_40_
+ sb_2__7_/right_bottom_grid_pin_40_ sb_3__7_/left_bottom_grid_pin_41_ sb_2__7_/right_bottom_grid_pin_41_
+ cbx_3__7_/bottom_grid_pin_4_ cbx_3__7_/bottom_grid_pin_5_ cbx_3__7_/bottom_grid_pin_6_
+ cbx_3__7_/bottom_grid_pin_7_ cbx_3__7_/bottom_grid_pin_8_ cbx_3__7_/bottom_grid_pin_9_
+ grid_clb
Xsb_8__4_ VGND VPWR sb_8__4_/bottom_left_grid_pin_42_ sb_8__4_/bottom_left_grid_pin_43_
+ sb_8__4_/bottom_left_grid_pin_44_ sb_8__4_/bottom_left_grid_pin_45_ sb_8__4_/bottom_left_grid_pin_46_
+ sb_8__4_/bottom_left_grid_pin_47_ sb_8__4_/bottom_left_grid_pin_48_ sb_8__4_/bottom_left_grid_pin_49_
+ sb_8__4_/bottom_right_grid_pin_1_ sb_8__4_/ccff_head sb_8__4_/ccff_tail sb_8__4_/chanx_left_in[0]
+ sb_8__4_/chanx_left_in[10] sb_8__4_/chanx_left_in[11] sb_8__4_/chanx_left_in[12]
+ sb_8__4_/chanx_left_in[13] sb_8__4_/chanx_left_in[14] sb_8__4_/chanx_left_in[15]
+ sb_8__4_/chanx_left_in[16] sb_8__4_/chanx_left_in[17] sb_8__4_/chanx_left_in[18]
+ sb_8__4_/chanx_left_in[19] sb_8__4_/chanx_left_in[1] sb_8__4_/chanx_left_in[2] sb_8__4_/chanx_left_in[3]
+ sb_8__4_/chanx_left_in[4] sb_8__4_/chanx_left_in[5] sb_8__4_/chanx_left_in[6] sb_8__4_/chanx_left_in[7]
+ sb_8__4_/chanx_left_in[8] sb_8__4_/chanx_left_in[9] sb_8__4_/chanx_left_out[0] sb_8__4_/chanx_left_out[10]
+ sb_8__4_/chanx_left_out[11] sb_8__4_/chanx_left_out[12] sb_8__4_/chanx_left_out[13]
+ sb_8__4_/chanx_left_out[14] sb_8__4_/chanx_left_out[15] sb_8__4_/chanx_left_out[16]
+ sb_8__4_/chanx_left_out[17] sb_8__4_/chanx_left_out[18] sb_8__4_/chanx_left_out[19]
+ sb_8__4_/chanx_left_out[1] sb_8__4_/chanx_left_out[2] sb_8__4_/chanx_left_out[3]
+ sb_8__4_/chanx_left_out[4] sb_8__4_/chanx_left_out[5] sb_8__4_/chanx_left_out[6]
+ sb_8__4_/chanx_left_out[7] sb_8__4_/chanx_left_out[8] sb_8__4_/chanx_left_out[9]
+ cby_8__4_/chany_top_out[0] cby_8__4_/chany_top_out[10] cby_8__4_/chany_top_out[11]
+ cby_8__4_/chany_top_out[12] cby_8__4_/chany_top_out[13] cby_8__4_/chany_top_out[14]
+ cby_8__4_/chany_top_out[15] cby_8__4_/chany_top_out[16] cby_8__4_/chany_top_out[17]
+ cby_8__4_/chany_top_out[18] cby_8__4_/chany_top_out[19] cby_8__4_/chany_top_out[1]
+ cby_8__4_/chany_top_out[2] cby_8__4_/chany_top_out[3] cby_8__4_/chany_top_out[4]
+ cby_8__4_/chany_top_out[5] cby_8__4_/chany_top_out[6] cby_8__4_/chany_top_out[7]
+ cby_8__4_/chany_top_out[8] cby_8__4_/chany_top_out[9] cby_8__4_/chany_top_in[0]
+ cby_8__4_/chany_top_in[10] cby_8__4_/chany_top_in[11] cby_8__4_/chany_top_in[12]
+ cby_8__4_/chany_top_in[13] cby_8__4_/chany_top_in[14] cby_8__4_/chany_top_in[15]
+ cby_8__4_/chany_top_in[16] cby_8__4_/chany_top_in[17] cby_8__4_/chany_top_in[18]
+ cby_8__4_/chany_top_in[19] cby_8__4_/chany_top_in[1] cby_8__4_/chany_top_in[2] cby_8__4_/chany_top_in[3]
+ cby_8__4_/chany_top_in[4] cby_8__4_/chany_top_in[5] cby_8__4_/chany_top_in[6] cby_8__4_/chany_top_in[7]
+ cby_8__4_/chany_top_in[8] cby_8__4_/chany_top_in[9] sb_8__4_/chany_top_in[0] sb_8__4_/chany_top_in[10]
+ sb_8__4_/chany_top_in[11] sb_8__4_/chany_top_in[12] sb_8__4_/chany_top_in[13] sb_8__4_/chany_top_in[14]
+ sb_8__4_/chany_top_in[15] sb_8__4_/chany_top_in[16] sb_8__4_/chany_top_in[17] sb_8__4_/chany_top_in[18]
+ sb_8__4_/chany_top_in[19] sb_8__4_/chany_top_in[1] sb_8__4_/chany_top_in[2] sb_8__4_/chany_top_in[3]
+ sb_8__4_/chany_top_in[4] sb_8__4_/chany_top_in[5] sb_8__4_/chany_top_in[6] sb_8__4_/chany_top_in[7]
+ sb_8__4_/chany_top_in[8] sb_8__4_/chany_top_in[9] sb_8__4_/chany_top_out[0] sb_8__4_/chany_top_out[10]
+ sb_8__4_/chany_top_out[11] sb_8__4_/chany_top_out[12] sb_8__4_/chany_top_out[13]
+ sb_8__4_/chany_top_out[14] sb_8__4_/chany_top_out[15] sb_8__4_/chany_top_out[16]
+ sb_8__4_/chany_top_out[17] sb_8__4_/chany_top_out[18] sb_8__4_/chany_top_out[19]
+ sb_8__4_/chany_top_out[1] sb_8__4_/chany_top_out[2] sb_8__4_/chany_top_out[3] sb_8__4_/chany_top_out[4]
+ sb_8__4_/chany_top_out[5] sb_8__4_/chany_top_out[6] sb_8__4_/chany_top_out[7] sb_8__4_/chany_top_out[8]
+ sb_8__4_/chany_top_out[9] sb_8__4_/left_bottom_grid_pin_34_ sb_8__4_/left_bottom_grid_pin_35_
+ sb_8__4_/left_bottom_grid_pin_36_ sb_8__4_/left_bottom_grid_pin_37_ sb_8__4_/left_bottom_grid_pin_38_
+ sb_8__4_/left_bottom_grid_pin_39_ sb_8__4_/left_bottom_grid_pin_40_ sb_8__4_/left_bottom_grid_pin_41_
+ sb_8__4_/prog_clk_0_N_in sb_8__4_/top_left_grid_pin_42_ sb_8__4_/top_left_grid_pin_43_
+ sb_8__4_/top_left_grid_pin_44_ sb_8__4_/top_left_grid_pin_45_ sb_8__4_/top_left_grid_pin_46_
+ sb_8__4_/top_left_grid_pin_47_ sb_8__4_/top_left_grid_pin_48_ sb_8__4_/top_left_grid_pin_49_
+ sb_8__4_/top_right_grid_pin_1_ sb_2__1_
Xcbx_1__4_ cbx_1__4_/REGIN_FEEDTHROUGH cbx_1__4_/REGOUT_FEEDTHROUGH cbx_1__4_/SC_IN_BOT
+ cbx_1__4_/SC_IN_TOP cbx_1__4_/SC_OUT_BOT cbx_1__4_/SC_OUT_TOP VGND VPWR cbx_1__4_/bottom_grid_pin_0_
+ cbx_1__4_/bottom_grid_pin_10_ cbx_1__4_/bottom_grid_pin_11_ cbx_1__4_/bottom_grid_pin_12_
+ cbx_1__4_/bottom_grid_pin_13_ cbx_1__4_/bottom_grid_pin_14_ cbx_1__4_/bottom_grid_pin_15_
+ cbx_1__4_/bottom_grid_pin_1_ cbx_1__4_/bottom_grid_pin_2_ cbx_1__4_/bottom_grid_pin_3_
+ cbx_1__4_/bottom_grid_pin_4_ cbx_1__4_/bottom_grid_pin_5_ cbx_1__4_/bottom_grid_pin_6_
+ cbx_1__4_/bottom_grid_pin_7_ cbx_1__4_/bottom_grid_pin_8_ cbx_1__4_/bottom_grid_pin_9_
+ sb_1__4_/ccff_tail sb_0__4_/ccff_head cbx_1__4_/chanx_left_in[0] cbx_1__4_/chanx_left_in[10]
+ cbx_1__4_/chanx_left_in[11] cbx_1__4_/chanx_left_in[12] cbx_1__4_/chanx_left_in[13]
+ cbx_1__4_/chanx_left_in[14] cbx_1__4_/chanx_left_in[15] cbx_1__4_/chanx_left_in[16]
+ cbx_1__4_/chanx_left_in[17] cbx_1__4_/chanx_left_in[18] cbx_1__4_/chanx_left_in[19]
+ cbx_1__4_/chanx_left_in[1] cbx_1__4_/chanx_left_in[2] cbx_1__4_/chanx_left_in[3]
+ cbx_1__4_/chanx_left_in[4] cbx_1__4_/chanx_left_in[5] cbx_1__4_/chanx_left_in[6]
+ cbx_1__4_/chanx_left_in[7] cbx_1__4_/chanx_left_in[8] cbx_1__4_/chanx_left_in[9]
+ sb_0__4_/chanx_right_in[0] sb_0__4_/chanx_right_in[10] sb_0__4_/chanx_right_in[11]
+ sb_0__4_/chanx_right_in[12] sb_0__4_/chanx_right_in[13] sb_0__4_/chanx_right_in[14]
+ sb_0__4_/chanx_right_in[15] sb_0__4_/chanx_right_in[16] sb_0__4_/chanx_right_in[17]
+ sb_0__4_/chanx_right_in[18] sb_0__4_/chanx_right_in[19] sb_0__4_/chanx_right_in[1]
+ sb_0__4_/chanx_right_in[2] sb_0__4_/chanx_right_in[3] sb_0__4_/chanx_right_in[4]
+ sb_0__4_/chanx_right_in[5] sb_0__4_/chanx_right_in[6] sb_0__4_/chanx_right_in[7]
+ sb_0__4_/chanx_right_in[8] sb_0__4_/chanx_right_in[9] sb_1__4_/chanx_left_out[0]
+ sb_1__4_/chanx_left_out[10] sb_1__4_/chanx_left_out[11] sb_1__4_/chanx_left_out[12]
+ sb_1__4_/chanx_left_out[13] sb_1__4_/chanx_left_out[14] sb_1__4_/chanx_left_out[15]
+ sb_1__4_/chanx_left_out[16] sb_1__4_/chanx_left_out[17] sb_1__4_/chanx_left_out[18]
+ sb_1__4_/chanx_left_out[19] sb_1__4_/chanx_left_out[1] sb_1__4_/chanx_left_out[2]
+ sb_1__4_/chanx_left_out[3] sb_1__4_/chanx_left_out[4] sb_1__4_/chanx_left_out[5]
+ sb_1__4_/chanx_left_out[6] sb_1__4_/chanx_left_out[7] sb_1__4_/chanx_left_out[8]
+ sb_1__4_/chanx_left_out[9] sb_1__4_/chanx_left_in[0] sb_1__4_/chanx_left_in[10]
+ sb_1__4_/chanx_left_in[11] sb_1__4_/chanx_left_in[12] sb_1__4_/chanx_left_in[13]
+ sb_1__4_/chanx_left_in[14] sb_1__4_/chanx_left_in[15] sb_1__4_/chanx_left_in[16]
+ sb_1__4_/chanx_left_in[17] sb_1__4_/chanx_left_in[18] sb_1__4_/chanx_left_in[19]
+ sb_1__4_/chanx_left_in[1] sb_1__4_/chanx_left_in[2] sb_1__4_/chanx_left_in[3] sb_1__4_/chanx_left_in[4]
+ sb_1__4_/chanx_left_in[5] sb_1__4_/chanx_left_in[6] sb_1__4_/chanx_left_in[7] sb_1__4_/chanx_left_in[8]
+ sb_1__4_/chanx_left_in[9] cbx_1__4_/clk_1_N_out cbx_1__4_/clk_1_S_out cbx_1__4_/clk_1_W_in
+ cbx_1__4_/clk_2_E_out cbx_1__4_/clk_2_W_in cbx_1__4_/clk_2_W_out cbx_1__4_/clk_3_E_out
+ cbx_1__4_/clk_3_W_in cbx_1__4_/clk_3_W_out cbx_1__4_/prog_clk_0_N_in sb_0__4_/prog_clk_0_E_in
+ cbx_1__4_/prog_clk_1_N_out cbx_1__4_/prog_clk_1_S_out cbx_1__4_/prog_clk_1_W_in
+ cbx_1__4_/prog_clk_2_E_out cbx_1__4_/prog_clk_2_W_in cbx_1__4_/prog_clk_2_W_out
+ cbx_1__4_/prog_clk_3_E_out cbx_1__4_/prog_clk_3_W_in cbx_1__4_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_5__1_ sb_5__1_/Test_en_N_out sb_5__1_/Test_en_S_in VGND VPWR sb_5__1_/bottom_left_grid_pin_42_
+ sb_5__1_/bottom_left_grid_pin_43_ sb_5__1_/bottom_left_grid_pin_44_ sb_5__1_/bottom_left_grid_pin_45_
+ sb_5__1_/bottom_left_grid_pin_46_ sb_5__1_/bottom_left_grid_pin_47_ sb_5__1_/bottom_left_grid_pin_48_
+ sb_5__1_/bottom_left_grid_pin_49_ sb_5__1_/ccff_head sb_5__1_/ccff_tail sb_5__1_/chanx_left_in[0]
+ sb_5__1_/chanx_left_in[10] sb_5__1_/chanx_left_in[11] sb_5__1_/chanx_left_in[12]
+ sb_5__1_/chanx_left_in[13] sb_5__1_/chanx_left_in[14] sb_5__1_/chanx_left_in[15]
+ sb_5__1_/chanx_left_in[16] sb_5__1_/chanx_left_in[17] sb_5__1_/chanx_left_in[18]
+ sb_5__1_/chanx_left_in[19] sb_5__1_/chanx_left_in[1] sb_5__1_/chanx_left_in[2] sb_5__1_/chanx_left_in[3]
+ sb_5__1_/chanx_left_in[4] sb_5__1_/chanx_left_in[5] sb_5__1_/chanx_left_in[6] sb_5__1_/chanx_left_in[7]
+ sb_5__1_/chanx_left_in[8] sb_5__1_/chanx_left_in[9] sb_5__1_/chanx_left_out[0] sb_5__1_/chanx_left_out[10]
+ sb_5__1_/chanx_left_out[11] sb_5__1_/chanx_left_out[12] sb_5__1_/chanx_left_out[13]
+ sb_5__1_/chanx_left_out[14] sb_5__1_/chanx_left_out[15] sb_5__1_/chanx_left_out[16]
+ sb_5__1_/chanx_left_out[17] sb_5__1_/chanx_left_out[18] sb_5__1_/chanx_left_out[19]
+ sb_5__1_/chanx_left_out[1] sb_5__1_/chanx_left_out[2] sb_5__1_/chanx_left_out[3]
+ sb_5__1_/chanx_left_out[4] sb_5__1_/chanx_left_out[5] sb_5__1_/chanx_left_out[6]
+ sb_5__1_/chanx_left_out[7] sb_5__1_/chanx_left_out[8] sb_5__1_/chanx_left_out[9]
+ sb_5__1_/chanx_right_in[0] sb_5__1_/chanx_right_in[10] sb_5__1_/chanx_right_in[11]
+ sb_5__1_/chanx_right_in[12] sb_5__1_/chanx_right_in[13] sb_5__1_/chanx_right_in[14]
+ sb_5__1_/chanx_right_in[15] sb_5__1_/chanx_right_in[16] sb_5__1_/chanx_right_in[17]
+ sb_5__1_/chanx_right_in[18] sb_5__1_/chanx_right_in[19] sb_5__1_/chanx_right_in[1]
+ sb_5__1_/chanx_right_in[2] sb_5__1_/chanx_right_in[3] sb_5__1_/chanx_right_in[4]
+ sb_5__1_/chanx_right_in[5] sb_5__1_/chanx_right_in[6] sb_5__1_/chanx_right_in[7]
+ sb_5__1_/chanx_right_in[8] sb_5__1_/chanx_right_in[9] cbx_6__1_/chanx_left_in[0]
+ cbx_6__1_/chanx_left_in[10] cbx_6__1_/chanx_left_in[11] cbx_6__1_/chanx_left_in[12]
+ cbx_6__1_/chanx_left_in[13] cbx_6__1_/chanx_left_in[14] cbx_6__1_/chanx_left_in[15]
+ cbx_6__1_/chanx_left_in[16] cbx_6__1_/chanx_left_in[17] cbx_6__1_/chanx_left_in[18]
+ cbx_6__1_/chanx_left_in[19] cbx_6__1_/chanx_left_in[1] cbx_6__1_/chanx_left_in[2]
+ cbx_6__1_/chanx_left_in[3] cbx_6__1_/chanx_left_in[4] cbx_6__1_/chanx_left_in[5]
+ cbx_6__1_/chanx_left_in[6] cbx_6__1_/chanx_left_in[7] cbx_6__1_/chanx_left_in[8]
+ cbx_6__1_/chanx_left_in[9] cby_5__1_/chany_top_out[0] cby_5__1_/chany_top_out[10]
+ cby_5__1_/chany_top_out[11] cby_5__1_/chany_top_out[12] cby_5__1_/chany_top_out[13]
+ cby_5__1_/chany_top_out[14] cby_5__1_/chany_top_out[15] cby_5__1_/chany_top_out[16]
+ cby_5__1_/chany_top_out[17] cby_5__1_/chany_top_out[18] cby_5__1_/chany_top_out[19]
+ cby_5__1_/chany_top_out[1] cby_5__1_/chany_top_out[2] cby_5__1_/chany_top_out[3]
+ cby_5__1_/chany_top_out[4] cby_5__1_/chany_top_out[5] cby_5__1_/chany_top_out[6]
+ cby_5__1_/chany_top_out[7] cby_5__1_/chany_top_out[8] cby_5__1_/chany_top_out[9]
+ cby_5__1_/chany_top_in[0] cby_5__1_/chany_top_in[10] cby_5__1_/chany_top_in[11]
+ cby_5__1_/chany_top_in[12] cby_5__1_/chany_top_in[13] cby_5__1_/chany_top_in[14]
+ cby_5__1_/chany_top_in[15] cby_5__1_/chany_top_in[16] cby_5__1_/chany_top_in[17]
+ cby_5__1_/chany_top_in[18] cby_5__1_/chany_top_in[19] cby_5__1_/chany_top_in[1]
+ cby_5__1_/chany_top_in[2] cby_5__1_/chany_top_in[3] cby_5__1_/chany_top_in[4] cby_5__1_/chany_top_in[5]
+ cby_5__1_/chany_top_in[6] cby_5__1_/chany_top_in[7] cby_5__1_/chany_top_in[8] cby_5__1_/chany_top_in[9]
+ sb_5__1_/chany_top_in[0] sb_5__1_/chany_top_in[10] sb_5__1_/chany_top_in[11] sb_5__1_/chany_top_in[12]
+ sb_5__1_/chany_top_in[13] sb_5__1_/chany_top_in[14] sb_5__1_/chany_top_in[15] sb_5__1_/chany_top_in[16]
+ sb_5__1_/chany_top_in[17] sb_5__1_/chany_top_in[18] sb_5__1_/chany_top_in[19] sb_5__1_/chany_top_in[1]
+ sb_5__1_/chany_top_in[2] sb_5__1_/chany_top_in[3] sb_5__1_/chany_top_in[4] sb_5__1_/chany_top_in[5]
+ sb_5__1_/chany_top_in[6] sb_5__1_/chany_top_in[7] sb_5__1_/chany_top_in[8] sb_5__1_/chany_top_in[9]
+ sb_5__1_/chany_top_out[0] sb_5__1_/chany_top_out[10] sb_5__1_/chany_top_out[11]
+ sb_5__1_/chany_top_out[12] sb_5__1_/chany_top_out[13] sb_5__1_/chany_top_out[14]
+ sb_5__1_/chany_top_out[15] sb_5__1_/chany_top_out[16] sb_5__1_/chany_top_out[17]
+ sb_5__1_/chany_top_out[18] sb_5__1_/chany_top_out[19] sb_5__1_/chany_top_out[1]
+ sb_5__1_/chany_top_out[2] sb_5__1_/chany_top_out[3] sb_5__1_/chany_top_out[4] sb_5__1_/chany_top_out[5]
+ sb_5__1_/chany_top_out[6] sb_5__1_/chany_top_out[7] sb_5__1_/chany_top_out[8] sb_5__1_/chany_top_out[9]
+ sb_5__1_/clk_1_E_out sb_5__1_/clk_1_N_in sb_5__1_/clk_1_W_out sb_5__1_/clk_2_E_out
+ sb_5__1_/clk_2_N_in sb_5__1_/clk_2_N_out sb_5__1_/clk_2_S_out sb_5__1_/clk_2_W_out
+ sb_5__1_/clk_3_E_out sb_5__1_/clk_3_N_in sb_5__1_/clk_3_N_out sb_5__1_/clk_3_S_out
+ sb_5__1_/clk_3_W_out sb_5__1_/left_bottom_grid_pin_34_ sb_5__1_/left_bottom_grid_pin_35_
+ sb_5__1_/left_bottom_grid_pin_36_ sb_5__1_/left_bottom_grid_pin_37_ sb_5__1_/left_bottom_grid_pin_38_
+ sb_5__1_/left_bottom_grid_pin_39_ sb_5__1_/left_bottom_grid_pin_40_ sb_5__1_/left_bottom_grid_pin_41_
+ sb_5__1_/prog_clk_0_N_in sb_5__1_/prog_clk_1_E_out sb_5__1_/prog_clk_1_N_in sb_5__1_/prog_clk_1_W_out
+ sb_5__1_/prog_clk_2_E_out sb_5__1_/prog_clk_2_N_in sb_5__1_/prog_clk_2_N_out sb_5__1_/prog_clk_2_S_out
+ sb_5__1_/prog_clk_2_W_out sb_5__1_/prog_clk_3_E_out sb_5__1_/prog_clk_3_N_in sb_5__1_/prog_clk_3_N_out
+ sb_5__1_/prog_clk_3_S_out sb_5__1_/prog_clk_3_W_out sb_5__1_/right_bottom_grid_pin_34_
+ sb_5__1_/right_bottom_grid_pin_35_ sb_5__1_/right_bottom_grid_pin_36_ sb_5__1_/right_bottom_grid_pin_37_
+ sb_5__1_/right_bottom_grid_pin_38_ sb_5__1_/right_bottom_grid_pin_39_ sb_5__1_/right_bottom_grid_pin_40_
+ sb_5__1_/right_bottom_grid_pin_41_ sb_5__1_/top_left_grid_pin_42_ sb_5__1_/top_left_grid_pin_43_
+ sb_5__1_/top_left_grid_pin_44_ sb_5__1_/top_left_grid_pin_45_ sb_5__1_/top_left_grid_pin_46_
+ sb_5__1_/top_left_grid_pin_47_ sb_5__1_/top_left_grid_pin_48_ sb_5__1_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_7__8_ cby_7__8_/Test_en_W_in cby_7__8_/Test_en_E_out cby_7__8_/Test_en_N_out
+ cby_7__8_/Test_en_W_in cby_7__8_/Test_en_W_in cby_7__8_/Test_en_W_out VGND VPWR
+ cby_7__8_/ccff_head cby_7__8_/ccff_tail sb_7__7_/chany_top_out[0] sb_7__7_/chany_top_out[10]
+ sb_7__7_/chany_top_out[11] sb_7__7_/chany_top_out[12] sb_7__7_/chany_top_out[13]
+ sb_7__7_/chany_top_out[14] sb_7__7_/chany_top_out[15] sb_7__7_/chany_top_out[16]
+ sb_7__7_/chany_top_out[17] sb_7__7_/chany_top_out[18] sb_7__7_/chany_top_out[19]
+ sb_7__7_/chany_top_out[1] sb_7__7_/chany_top_out[2] sb_7__7_/chany_top_out[3] sb_7__7_/chany_top_out[4]
+ sb_7__7_/chany_top_out[5] sb_7__7_/chany_top_out[6] sb_7__7_/chany_top_out[7] sb_7__7_/chany_top_out[8]
+ sb_7__7_/chany_top_out[9] sb_7__7_/chany_top_in[0] sb_7__7_/chany_top_in[10] sb_7__7_/chany_top_in[11]
+ sb_7__7_/chany_top_in[12] sb_7__7_/chany_top_in[13] sb_7__7_/chany_top_in[14] sb_7__7_/chany_top_in[15]
+ sb_7__7_/chany_top_in[16] sb_7__7_/chany_top_in[17] sb_7__7_/chany_top_in[18] sb_7__7_/chany_top_in[19]
+ sb_7__7_/chany_top_in[1] sb_7__7_/chany_top_in[2] sb_7__7_/chany_top_in[3] sb_7__7_/chany_top_in[4]
+ sb_7__7_/chany_top_in[5] sb_7__7_/chany_top_in[6] sb_7__7_/chany_top_in[7] sb_7__7_/chany_top_in[8]
+ sb_7__7_/chany_top_in[9] cby_7__8_/chany_top_in[0] cby_7__8_/chany_top_in[10] cby_7__8_/chany_top_in[11]
+ cby_7__8_/chany_top_in[12] cby_7__8_/chany_top_in[13] cby_7__8_/chany_top_in[14]
+ cby_7__8_/chany_top_in[15] cby_7__8_/chany_top_in[16] cby_7__8_/chany_top_in[17]
+ cby_7__8_/chany_top_in[18] cby_7__8_/chany_top_in[19] cby_7__8_/chany_top_in[1]
+ cby_7__8_/chany_top_in[2] cby_7__8_/chany_top_in[3] cby_7__8_/chany_top_in[4] cby_7__8_/chany_top_in[5]
+ cby_7__8_/chany_top_in[6] cby_7__8_/chany_top_in[7] cby_7__8_/chany_top_in[8] cby_7__8_/chany_top_in[9]
+ cby_7__8_/chany_top_out[0] cby_7__8_/chany_top_out[10] cby_7__8_/chany_top_out[11]
+ cby_7__8_/chany_top_out[12] cby_7__8_/chany_top_out[13] cby_7__8_/chany_top_out[14]
+ cby_7__8_/chany_top_out[15] cby_7__8_/chany_top_out[16] cby_7__8_/chany_top_out[17]
+ cby_7__8_/chany_top_out[18] cby_7__8_/chany_top_out[19] cby_7__8_/chany_top_out[1]
+ cby_7__8_/chany_top_out[2] cby_7__8_/chany_top_out[3] cby_7__8_/chany_top_out[4]
+ cby_7__8_/chany_top_out[5] cby_7__8_/chany_top_out[6] cby_7__8_/chany_top_out[7]
+ cby_7__8_/chany_top_out[8] cby_7__8_/chany_top_out[9] cby_7__8_/clk_2_N_out cby_7__8_/clk_2_S_in
+ cby_7__8_/clk_2_S_out cby_7__8_/clk_3_N_out cby_7__8_/clk_3_S_in cby_7__8_/clk_3_S_out
+ cby_7__8_/left_grid_pin_16_ cby_7__8_/left_grid_pin_17_ cby_7__8_/left_grid_pin_18_
+ cby_7__8_/left_grid_pin_19_ cby_7__8_/left_grid_pin_20_ cby_7__8_/left_grid_pin_21_
+ cby_7__8_/left_grid_pin_22_ cby_7__8_/left_grid_pin_23_ cby_7__8_/left_grid_pin_24_
+ cby_7__8_/left_grid_pin_25_ cby_7__8_/left_grid_pin_26_ cby_7__8_/left_grid_pin_27_
+ cby_7__8_/left_grid_pin_28_ cby_7__8_/left_grid_pin_29_ cby_7__8_/left_grid_pin_30_
+ cby_7__8_/left_grid_pin_31_ sb_7__8_/prog_clk_0_S_in sb_7__7_/prog_clk_0_N_in cby_7__8_/prog_clk_0_W_in
+ cby_7__8_/prog_clk_2_N_out cby_7__8_/prog_clk_2_S_in cby_7__8_/prog_clk_2_S_out
+ cby_7__8_/prog_clk_3_N_out cby_7__8_/prog_clk_3_S_in cby_7__8_/prog_clk_3_S_out
+ cby_1__1_
Xcby_4__5_ sb_4__4_/Test_en_N_out cby_4__5_/Test_en_E_out sb_4__5_/Test_en_S_in sb_4__4_/Test_en_N_out
+ sb_4__4_/Test_en_N_out cby_4__5_/Test_en_W_out VGND VPWR cby_4__5_/ccff_head cby_4__5_/ccff_tail
+ sb_4__4_/chany_top_out[0] sb_4__4_/chany_top_out[10] sb_4__4_/chany_top_out[11]
+ sb_4__4_/chany_top_out[12] sb_4__4_/chany_top_out[13] sb_4__4_/chany_top_out[14]
+ sb_4__4_/chany_top_out[15] sb_4__4_/chany_top_out[16] sb_4__4_/chany_top_out[17]
+ sb_4__4_/chany_top_out[18] sb_4__4_/chany_top_out[19] sb_4__4_/chany_top_out[1]
+ sb_4__4_/chany_top_out[2] sb_4__4_/chany_top_out[3] sb_4__4_/chany_top_out[4] sb_4__4_/chany_top_out[5]
+ sb_4__4_/chany_top_out[6] sb_4__4_/chany_top_out[7] sb_4__4_/chany_top_out[8] sb_4__4_/chany_top_out[9]
+ sb_4__4_/chany_top_in[0] sb_4__4_/chany_top_in[10] sb_4__4_/chany_top_in[11] sb_4__4_/chany_top_in[12]
+ sb_4__4_/chany_top_in[13] sb_4__4_/chany_top_in[14] sb_4__4_/chany_top_in[15] sb_4__4_/chany_top_in[16]
+ sb_4__4_/chany_top_in[17] sb_4__4_/chany_top_in[18] sb_4__4_/chany_top_in[19] sb_4__4_/chany_top_in[1]
+ sb_4__4_/chany_top_in[2] sb_4__4_/chany_top_in[3] sb_4__4_/chany_top_in[4] sb_4__4_/chany_top_in[5]
+ sb_4__4_/chany_top_in[6] sb_4__4_/chany_top_in[7] sb_4__4_/chany_top_in[8] sb_4__4_/chany_top_in[9]
+ cby_4__5_/chany_top_in[0] cby_4__5_/chany_top_in[10] cby_4__5_/chany_top_in[11]
+ cby_4__5_/chany_top_in[12] cby_4__5_/chany_top_in[13] cby_4__5_/chany_top_in[14]
+ cby_4__5_/chany_top_in[15] cby_4__5_/chany_top_in[16] cby_4__5_/chany_top_in[17]
+ cby_4__5_/chany_top_in[18] cby_4__5_/chany_top_in[19] cby_4__5_/chany_top_in[1]
+ cby_4__5_/chany_top_in[2] cby_4__5_/chany_top_in[3] cby_4__5_/chany_top_in[4] cby_4__5_/chany_top_in[5]
+ cby_4__5_/chany_top_in[6] cby_4__5_/chany_top_in[7] cby_4__5_/chany_top_in[8] cby_4__5_/chany_top_in[9]
+ cby_4__5_/chany_top_out[0] cby_4__5_/chany_top_out[10] cby_4__5_/chany_top_out[11]
+ cby_4__5_/chany_top_out[12] cby_4__5_/chany_top_out[13] cby_4__5_/chany_top_out[14]
+ cby_4__5_/chany_top_out[15] cby_4__5_/chany_top_out[16] cby_4__5_/chany_top_out[17]
+ cby_4__5_/chany_top_out[18] cby_4__5_/chany_top_out[19] cby_4__5_/chany_top_out[1]
+ cby_4__5_/chany_top_out[2] cby_4__5_/chany_top_out[3] cby_4__5_/chany_top_out[4]
+ cby_4__5_/chany_top_out[5] cby_4__5_/chany_top_out[6] cby_4__5_/chany_top_out[7]
+ cby_4__5_/chany_top_out[8] cby_4__5_/chany_top_out[9] cby_4__5_/clk_2_N_out cby_4__5_/clk_2_S_in
+ cby_4__5_/clk_2_S_out cby_4__5_/clk_3_N_out cby_4__5_/clk_3_S_in cby_4__5_/clk_3_S_out
+ cby_4__5_/left_grid_pin_16_ cby_4__5_/left_grid_pin_17_ cby_4__5_/left_grid_pin_18_
+ cby_4__5_/left_grid_pin_19_ cby_4__5_/left_grid_pin_20_ cby_4__5_/left_grid_pin_21_
+ cby_4__5_/left_grid_pin_22_ cby_4__5_/left_grid_pin_23_ cby_4__5_/left_grid_pin_24_
+ cby_4__5_/left_grid_pin_25_ cby_4__5_/left_grid_pin_26_ cby_4__5_/left_grid_pin_27_
+ cby_4__5_/left_grid_pin_28_ cby_4__5_/left_grid_pin_29_ cby_4__5_/left_grid_pin_30_
+ cby_4__5_/left_grid_pin_31_ cby_4__5_/prog_clk_0_N_out sb_4__4_/prog_clk_0_N_in
+ cby_4__5_/prog_clk_0_W_in cby_4__5_/prog_clk_2_N_out cby_4__5_/prog_clk_2_S_in cby_4__5_/prog_clk_2_S_out
+ cby_4__5_/prog_clk_3_N_out cby_4__5_/prog_clk_3_S_in cby_4__5_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_4__6_ cbx_4__6_/REGIN_FEEDTHROUGH cbx_4__6_/REGOUT_FEEDTHROUGH cbx_4__6_/SC_IN_BOT
+ cbx_4__6_/SC_IN_TOP cbx_4__6_/SC_OUT_BOT cbx_4__6_/SC_OUT_TOP VGND VPWR cbx_4__6_/bottom_grid_pin_0_
+ cbx_4__6_/bottom_grid_pin_10_ cbx_4__6_/bottom_grid_pin_11_ cbx_4__6_/bottom_grid_pin_12_
+ cbx_4__6_/bottom_grid_pin_13_ cbx_4__6_/bottom_grid_pin_14_ cbx_4__6_/bottom_grid_pin_15_
+ cbx_4__6_/bottom_grid_pin_1_ cbx_4__6_/bottom_grid_pin_2_ cbx_4__6_/bottom_grid_pin_3_
+ cbx_4__6_/bottom_grid_pin_4_ cbx_4__6_/bottom_grid_pin_5_ cbx_4__6_/bottom_grid_pin_6_
+ cbx_4__6_/bottom_grid_pin_7_ cbx_4__6_/bottom_grid_pin_8_ cbx_4__6_/bottom_grid_pin_9_
+ sb_4__6_/ccff_tail sb_3__6_/ccff_head cbx_4__6_/chanx_left_in[0] cbx_4__6_/chanx_left_in[10]
+ cbx_4__6_/chanx_left_in[11] cbx_4__6_/chanx_left_in[12] cbx_4__6_/chanx_left_in[13]
+ cbx_4__6_/chanx_left_in[14] cbx_4__6_/chanx_left_in[15] cbx_4__6_/chanx_left_in[16]
+ cbx_4__6_/chanx_left_in[17] cbx_4__6_/chanx_left_in[18] cbx_4__6_/chanx_left_in[19]
+ cbx_4__6_/chanx_left_in[1] cbx_4__6_/chanx_left_in[2] cbx_4__6_/chanx_left_in[3]
+ cbx_4__6_/chanx_left_in[4] cbx_4__6_/chanx_left_in[5] cbx_4__6_/chanx_left_in[6]
+ cbx_4__6_/chanx_left_in[7] cbx_4__6_/chanx_left_in[8] cbx_4__6_/chanx_left_in[9]
+ sb_3__6_/chanx_right_in[0] sb_3__6_/chanx_right_in[10] sb_3__6_/chanx_right_in[11]
+ sb_3__6_/chanx_right_in[12] sb_3__6_/chanx_right_in[13] sb_3__6_/chanx_right_in[14]
+ sb_3__6_/chanx_right_in[15] sb_3__6_/chanx_right_in[16] sb_3__6_/chanx_right_in[17]
+ sb_3__6_/chanx_right_in[18] sb_3__6_/chanx_right_in[19] sb_3__6_/chanx_right_in[1]
+ sb_3__6_/chanx_right_in[2] sb_3__6_/chanx_right_in[3] sb_3__6_/chanx_right_in[4]
+ sb_3__6_/chanx_right_in[5] sb_3__6_/chanx_right_in[6] sb_3__6_/chanx_right_in[7]
+ sb_3__6_/chanx_right_in[8] sb_3__6_/chanx_right_in[9] sb_4__6_/chanx_left_out[0]
+ sb_4__6_/chanx_left_out[10] sb_4__6_/chanx_left_out[11] sb_4__6_/chanx_left_out[12]
+ sb_4__6_/chanx_left_out[13] sb_4__6_/chanx_left_out[14] sb_4__6_/chanx_left_out[15]
+ sb_4__6_/chanx_left_out[16] sb_4__6_/chanx_left_out[17] sb_4__6_/chanx_left_out[18]
+ sb_4__6_/chanx_left_out[19] sb_4__6_/chanx_left_out[1] sb_4__6_/chanx_left_out[2]
+ sb_4__6_/chanx_left_out[3] sb_4__6_/chanx_left_out[4] sb_4__6_/chanx_left_out[5]
+ sb_4__6_/chanx_left_out[6] sb_4__6_/chanx_left_out[7] sb_4__6_/chanx_left_out[8]
+ sb_4__6_/chanx_left_out[9] sb_4__6_/chanx_left_in[0] sb_4__6_/chanx_left_in[10]
+ sb_4__6_/chanx_left_in[11] sb_4__6_/chanx_left_in[12] sb_4__6_/chanx_left_in[13]
+ sb_4__6_/chanx_left_in[14] sb_4__6_/chanx_left_in[15] sb_4__6_/chanx_left_in[16]
+ sb_4__6_/chanx_left_in[17] sb_4__6_/chanx_left_in[18] sb_4__6_/chanx_left_in[19]
+ sb_4__6_/chanx_left_in[1] sb_4__6_/chanx_left_in[2] sb_4__6_/chanx_left_in[3] sb_4__6_/chanx_left_in[4]
+ sb_4__6_/chanx_left_in[5] sb_4__6_/chanx_left_in[6] sb_4__6_/chanx_left_in[7] sb_4__6_/chanx_left_in[8]
+ sb_4__6_/chanx_left_in[9] cbx_4__6_/clk_1_N_out cbx_4__6_/clk_1_S_out cbx_4__6_/clk_1_W_in
+ cbx_4__6_/clk_2_E_out cbx_4__6_/clk_2_W_in cbx_4__6_/clk_2_W_out cbx_4__6_/clk_3_E_out
+ cbx_4__6_/clk_3_W_in cbx_4__6_/clk_3_W_out cbx_4__6_/prog_clk_0_N_in cbx_4__6_/prog_clk_0_W_out
+ cbx_4__6_/prog_clk_1_N_out cbx_4__6_/prog_clk_1_S_out cbx_4__6_/prog_clk_1_W_in
+ cbx_4__6_/prog_clk_2_E_out cbx_4__6_/prog_clk_2_W_in cbx_4__6_/prog_clk_2_W_out
+ cbx_4__6_/prog_clk_3_E_out cbx_4__6_/prog_clk_3_W_in cbx_4__6_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_8__3_ VGND VPWR sb_8__3_/bottom_left_grid_pin_42_ sb_8__3_/bottom_left_grid_pin_43_
+ sb_8__3_/bottom_left_grid_pin_44_ sb_8__3_/bottom_left_grid_pin_45_ sb_8__3_/bottom_left_grid_pin_46_
+ sb_8__3_/bottom_left_grid_pin_47_ sb_8__3_/bottom_left_grid_pin_48_ sb_8__3_/bottom_left_grid_pin_49_
+ sb_8__3_/bottom_right_grid_pin_1_ sb_8__3_/ccff_head sb_8__3_/ccff_tail sb_8__3_/chanx_left_in[0]
+ sb_8__3_/chanx_left_in[10] sb_8__3_/chanx_left_in[11] sb_8__3_/chanx_left_in[12]
+ sb_8__3_/chanx_left_in[13] sb_8__3_/chanx_left_in[14] sb_8__3_/chanx_left_in[15]
+ sb_8__3_/chanx_left_in[16] sb_8__3_/chanx_left_in[17] sb_8__3_/chanx_left_in[18]
+ sb_8__3_/chanx_left_in[19] sb_8__3_/chanx_left_in[1] sb_8__3_/chanx_left_in[2] sb_8__3_/chanx_left_in[3]
+ sb_8__3_/chanx_left_in[4] sb_8__3_/chanx_left_in[5] sb_8__3_/chanx_left_in[6] sb_8__3_/chanx_left_in[7]
+ sb_8__3_/chanx_left_in[8] sb_8__3_/chanx_left_in[9] sb_8__3_/chanx_left_out[0] sb_8__3_/chanx_left_out[10]
+ sb_8__3_/chanx_left_out[11] sb_8__3_/chanx_left_out[12] sb_8__3_/chanx_left_out[13]
+ sb_8__3_/chanx_left_out[14] sb_8__3_/chanx_left_out[15] sb_8__3_/chanx_left_out[16]
+ sb_8__3_/chanx_left_out[17] sb_8__3_/chanx_left_out[18] sb_8__3_/chanx_left_out[19]
+ sb_8__3_/chanx_left_out[1] sb_8__3_/chanx_left_out[2] sb_8__3_/chanx_left_out[3]
+ sb_8__3_/chanx_left_out[4] sb_8__3_/chanx_left_out[5] sb_8__3_/chanx_left_out[6]
+ sb_8__3_/chanx_left_out[7] sb_8__3_/chanx_left_out[8] sb_8__3_/chanx_left_out[9]
+ cby_8__3_/chany_top_out[0] cby_8__3_/chany_top_out[10] cby_8__3_/chany_top_out[11]
+ cby_8__3_/chany_top_out[12] cby_8__3_/chany_top_out[13] cby_8__3_/chany_top_out[14]
+ cby_8__3_/chany_top_out[15] cby_8__3_/chany_top_out[16] cby_8__3_/chany_top_out[17]
+ cby_8__3_/chany_top_out[18] cby_8__3_/chany_top_out[19] cby_8__3_/chany_top_out[1]
+ cby_8__3_/chany_top_out[2] cby_8__3_/chany_top_out[3] cby_8__3_/chany_top_out[4]
+ cby_8__3_/chany_top_out[5] cby_8__3_/chany_top_out[6] cby_8__3_/chany_top_out[7]
+ cby_8__3_/chany_top_out[8] cby_8__3_/chany_top_out[9] cby_8__3_/chany_top_in[0]
+ cby_8__3_/chany_top_in[10] cby_8__3_/chany_top_in[11] cby_8__3_/chany_top_in[12]
+ cby_8__3_/chany_top_in[13] cby_8__3_/chany_top_in[14] cby_8__3_/chany_top_in[15]
+ cby_8__3_/chany_top_in[16] cby_8__3_/chany_top_in[17] cby_8__3_/chany_top_in[18]
+ cby_8__3_/chany_top_in[19] cby_8__3_/chany_top_in[1] cby_8__3_/chany_top_in[2] cby_8__3_/chany_top_in[3]
+ cby_8__3_/chany_top_in[4] cby_8__3_/chany_top_in[5] cby_8__3_/chany_top_in[6] cby_8__3_/chany_top_in[7]
+ cby_8__3_/chany_top_in[8] cby_8__3_/chany_top_in[9] sb_8__3_/chany_top_in[0] sb_8__3_/chany_top_in[10]
+ sb_8__3_/chany_top_in[11] sb_8__3_/chany_top_in[12] sb_8__3_/chany_top_in[13] sb_8__3_/chany_top_in[14]
+ sb_8__3_/chany_top_in[15] sb_8__3_/chany_top_in[16] sb_8__3_/chany_top_in[17] sb_8__3_/chany_top_in[18]
+ sb_8__3_/chany_top_in[19] sb_8__3_/chany_top_in[1] sb_8__3_/chany_top_in[2] sb_8__3_/chany_top_in[3]
+ sb_8__3_/chany_top_in[4] sb_8__3_/chany_top_in[5] sb_8__3_/chany_top_in[6] sb_8__3_/chany_top_in[7]
+ sb_8__3_/chany_top_in[8] sb_8__3_/chany_top_in[9] sb_8__3_/chany_top_out[0] sb_8__3_/chany_top_out[10]
+ sb_8__3_/chany_top_out[11] sb_8__3_/chany_top_out[12] sb_8__3_/chany_top_out[13]
+ sb_8__3_/chany_top_out[14] sb_8__3_/chany_top_out[15] sb_8__3_/chany_top_out[16]
+ sb_8__3_/chany_top_out[17] sb_8__3_/chany_top_out[18] sb_8__3_/chany_top_out[19]
+ sb_8__3_/chany_top_out[1] sb_8__3_/chany_top_out[2] sb_8__3_/chany_top_out[3] sb_8__3_/chany_top_out[4]
+ sb_8__3_/chany_top_out[5] sb_8__3_/chany_top_out[6] sb_8__3_/chany_top_out[7] sb_8__3_/chany_top_out[8]
+ sb_8__3_/chany_top_out[9] sb_8__3_/left_bottom_grid_pin_34_ sb_8__3_/left_bottom_grid_pin_35_
+ sb_8__3_/left_bottom_grid_pin_36_ sb_8__3_/left_bottom_grid_pin_37_ sb_8__3_/left_bottom_grid_pin_38_
+ sb_8__3_/left_bottom_grid_pin_39_ sb_8__3_/left_bottom_grid_pin_40_ sb_8__3_/left_bottom_grid_pin_41_
+ sb_8__3_/prog_clk_0_N_in sb_8__3_/top_left_grid_pin_42_ sb_8__3_/top_left_grid_pin_43_
+ sb_8__3_/top_left_grid_pin_44_ sb_8__3_/top_left_grid_pin_45_ sb_8__3_/top_left_grid_pin_46_
+ sb_8__3_/top_left_grid_pin_47_ sb_8__3_/top_left_grid_pin_48_ sb_8__3_/top_left_grid_pin_49_
+ sb_8__3_/top_right_grid_pin_1_ sb_2__1_
Xcby_1__2_ cby_1__2_/Test_en_W_in cby_1__2_/Test_en_E_out cby_1__2_/Test_en_N_out
+ cby_1__2_/Test_en_W_in cby_1__2_/Test_en_W_in cby_1__2_/Test_en_W_out VGND VPWR
+ cby_1__2_/ccff_head cby_1__2_/ccff_tail sb_1__1_/chany_top_out[0] sb_1__1_/chany_top_out[10]
+ sb_1__1_/chany_top_out[11] sb_1__1_/chany_top_out[12] sb_1__1_/chany_top_out[13]
+ sb_1__1_/chany_top_out[14] sb_1__1_/chany_top_out[15] sb_1__1_/chany_top_out[16]
+ sb_1__1_/chany_top_out[17] sb_1__1_/chany_top_out[18] sb_1__1_/chany_top_out[19]
+ sb_1__1_/chany_top_out[1] sb_1__1_/chany_top_out[2] sb_1__1_/chany_top_out[3] sb_1__1_/chany_top_out[4]
+ sb_1__1_/chany_top_out[5] sb_1__1_/chany_top_out[6] sb_1__1_/chany_top_out[7] sb_1__1_/chany_top_out[8]
+ sb_1__1_/chany_top_out[9] sb_1__1_/chany_top_in[0] sb_1__1_/chany_top_in[10] sb_1__1_/chany_top_in[11]
+ sb_1__1_/chany_top_in[12] sb_1__1_/chany_top_in[13] sb_1__1_/chany_top_in[14] sb_1__1_/chany_top_in[15]
+ sb_1__1_/chany_top_in[16] sb_1__1_/chany_top_in[17] sb_1__1_/chany_top_in[18] sb_1__1_/chany_top_in[19]
+ sb_1__1_/chany_top_in[1] sb_1__1_/chany_top_in[2] sb_1__1_/chany_top_in[3] sb_1__1_/chany_top_in[4]
+ sb_1__1_/chany_top_in[5] sb_1__1_/chany_top_in[6] sb_1__1_/chany_top_in[7] sb_1__1_/chany_top_in[8]
+ sb_1__1_/chany_top_in[9] cby_1__2_/chany_top_in[0] cby_1__2_/chany_top_in[10] cby_1__2_/chany_top_in[11]
+ cby_1__2_/chany_top_in[12] cby_1__2_/chany_top_in[13] cby_1__2_/chany_top_in[14]
+ cby_1__2_/chany_top_in[15] cby_1__2_/chany_top_in[16] cby_1__2_/chany_top_in[17]
+ cby_1__2_/chany_top_in[18] cby_1__2_/chany_top_in[19] cby_1__2_/chany_top_in[1]
+ cby_1__2_/chany_top_in[2] cby_1__2_/chany_top_in[3] cby_1__2_/chany_top_in[4] cby_1__2_/chany_top_in[5]
+ cby_1__2_/chany_top_in[6] cby_1__2_/chany_top_in[7] cby_1__2_/chany_top_in[8] cby_1__2_/chany_top_in[9]
+ cby_1__2_/chany_top_out[0] cby_1__2_/chany_top_out[10] cby_1__2_/chany_top_out[11]
+ cby_1__2_/chany_top_out[12] cby_1__2_/chany_top_out[13] cby_1__2_/chany_top_out[14]
+ cby_1__2_/chany_top_out[15] cby_1__2_/chany_top_out[16] cby_1__2_/chany_top_out[17]
+ cby_1__2_/chany_top_out[18] cby_1__2_/chany_top_out[19] cby_1__2_/chany_top_out[1]
+ cby_1__2_/chany_top_out[2] cby_1__2_/chany_top_out[3] cby_1__2_/chany_top_out[4]
+ cby_1__2_/chany_top_out[5] cby_1__2_/chany_top_out[6] cby_1__2_/chany_top_out[7]
+ cby_1__2_/chany_top_out[8] cby_1__2_/chany_top_out[9] cby_1__2_/clk_2_N_out sb_1__2_/clk_2_S_out
+ sb_1__1_/clk_1_N_in cby_1__2_/clk_3_N_out cby_1__2_/clk_3_S_in cby_1__2_/clk_3_S_out
+ cby_1__2_/left_grid_pin_16_ cby_1__2_/left_grid_pin_17_ cby_1__2_/left_grid_pin_18_
+ cby_1__2_/left_grid_pin_19_ cby_1__2_/left_grid_pin_20_ cby_1__2_/left_grid_pin_21_
+ cby_1__2_/left_grid_pin_22_ cby_1__2_/left_grid_pin_23_ cby_1__2_/left_grid_pin_24_
+ cby_1__2_/left_grid_pin_25_ cby_1__2_/left_grid_pin_26_ cby_1__2_/left_grid_pin_27_
+ cby_1__2_/left_grid_pin_28_ cby_1__2_/left_grid_pin_29_ cby_1__2_/left_grid_pin_30_
+ cby_1__2_/left_grid_pin_31_ cby_1__2_/prog_clk_0_N_out sb_1__1_/prog_clk_0_N_in
+ cby_1__2_/prog_clk_0_W_in cby_1__2_/prog_clk_2_N_out sb_1__2_/prog_clk_2_S_out sb_1__1_/prog_clk_1_N_in
+ cby_1__2_/prog_clk_3_N_out cby_1__2_/prog_clk_3_S_in cby_1__2_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_3__6_ cbx_3__6_/SC_OUT_BOT cbx_3__5_/SC_IN_TOP grid_clb_3__6_/SC_OUT_TOP
+ cby_3__6_/Test_en_W_out grid_clb_3__6_/Test_en_E_out cby_3__6_/Test_en_W_out cby_2__6_/Test_en_W_in
+ VGND VPWR cbx_3__5_/REGIN_FEEDTHROUGH grid_clb_3__6_/bottom_width_0_height_0__pin_51_
+ cby_2__6_/ccff_tail cby_3__6_/ccff_head cbx_3__5_/clk_1_N_out cbx_3__5_/clk_1_N_out
+ cby_3__6_/prog_clk_0_W_in cbx_3__5_/prog_clk_1_N_out grid_clb_3__6_/prog_clk_0_N_out
+ cbx_3__5_/prog_clk_1_N_out cbx_3__5_/prog_clk_0_N_in grid_clb_3__6_/prog_clk_0_W_out
+ cby_3__6_/left_grid_pin_16_ cby_3__6_/left_grid_pin_17_ cby_3__6_/left_grid_pin_18_
+ cby_3__6_/left_grid_pin_19_ cby_3__6_/left_grid_pin_20_ cby_3__6_/left_grid_pin_21_
+ cby_3__6_/left_grid_pin_22_ cby_3__6_/left_grid_pin_23_ cby_3__6_/left_grid_pin_24_
+ cby_3__6_/left_grid_pin_25_ cby_3__6_/left_grid_pin_26_ cby_3__6_/left_grid_pin_27_
+ cby_3__6_/left_grid_pin_28_ cby_3__6_/left_grid_pin_29_ cby_3__6_/left_grid_pin_30_
+ cby_3__6_/left_grid_pin_31_ sb_3__5_/top_left_grid_pin_42_ sb_3__6_/bottom_left_grid_pin_42_
+ sb_3__5_/top_left_grid_pin_43_ sb_3__6_/bottom_left_grid_pin_43_ sb_3__5_/top_left_grid_pin_44_
+ sb_3__6_/bottom_left_grid_pin_44_ sb_3__5_/top_left_grid_pin_45_ sb_3__6_/bottom_left_grid_pin_45_
+ sb_3__5_/top_left_grid_pin_46_ sb_3__6_/bottom_left_grid_pin_46_ sb_3__5_/top_left_grid_pin_47_
+ sb_3__6_/bottom_left_grid_pin_47_ sb_3__5_/top_left_grid_pin_48_ sb_3__6_/bottom_left_grid_pin_48_
+ sb_3__5_/top_left_grid_pin_49_ sb_3__6_/bottom_left_grid_pin_49_ cbx_3__6_/bottom_grid_pin_0_
+ cbx_3__6_/bottom_grid_pin_10_ cbx_3__6_/bottom_grid_pin_11_ cbx_3__6_/bottom_grid_pin_12_
+ cbx_3__6_/bottom_grid_pin_13_ cbx_3__6_/bottom_grid_pin_14_ cbx_3__6_/bottom_grid_pin_15_
+ cbx_3__6_/bottom_grid_pin_1_ cbx_3__6_/bottom_grid_pin_2_ cbx_3__6_/REGOUT_FEEDTHROUGH
+ grid_clb_3__6_/top_width_0_height_0__pin_33_ sb_3__6_/left_bottom_grid_pin_34_ sb_2__6_/right_bottom_grid_pin_34_
+ sb_3__6_/left_bottom_grid_pin_35_ sb_2__6_/right_bottom_grid_pin_35_ sb_3__6_/left_bottom_grid_pin_36_
+ sb_2__6_/right_bottom_grid_pin_36_ sb_3__6_/left_bottom_grid_pin_37_ sb_2__6_/right_bottom_grid_pin_37_
+ sb_3__6_/left_bottom_grid_pin_38_ sb_2__6_/right_bottom_grid_pin_38_ sb_3__6_/left_bottom_grid_pin_39_
+ sb_2__6_/right_bottom_grid_pin_39_ cbx_3__6_/bottom_grid_pin_3_ sb_3__6_/left_bottom_grid_pin_40_
+ sb_2__6_/right_bottom_grid_pin_40_ sb_3__6_/left_bottom_grid_pin_41_ sb_2__6_/right_bottom_grid_pin_41_
+ cbx_3__6_/bottom_grid_pin_4_ cbx_3__6_/bottom_grid_pin_5_ cbx_3__6_/bottom_grid_pin_6_
+ cbx_3__6_/bottom_grid_pin_7_ cbx_3__6_/bottom_grid_pin_8_ cbx_3__6_/bottom_grid_pin_9_
+ grid_clb
Xcbx_1__3_ cbx_1__3_/REGIN_FEEDTHROUGH cbx_1__3_/REGOUT_FEEDTHROUGH cbx_1__3_/SC_IN_BOT
+ cbx_1__3_/SC_IN_TOP cbx_1__3_/SC_OUT_BOT cbx_1__3_/SC_OUT_TOP VGND VPWR cbx_1__3_/bottom_grid_pin_0_
+ cbx_1__3_/bottom_grid_pin_10_ cbx_1__3_/bottom_grid_pin_11_ cbx_1__3_/bottom_grid_pin_12_
+ cbx_1__3_/bottom_grid_pin_13_ cbx_1__3_/bottom_grid_pin_14_ cbx_1__3_/bottom_grid_pin_15_
+ cbx_1__3_/bottom_grid_pin_1_ cbx_1__3_/bottom_grid_pin_2_ cbx_1__3_/bottom_grid_pin_3_
+ cbx_1__3_/bottom_grid_pin_4_ cbx_1__3_/bottom_grid_pin_5_ cbx_1__3_/bottom_grid_pin_6_
+ cbx_1__3_/bottom_grid_pin_7_ cbx_1__3_/bottom_grid_pin_8_ cbx_1__3_/bottom_grid_pin_9_
+ sb_1__3_/ccff_tail sb_0__3_/ccff_head cbx_1__3_/chanx_left_in[0] cbx_1__3_/chanx_left_in[10]
+ cbx_1__3_/chanx_left_in[11] cbx_1__3_/chanx_left_in[12] cbx_1__3_/chanx_left_in[13]
+ cbx_1__3_/chanx_left_in[14] cbx_1__3_/chanx_left_in[15] cbx_1__3_/chanx_left_in[16]
+ cbx_1__3_/chanx_left_in[17] cbx_1__3_/chanx_left_in[18] cbx_1__3_/chanx_left_in[19]
+ cbx_1__3_/chanx_left_in[1] cbx_1__3_/chanx_left_in[2] cbx_1__3_/chanx_left_in[3]
+ cbx_1__3_/chanx_left_in[4] cbx_1__3_/chanx_left_in[5] cbx_1__3_/chanx_left_in[6]
+ cbx_1__3_/chanx_left_in[7] cbx_1__3_/chanx_left_in[8] cbx_1__3_/chanx_left_in[9]
+ sb_0__3_/chanx_right_in[0] sb_0__3_/chanx_right_in[10] sb_0__3_/chanx_right_in[11]
+ sb_0__3_/chanx_right_in[12] sb_0__3_/chanx_right_in[13] sb_0__3_/chanx_right_in[14]
+ sb_0__3_/chanx_right_in[15] sb_0__3_/chanx_right_in[16] sb_0__3_/chanx_right_in[17]
+ sb_0__3_/chanx_right_in[18] sb_0__3_/chanx_right_in[19] sb_0__3_/chanx_right_in[1]
+ sb_0__3_/chanx_right_in[2] sb_0__3_/chanx_right_in[3] sb_0__3_/chanx_right_in[4]
+ sb_0__3_/chanx_right_in[5] sb_0__3_/chanx_right_in[6] sb_0__3_/chanx_right_in[7]
+ sb_0__3_/chanx_right_in[8] sb_0__3_/chanx_right_in[9] sb_1__3_/chanx_left_out[0]
+ sb_1__3_/chanx_left_out[10] sb_1__3_/chanx_left_out[11] sb_1__3_/chanx_left_out[12]
+ sb_1__3_/chanx_left_out[13] sb_1__3_/chanx_left_out[14] sb_1__3_/chanx_left_out[15]
+ sb_1__3_/chanx_left_out[16] sb_1__3_/chanx_left_out[17] sb_1__3_/chanx_left_out[18]
+ sb_1__3_/chanx_left_out[19] sb_1__3_/chanx_left_out[1] sb_1__3_/chanx_left_out[2]
+ sb_1__3_/chanx_left_out[3] sb_1__3_/chanx_left_out[4] sb_1__3_/chanx_left_out[5]
+ sb_1__3_/chanx_left_out[6] sb_1__3_/chanx_left_out[7] sb_1__3_/chanx_left_out[8]
+ sb_1__3_/chanx_left_out[9] sb_1__3_/chanx_left_in[0] sb_1__3_/chanx_left_in[10]
+ sb_1__3_/chanx_left_in[11] sb_1__3_/chanx_left_in[12] sb_1__3_/chanx_left_in[13]
+ sb_1__3_/chanx_left_in[14] sb_1__3_/chanx_left_in[15] sb_1__3_/chanx_left_in[16]
+ sb_1__3_/chanx_left_in[17] sb_1__3_/chanx_left_in[18] sb_1__3_/chanx_left_in[19]
+ sb_1__3_/chanx_left_in[1] sb_1__3_/chanx_left_in[2] sb_1__3_/chanx_left_in[3] sb_1__3_/chanx_left_in[4]
+ sb_1__3_/chanx_left_in[5] sb_1__3_/chanx_left_in[6] sb_1__3_/chanx_left_in[7] sb_1__3_/chanx_left_in[8]
+ sb_1__3_/chanx_left_in[9] cbx_1__3_/clk_1_N_out cbx_1__3_/clk_1_S_out sb_1__3_/clk_1_W_out
+ cbx_1__3_/clk_2_E_out cbx_1__3_/clk_2_W_in cbx_1__3_/clk_2_W_out cbx_1__3_/clk_3_E_out
+ cbx_1__3_/clk_3_W_in cbx_1__3_/clk_3_W_out cbx_1__3_/prog_clk_0_N_in sb_0__3_/prog_clk_0_E_in
+ cbx_1__3_/prog_clk_1_N_out cbx_1__3_/prog_clk_1_S_out sb_1__3_/prog_clk_1_W_out
+ cbx_1__3_/prog_clk_2_E_out cbx_1__3_/prog_clk_2_W_in cbx_1__3_/prog_clk_2_W_out
+ cbx_1__3_/prog_clk_3_E_out cbx_1__3_/prog_clk_3_W_in cbx_1__3_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_5__0_ sb_5__0_/SC_IN_TOP sb_5__0_/SC_OUT_TOP sb_5__0_/Test_en_N_out sb_5__0_/Test_en_S_in
+ VGND VPWR sb_5__0_/ccff_head sb_5__0_/ccff_tail sb_5__0_/chanx_left_in[0] sb_5__0_/chanx_left_in[10]
+ sb_5__0_/chanx_left_in[11] sb_5__0_/chanx_left_in[12] sb_5__0_/chanx_left_in[13]
+ sb_5__0_/chanx_left_in[14] sb_5__0_/chanx_left_in[15] sb_5__0_/chanx_left_in[16]
+ sb_5__0_/chanx_left_in[17] sb_5__0_/chanx_left_in[18] sb_5__0_/chanx_left_in[19]
+ sb_5__0_/chanx_left_in[1] sb_5__0_/chanx_left_in[2] sb_5__0_/chanx_left_in[3] sb_5__0_/chanx_left_in[4]
+ sb_5__0_/chanx_left_in[5] sb_5__0_/chanx_left_in[6] sb_5__0_/chanx_left_in[7] sb_5__0_/chanx_left_in[8]
+ sb_5__0_/chanx_left_in[9] sb_5__0_/chanx_left_out[0] sb_5__0_/chanx_left_out[10]
+ sb_5__0_/chanx_left_out[11] sb_5__0_/chanx_left_out[12] sb_5__0_/chanx_left_out[13]
+ sb_5__0_/chanx_left_out[14] sb_5__0_/chanx_left_out[15] sb_5__0_/chanx_left_out[16]
+ sb_5__0_/chanx_left_out[17] sb_5__0_/chanx_left_out[18] sb_5__0_/chanx_left_out[19]
+ sb_5__0_/chanx_left_out[1] sb_5__0_/chanx_left_out[2] sb_5__0_/chanx_left_out[3]
+ sb_5__0_/chanx_left_out[4] sb_5__0_/chanx_left_out[5] sb_5__0_/chanx_left_out[6]
+ sb_5__0_/chanx_left_out[7] sb_5__0_/chanx_left_out[8] sb_5__0_/chanx_left_out[9]
+ sb_5__0_/chanx_right_in[0] sb_5__0_/chanx_right_in[10] sb_5__0_/chanx_right_in[11]
+ sb_5__0_/chanx_right_in[12] sb_5__0_/chanx_right_in[13] sb_5__0_/chanx_right_in[14]
+ sb_5__0_/chanx_right_in[15] sb_5__0_/chanx_right_in[16] sb_5__0_/chanx_right_in[17]
+ sb_5__0_/chanx_right_in[18] sb_5__0_/chanx_right_in[19] sb_5__0_/chanx_right_in[1]
+ sb_5__0_/chanx_right_in[2] sb_5__0_/chanx_right_in[3] sb_5__0_/chanx_right_in[4]
+ sb_5__0_/chanx_right_in[5] sb_5__0_/chanx_right_in[6] sb_5__0_/chanx_right_in[7]
+ sb_5__0_/chanx_right_in[8] sb_5__0_/chanx_right_in[9] cbx_6__0_/chanx_left_in[0]
+ cbx_6__0_/chanx_left_in[10] cbx_6__0_/chanx_left_in[11] cbx_6__0_/chanx_left_in[12]
+ cbx_6__0_/chanx_left_in[13] cbx_6__0_/chanx_left_in[14] cbx_6__0_/chanx_left_in[15]
+ cbx_6__0_/chanx_left_in[16] cbx_6__0_/chanx_left_in[17] cbx_6__0_/chanx_left_in[18]
+ cbx_6__0_/chanx_left_in[19] cbx_6__0_/chanx_left_in[1] cbx_6__0_/chanx_left_in[2]
+ cbx_6__0_/chanx_left_in[3] cbx_6__0_/chanx_left_in[4] cbx_6__0_/chanx_left_in[5]
+ cbx_6__0_/chanx_left_in[6] cbx_6__0_/chanx_left_in[7] cbx_6__0_/chanx_left_in[8]
+ cbx_6__0_/chanx_left_in[9] sb_5__0_/chany_top_in[0] sb_5__0_/chany_top_in[10] sb_5__0_/chany_top_in[11]
+ sb_5__0_/chany_top_in[12] sb_5__0_/chany_top_in[13] sb_5__0_/chany_top_in[14] sb_5__0_/chany_top_in[15]
+ sb_5__0_/chany_top_in[16] sb_5__0_/chany_top_in[17] sb_5__0_/chany_top_in[18] sb_5__0_/chany_top_in[19]
+ sb_5__0_/chany_top_in[1] sb_5__0_/chany_top_in[2] sb_5__0_/chany_top_in[3] sb_5__0_/chany_top_in[4]
+ sb_5__0_/chany_top_in[5] sb_5__0_/chany_top_in[6] sb_5__0_/chany_top_in[7] sb_5__0_/chany_top_in[8]
+ sb_5__0_/chany_top_in[9] sb_5__0_/chany_top_out[0] sb_5__0_/chany_top_out[10] sb_5__0_/chany_top_out[11]
+ sb_5__0_/chany_top_out[12] sb_5__0_/chany_top_out[13] sb_5__0_/chany_top_out[14]
+ sb_5__0_/chany_top_out[15] sb_5__0_/chany_top_out[16] sb_5__0_/chany_top_out[17]
+ sb_5__0_/chany_top_out[18] sb_5__0_/chany_top_out[19] sb_5__0_/chany_top_out[1]
+ sb_5__0_/chany_top_out[2] sb_5__0_/chany_top_out[3] sb_5__0_/chany_top_out[4] sb_5__0_/chany_top_out[5]
+ sb_5__0_/chany_top_out[6] sb_5__0_/chany_top_out[7] sb_5__0_/chany_top_out[8] sb_5__0_/chany_top_out[9]
+ sb_5__0_/clk_3_N_out sb_5__0_/clk_3_S_in sb_5__0_/left_bottom_grid_pin_11_ sb_5__0_/left_bottom_grid_pin_13_
+ sb_5__0_/left_bottom_grid_pin_15_ sb_5__0_/left_bottom_grid_pin_17_ sb_5__0_/left_bottom_grid_pin_1_
+ sb_5__0_/left_bottom_grid_pin_3_ sb_5__0_/left_bottom_grid_pin_5_ sb_5__0_/left_bottom_grid_pin_7_
+ sb_5__0_/left_bottom_grid_pin_9_ sb_5__0_/prog_clk_0_N_in sb_5__0_/prog_clk_3_N_out
+ sb_5__0_/prog_clk_3_S_in sb_5__0_/right_bottom_grid_pin_11_ sb_5__0_/right_bottom_grid_pin_13_
+ sb_5__0_/right_bottom_grid_pin_15_ sb_5__0_/right_bottom_grid_pin_17_ sb_5__0_/right_bottom_grid_pin_1_
+ sb_5__0_/right_bottom_grid_pin_3_ sb_5__0_/right_bottom_grid_pin_5_ sb_5__0_/right_bottom_grid_pin_7_
+ sb_5__0_/right_bottom_grid_pin_9_ sb_5__0_/top_left_grid_pin_42_ sb_5__0_/top_left_grid_pin_43_
+ sb_5__0_/top_left_grid_pin_44_ sb_5__0_/top_left_grid_pin_45_ sb_5__0_/top_left_grid_pin_46_
+ sb_5__0_/top_left_grid_pin_47_ sb_5__0_/top_left_grid_pin_48_ sb_5__0_/top_left_grid_pin_49_
+ sb_1__0_
Xsb_1__8_ sb_1__8_/SC_IN_BOT sb_1__8_/SC_OUT_BOT VGND VPWR sb_1__8_/bottom_left_grid_pin_42_
+ sb_1__8_/bottom_left_grid_pin_43_ sb_1__8_/bottom_left_grid_pin_44_ sb_1__8_/bottom_left_grid_pin_45_
+ sb_1__8_/bottom_left_grid_pin_46_ sb_1__8_/bottom_left_grid_pin_47_ sb_1__8_/bottom_left_grid_pin_48_
+ sb_1__8_/bottom_left_grid_pin_49_ sb_1__8_/ccff_head sb_1__8_/ccff_tail sb_1__8_/chanx_left_in[0]
+ sb_1__8_/chanx_left_in[10] sb_1__8_/chanx_left_in[11] sb_1__8_/chanx_left_in[12]
+ sb_1__8_/chanx_left_in[13] sb_1__8_/chanx_left_in[14] sb_1__8_/chanx_left_in[15]
+ sb_1__8_/chanx_left_in[16] sb_1__8_/chanx_left_in[17] sb_1__8_/chanx_left_in[18]
+ sb_1__8_/chanx_left_in[19] sb_1__8_/chanx_left_in[1] sb_1__8_/chanx_left_in[2] sb_1__8_/chanx_left_in[3]
+ sb_1__8_/chanx_left_in[4] sb_1__8_/chanx_left_in[5] sb_1__8_/chanx_left_in[6] sb_1__8_/chanx_left_in[7]
+ sb_1__8_/chanx_left_in[8] sb_1__8_/chanx_left_in[9] sb_1__8_/chanx_left_out[0] sb_1__8_/chanx_left_out[10]
+ sb_1__8_/chanx_left_out[11] sb_1__8_/chanx_left_out[12] sb_1__8_/chanx_left_out[13]
+ sb_1__8_/chanx_left_out[14] sb_1__8_/chanx_left_out[15] sb_1__8_/chanx_left_out[16]
+ sb_1__8_/chanx_left_out[17] sb_1__8_/chanx_left_out[18] sb_1__8_/chanx_left_out[19]
+ sb_1__8_/chanx_left_out[1] sb_1__8_/chanx_left_out[2] sb_1__8_/chanx_left_out[3]
+ sb_1__8_/chanx_left_out[4] sb_1__8_/chanx_left_out[5] sb_1__8_/chanx_left_out[6]
+ sb_1__8_/chanx_left_out[7] sb_1__8_/chanx_left_out[8] sb_1__8_/chanx_left_out[9]
+ sb_1__8_/chanx_right_in[0] sb_1__8_/chanx_right_in[10] sb_1__8_/chanx_right_in[11]
+ sb_1__8_/chanx_right_in[12] sb_1__8_/chanx_right_in[13] sb_1__8_/chanx_right_in[14]
+ sb_1__8_/chanx_right_in[15] sb_1__8_/chanx_right_in[16] sb_1__8_/chanx_right_in[17]
+ sb_1__8_/chanx_right_in[18] sb_1__8_/chanx_right_in[19] sb_1__8_/chanx_right_in[1]
+ sb_1__8_/chanx_right_in[2] sb_1__8_/chanx_right_in[3] sb_1__8_/chanx_right_in[4]
+ sb_1__8_/chanx_right_in[5] sb_1__8_/chanx_right_in[6] sb_1__8_/chanx_right_in[7]
+ sb_1__8_/chanx_right_in[8] sb_1__8_/chanx_right_in[9] cbx_2__8_/chanx_left_in[0]
+ cbx_2__8_/chanx_left_in[10] cbx_2__8_/chanx_left_in[11] cbx_2__8_/chanx_left_in[12]
+ cbx_2__8_/chanx_left_in[13] cbx_2__8_/chanx_left_in[14] cbx_2__8_/chanx_left_in[15]
+ cbx_2__8_/chanx_left_in[16] cbx_2__8_/chanx_left_in[17] cbx_2__8_/chanx_left_in[18]
+ cbx_2__8_/chanx_left_in[19] cbx_2__8_/chanx_left_in[1] cbx_2__8_/chanx_left_in[2]
+ cbx_2__8_/chanx_left_in[3] cbx_2__8_/chanx_left_in[4] cbx_2__8_/chanx_left_in[5]
+ cbx_2__8_/chanx_left_in[6] cbx_2__8_/chanx_left_in[7] cbx_2__8_/chanx_left_in[8]
+ cbx_2__8_/chanx_left_in[9] cby_1__8_/chany_top_out[0] cby_1__8_/chany_top_out[10]
+ cby_1__8_/chany_top_out[11] cby_1__8_/chany_top_out[12] cby_1__8_/chany_top_out[13]
+ cby_1__8_/chany_top_out[14] cby_1__8_/chany_top_out[15] cby_1__8_/chany_top_out[16]
+ cby_1__8_/chany_top_out[17] cby_1__8_/chany_top_out[18] cby_1__8_/chany_top_out[19]
+ cby_1__8_/chany_top_out[1] cby_1__8_/chany_top_out[2] cby_1__8_/chany_top_out[3]
+ cby_1__8_/chany_top_out[4] cby_1__8_/chany_top_out[5] cby_1__8_/chany_top_out[6]
+ cby_1__8_/chany_top_out[7] cby_1__8_/chany_top_out[8] cby_1__8_/chany_top_out[9]
+ cby_1__8_/chany_top_in[0] cby_1__8_/chany_top_in[10] cby_1__8_/chany_top_in[11]
+ cby_1__8_/chany_top_in[12] cby_1__8_/chany_top_in[13] cby_1__8_/chany_top_in[14]
+ cby_1__8_/chany_top_in[15] cby_1__8_/chany_top_in[16] cby_1__8_/chany_top_in[17]
+ cby_1__8_/chany_top_in[18] cby_1__8_/chany_top_in[19] cby_1__8_/chany_top_in[1]
+ cby_1__8_/chany_top_in[2] cby_1__8_/chany_top_in[3] cby_1__8_/chany_top_in[4] cby_1__8_/chany_top_in[5]
+ cby_1__8_/chany_top_in[6] cby_1__8_/chany_top_in[7] cby_1__8_/chany_top_in[8] cby_1__8_/chany_top_in[9]
+ sb_1__8_/left_bottom_grid_pin_34_ sb_1__8_/left_bottom_grid_pin_35_ sb_1__8_/left_bottom_grid_pin_36_
+ sb_1__8_/left_bottom_grid_pin_37_ sb_1__8_/left_bottom_grid_pin_38_ sb_1__8_/left_bottom_grid_pin_39_
+ sb_1__8_/left_bottom_grid_pin_40_ sb_1__8_/left_bottom_grid_pin_41_ sb_1__8_/left_top_grid_pin_1_
+ sb_1__8_/prog_clk_0_S_in sb_1__8_/right_bottom_grid_pin_34_ sb_1__8_/right_bottom_grid_pin_35_
+ sb_1__8_/right_bottom_grid_pin_36_ sb_1__8_/right_bottom_grid_pin_37_ sb_1__8_/right_bottom_grid_pin_38_
+ sb_1__8_/right_bottom_grid_pin_39_ sb_1__8_/right_bottom_grid_pin_40_ sb_1__8_/right_bottom_grid_pin_41_
+ sb_1__8_/right_top_grid_pin_1_ sb_1__2_
Xcby_7__7_ cby_7__7_/Test_en_W_in cby_7__7_/Test_en_E_out cby_7__7_/Test_en_N_out
+ cby_7__7_/Test_en_W_in cby_7__7_/Test_en_W_in cby_7__7_/Test_en_W_out VGND VPWR
+ cby_7__7_/ccff_head cby_7__7_/ccff_tail sb_7__6_/chany_top_out[0] sb_7__6_/chany_top_out[10]
+ sb_7__6_/chany_top_out[11] sb_7__6_/chany_top_out[12] sb_7__6_/chany_top_out[13]
+ sb_7__6_/chany_top_out[14] sb_7__6_/chany_top_out[15] sb_7__6_/chany_top_out[16]
+ sb_7__6_/chany_top_out[17] sb_7__6_/chany_top_out[18] sb_7__6_/chany_top_out[19]
+ sb_7__6_/chany_top_out[1] sb_7__6_/chany_top_out[2] sb_7__6_/chany_top_out[3] sb_7__6_/chany_top_out[4]
+ sb_7__6_/chany_top_out[5] sb_7__6_/chany_top_out[6] sb_7__6_/chany_top_out[7] sb_7__6_/chany_top_out[8]
+ sb_7__6_/chany_top_out[9] sb_7__6_/chany_top_in[0] sb_7__6_/chany_top_in[10] sb_7__6_/chany_top_in[11]
+ sb_7__6_/chany_top_in[12] sb_7__6_/chany_top_in[13] sb_7__6_/chany_top_in[14] sb_7__6_/chany_top_in[15]
+ sb_7__6_/chany_top_in[16] sb_7__6_/chany_top_in[17] sb_7__6_/chany_top_in[18] sb_7__6_/chany_top_in[19]
+ sb_7__6_/chany_top_in[1] sb_7__6_/chany_top_in[2] sb_7__6_/chany_top_in[3] sb_7__6_/chany_top_in[4]
+ sb_7__6_/chany_top_in[5] sb_7__6_/chany_top_in[6] sb_7__6_/chany_top_in[7] sb_7__6_/chany_top_in[8]
+ sb_7__6_/chany_top_in[9] cby_7__7_/chany_top_in[0] cby_7__7_/chany_top_in[10] cby_7__7_/chany_top_in[11]
+ cby_7__7_/chany_top_in[12] cby_7__7_/chany_top_in[13] cby_7__7_/chany_top_in[14]
+ cby_7__7_/chany_top_in[15] cby_7__7_/chany_top_in[16] cby_7__7_/chany_top_in[17]
+ cby_7__7_/chany_top_in[18] cby_7__7_/chany_top_in[19] cby_7__7_/chany_top_in[1]
+ cby_7__7_/chany_top_in[2] cby_7__7_/chany_top_in[3] cby_7__7_/chany_top_in[4] cby_7__7_/chany_top_in[5]
+ cby_7__7_/chany_top_in[6] cby_7__7_/chany_top_in[7] cby_7__7_/chany_top_in[8] cby_7__7_/chany_top_in[9]
+ cby_7__7_/chany_top_out[0] cby_7__7_/chany_top_out[10] cby_7__7_/chany_top_out[11]
+ cby_7__7_/chany_top_out[12] cby_7__7_/chany_top_out[13] cby_7__7_/chany_top_out[14]
+ cby_7__7_/chany_top_out[15] cby_7__7_/chany_top_out[16] cby_7__7_/chany_top_out[17]
+ cby_7__7_/chany_top_out[18] cby_7__7_/chany_top_out[19] cby_7__7_/chany_top_out[1]
+ cby_7__7_/chany_top_out[2] cby_7__7_/chany_top_out[3] cby_7__7_/chany_top_out[4]
+ cby_7__7_/chany_top_out[5] cby_7__7_/chany_top_out[6] cby_7__7_/chany_top_out[7]
+ cby_7__7_/chany_top_out[8] cby_7__7_/chany_top_out[9] sb_7__7_/clk_1_N_in sb_7__6_/clk_2_N_out
+ cby_7__7_/clk_2_S_out cby_7__7_/clk_3_N_out cby_7__7_/clk_3_S_in cby_7__7_/clk_3_S_out
+ cby_7__7_/left_grid_pin_16_ cby_7__7_/left_grid_pin_17_ cby_7__7_/left_grid_pin_18_
+ cby_7__7_/left_grid_pin_19_ cby_7__7_/left_grid_pin_20_ cby_7__7_/left_grid_pin_21_
+ cby_7__7_/left_grid_pin_22_ cby_7__7_/left_grid_pin_23_ cby_7__7_/left_grid_pin_24_
+ cby_7__7_/left_grid_pin_25_ cby_7__7_/left_grid_pin_26_ cby_7__7_/left_grid_pin_27_
+ cby_7__7_/left_grid_pin_28_ cby_7__7_/left_grid_pin_29_ cby_7__7_/left_grid_pin_30_
+ cby_7__7_/left_grid_pin_31_ cby_7__7_/prog_clk_0_N_out sb_7__6_/prog_clk_0_N_in
+ cby_7__7_/prog_clk_0_W_in sb_7__7_/prog_clk_1_N_in sb_7__6_/prog_clk_2_N_out cby_7__7_/prog_clk_2_S_out
+ cby_7__7_/prog_clk_3_N_out cby_7__7_/prog_clk_3_S_in cby_7__7_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_7__8_ IO_ISOL_N cbx_7__8_/SC_IN_BOT sb_6__8_/SC_OUT_BOT cbx_7__8_/SC_OUT_BOT
+ cbx_7__8_/SC_OUT_TOP VGND VPWR cbx_7__8_/bottom_grid_pin_0_ cbx_7__8_/bottom_grid_pin_10_
+ cbx_7__8_/bottom_grid_pin_11_ cbx_7__8_/bottom_grid_pin_12_ cbx_7__8_/bottom_grid_pin_13_
+ cbx_7__8_/bottom_grid_pin_14_ cbx_7__8_/bottom_grid_pin_15_ cbx_7__8_/bottom_grid_pin_1_
+ cbx_7__8_/bottom_grid_pin_2_ cbx_7__8_/bottom_grid_pin_3_ cbx_7__8_/bottom_grid_pin_4_
+ cbx_7__8_/bottom_grid_pin_5_ cbx_7__8_/bottom_grid_pin_6_ cbx_7__8_/bottom_grid_pin_7_
+ cbx_7__8_/bottom_grid_pin_8_ cbx_7__8_/bottom_grid_pin_9_ cbx_7__8_/top_grid_pin_0_
+ sb_7__8_/left_top_grid_pin_1_ sb_6__8_/right_top_grid_pin_1_ sb_7__8_/ccff_tail
+ sb_6__8_/ccff_head cbx_7__8_/chanx_left_in[0] cbx_7__8_/chanx_left_in[10] cbx_7__8_/chanx_left_in[11]
+ cbx_7__8_/chanx_left_in[12] cbx_7__8_/chanx_left_in[13] cbx_7__8_/chanx_left_in[14]
+ cbx_7__8_/chanx_left_in[15] cbx_7__8_/chanx_left_in[16] cbx_7__8_/chanx_left_in[17]
+ cbx_7__8_/chanx_left_in[18] cbx_7__8_/chanx_left_in[19] cbx_7__8_/chanx_left_in[1]
+ cbx_7__8_/chanx_left_in[2] cbx_7__8_/chanx_left_in[3] cbx_7__8_/chanx_left_in[4]
+ cbx_7__8_/chanx_left_in[5] cbx_7__8_/chanx_left_in[6] cbx_7__8_/chanx_left_in[7]
+ cbx_7__8_/chanx_left_in[8] cbx_7__8_/chanx_left_in[9] sb_6__8_/chanx_right_in[0]
+ sb_6__8_/chanx_right_in[10] sb_6__8_/chanx_right_in[11] sb_6__8_/chanx_right_in[12]
+ sb_6__8_/chanx_right_in[13] sb_6__8_/chanx_right_in[14] sb_6__8_/chanx_right_in[15]
+ sb_6__8_/chanx_right_in[16] sb_6__8_/chanx_right_in[17] sb_6__8_/chanx_right_in[18]
+ sb_6__8_/chanx_right_in[19] sb_6__8_/chanx_right_in[1] sb_6__8_/chanx_right_in[2]
+ sb_6__8_/chanx_right_in[3] sb_6__8_/chanx_right_in[4] sb_6__8_/chanx_right_in[5]
+ sb_6__8_/chanx_right_in[6] sb_6__8_/chanx_right_in[7] sb_6__8_/chanx_right_in[8]
+ sb_6__8_/chanx_right_in[9] sb_7__8_/chanx_left_out[0] sb_7__8_/chanx_left_out[10]
+ sb_7__8_/chanx_left_out[11] sb_7__8_/chanx_left_out[12] sb_7__8_/chanx_left_out[13]
+ sb_7__8_/chanx_left_out[14] sb_7__8_/chanx_left_out[15] sb_7__8_/chanx_left_out[16]
+ sb_7__8_/chanx_left_out[17] sb_7__8_/chanx_left_out[18] sb_7__8_/chanx_left_out[19]
+ sb_7__8_/chanx_left_out[1] sb_7__8_/chanx_left_out[2] sb_7__8_/chanx_left_out[3]
+ sb_7__8_/chanx_left_out[4] sb_7__8_/chanx_left_out[5] sb_7__8_/chanx_left_out[6]
+ sb_7__8_/chanx_left_out[7] sb_7__8_/chanx_left_out[8] sb_7__8_/chanx_left_out[9]
+ sb_7__8_/chanx_left_in[0] sb_7__8_/chanx_left_in[10] sb_7__8_/chanx_left_in[11]
+ sb_7__8_/chanx_left_in[12] sb_7__8_/chanx_left_in[13] sb_7__8_/chanx_left_in[14]
+ sb_7__8_/chanx_left_in[15] sb_7__8_/chanx_left_in[16] sb_7__8_/chanx_left_in[17]
+ sb_7__8_/chanx_left_in[18] sb_7__8_/chanx_left_in[19] sb_7__8_/chanx_left_in[1]
+ sb_7__8_/chanx_left_in[2] sb_7__8_/chanx_left_in[3] sb_7__8_/chanx_left_in[4] sb_7__8_/chanx_left_in[5]
+ sb_7__8_/chanx_left_in[6] sb_7__8_/chanx_left_in[7] sb_7__8_/chanx_left_in[8] sb_7__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
+ cbx_7__8_/prog_clk_0_S_in cbx_7__8_/prog_clk_0_W_out cbx_7__8_/top_grid_pin_0_ cbx_1__2_
Xcby_4__4_ sb_4__3_/Test_en_N_out cby_4__4_/Test_en_E_out sb_4__4_/Test_en_S_in sb_4__3_/Test_en_N_out
+ sb_4__3_/Test_en_N_out cby_4__4_/Test_en_W_out VGND VPWR cby_4__4_/ccff_head cby_4__4_/ccff_tail
+ sb_4__3_/chany_top_out[0] sb_4__3_/chany_top_out[10] sb_4__3_/chany_top_out[11]
+ sb_4__3_/chany_top_out[12] sb_4__3_/chany_top_out[13] sb_4__3_/chany_top_out[14]
+ sb_4__3_/chany_top_out[15] sb_4__3_/chany_top_out[16] sb_4__3_/chany_top_out[17]
+ sb_4__3_/chany_top_out[18] sb_4__3_/chany_top_out[19] sb_4__3_/chany_top_out[1]
+ sb_4__3_/chany_top_out[2] sb_4__3_/chany_top_out[3] sb_4__3_/chany_top_out[4] sb_4__3_/chany_top_out[5]
+ sb_4__3_/chany_top_out[6] sb_4__3_/chany_top_out[7] sb_4__3_/chany_top_out[8] sb_4__3_/chany_top_out[9]
+ sb_4__3_/chany_top_in[0] sb_4__3_/chany_top_in[10] sb_4__3_/chany_top_in[11] sb_4__3_/chany_top_in[12]
+ sb_4__3_/chany_top_in[13] sb_4__3_/chany_top_in[14] sb_4__3_/chany_top_in[15] sb_4__3_/chany_top_in[16]
+ sb_4__3_/chany_top_in[17] sb_4__3_/chany_top_in[18] sb_4__3_/chany_top_in[19] sb_4__3_/chany_top_in[1]
+ sb_4__3_/chany_top_in[2] sb_4__3_/chany_top_in[3] sb_4__3_/chany_top_in[4] sb_4__3_/chany_top_in[5]
+ sb_4__3_/chany_top_in[6] sb_4__3_/chany_top_in[7] sb_4__3_/chany_top_in[8] sb_4__3_/chany_top_in[9]
+ cby_4__4_/chany_top_in[0] cby_4__4_/chany_top_in[10] cby_4__4_/chany_top_in[11]
+ cby_4__4_/chany_top_in[12] cby_4__4_/chany_top_in[13] cby_4__4_/chany_top_in[14]
+ cby_4__4_/chany_top_in[15] cby_4__4_/chany_top_in[16] cby_4__4_/chany_top_in[17]
+ cby_4__4_/chany_top_in[18] cby_4__4_/chany_top_in[19] cby_4__4_/chany_top_in[1]
+ cby_4__4_/chany_top_in[2] cby_4__4_/chany_top_in[3] cby_4__4_/chany_top_in[4] cby_4__4_/chany_top_in[5]
+ cby_4__4_/chany_top_in[6] cby_4__4_/chany_top_in[7] cby_4__4_/chany_top_in[8] cby_4__4_/chany_top_in[9]
+ cby_4__4_/chany_top_out[0] cby_4__4_/chany_top_out[10] cby_4__4_/chany_top_out[11]
+ cby_4__4_/chany_top_out[12] cby_4__4_/chany_top_out[13] cby_4__4_/chany_top_out[14]
+ cby_4__4_/chany_top_out[15] cby_4__4_/chany_top_out[16] cby_4__4_/chany_top_out[17]
+ cby_4__4_/chany_top_out[18] cby_4__4_/chany_top_out[19] cby_4__4_/chany_top_out[1]
+ cby_4__4_/chany_top_out[2] cby_4__4_/chany_top_out[3] cby_4__4_/chany_top_out[4]
+ cby_4__4_/chany_top_out[5] cby_4__4_/chany_top_out[6] cby_4__4_/chany_top_out[7]
+ cby_4__4_/chany_top_out[8] cby_4__4_/chany_top_out[9] cby_4__4_/clk_2_N_out cby_4__4_/clk_2_S_in
+ cby_4__4_/clk_2_S_out sb_4__4_/clk_3_N_in sb_4__3_/clk_3_N_out cby_4__4_/clk_3_S_out
+ cby_4__4_/left_grid_pin_16_ cby_4__4_/left_grid_pin_17_ cby_4__4_/left_grid_pin_18_
+ cby_4__4_/left_grid_pin_19_ cby_4__4_/left_grid_pin_20_ cby_4__4_/left_grid_pin_21_
+ cby_4__4_/left_grid_pin_22_ cby_4__4_/left_grid_pin_23_ cby_4__4_/left_grid_pin_24_
+ cby_4__4_/left_grid_pin_25_ cby_4__4_/left_grid_pin_26_ cby_4__4_/left_grid_pin_27_
+ cby_4__4_/left_grid_pin_28_ cby_4__4_/left_grid_pin_29_ cby_4__4_/left_grid_pin_30_
+ cby_4__4_/left_grid_pin_31_ cby_4__4_/prog_clk_0_N_out sb_4__3_/prog_clk_0_N_in
+ cby_4__4_/prog_clk_0_W_in cby_4__4_/prog_clk_2_N_out cby_4__4_/prog_clk_2_S_in cby_4__4_/prog_clk_2_S_out
+ sb_4__4_/prog_clk_3_N_in sb_4__3_/prog_clk_3_N_out cby_4__4_/prog_clk_3_S_out cby_1__1_
Xcby_1__1_ cby_1__1_/Test_en_W_in cby_1__1_/Test_en_E_out cby_1__1_/Test_en_N_out
+ cby_1__1_/Test_en_W_in cby_1__1_/Test_en_W_in cby_1__1_/Test_en_W_out VGND VPWR
+ cby_1__1_/ccff_head cby_1__1_/ccff_tail sb_1__0_/chany_top_out[0] sb_1__0_/chany_top_out[10]
+ sb_1__0_/chany_top_out[11] sb_1__0_/chany_top_out[12] sb_1__0_/chany_top_out[13]
+ sb_1__0_/chany_top_out[14] sb_1__0_/chany_top_out[15] sb_1__0_/chany_top_out[16]
+ sb_1__0_/chany_top_out[17] sb_1__0_/chany_top_out[18] sb_1__0_/chany_top_out[19]
+ sb_1__0_/chany_top_out[1] sb_1__0_/chany_top_out[2] sb_1__0_/chany_top_out[3] sb_1__0_/chany_top_out[4]
+ sb_1__0_/chany_top_out[5] sb_1__0_/chany_top_out[6] sb_1__0_/chany_top_out[7] sb_1__0_/chany_top_out[8]
+ sb_1__0_/chany_top_out[9] sb_1__0_/chany_top_in[0] sb_1__0_/chany_top_in[10] sb_1__0_/chany_top_in[11]
+ sb_1__0_/chany_top_in[12] sb_1__0_/chany_top_in[13] sb_1__0_/chany_top_in[14] sb_1__0_/chany_top_in[15]
+ sb_1__0_/chany_top_in[16] sb_1__0_/chany_top_in[17] sb_1__0_/chany_top_in[18] sb_1__0_/chany_top_in[19]
+ sb_1__0_/chany_top_in[1] sb_1__0_/chany_top_in[2] sb_1__0_/chany_top_in[3] sb_1__0_/chany_top_in[4]
+ sb_1__0_/chany_top_in[5] sb_1__0_/chany_top_in[6] sb_1__0_/chany_top_in[7] sb_1__0_/chany_top_in[8]
+ sb_1__0_/chany_top_in[9] cby_1__1_/chany_top_in[0] cby_1__1_/chany_top_in[10] cby_1__1_/chany_top_in[11]
+ cby_1__1_/chany_top_in[12] cby_1__1_/chany_top_in[13] cby_1__1_/chany_top_in[14]
+ cby_1__1_/chany_top_in[15] cby_1__1_/chany_top_in[16] cby_1__1_/chany_top_in[17]
+ cby_1__1_/chany_top_in[18] cby_1__1_/chany_top_in[19] cby_1__1_/chany_top_in[1]
+ cby_1__1_/chany_top_in[2] cby_1__1_/chany_top_in[3] cby_1__1_/chany_top_in[4] cby_1__1_/chany_top_in[5]
+ cby_1__1_/chany_top_in[6] cby_1__1_/chany_top_in[7] cby_1__1_/chany_top_in[8] cby_1__1_/chany_top_in[9]
+ cby_1__1_/chany_top_out[0] cby_1__1_/chany_top_out[10] cby_1__1_/chany_top_out[11]
+ cby_1__1_/chany_top_out[12] cby_1__1_/chany_top_out[13] cby_1__1_/chany_top_out[14]
+ cby_1__1_/chany_top_out[15] cby_1__1_/chany_top_out[16] cby_1__1_/chany_top_out[17]
+ cby_1__1_/chany_top_out[18] cby_1__1_/chany_top_out[19] cby_1__1_/chany_top_out[1]
+ cby_1__1_/chany_top_out[2] cby_1__1_/chany_top_out[3] cby_1__1_/chany_top_out[4]
+ cby_1__1_/chany_top_out[5] cby_1__1_/chany_top_out[6] cby_1__1_/chany_top_out[7]
+ cby_1__1_/chany_top_out[8] cby_1__1_/chany_top_out[9] cby_1__1_/clk_2_N_out cby_1__1_/clk_2_S_in
+ cby_1__1_/clk_2_S_out cby_1__1_/clk_3_N_out cby_1__1_/clk_3_S_in cby_1__1_/clk_3_S_out
+ cby_1__1_/left_grid_pin_16_ cby_1__1_/left_grid_pin_17_ cby_1__1_/left_grid_pin_18_
+ cby_1__1_/left_grid_pin_19_ cby_1__1_/left_grid_pin_20_ cby_1__1_/left_grid_pin_21_
+ cby_1__1_/left_grid_pin_22_ cby_1__1_/left_grid_pin_23_ cby_1__1_/left_grid_pin_24_
+ cby_1__1_/left_grid_pin_25_ cby_1__1_/left_grid_pin_26_ cby_1__1_/left_grid_pin_27_
+ cby_1__1_/left_grid_pin_28_ cby_1__1_/left_grid_pin_29_ cby_1__1_/left_grid_pin_30_
+ cby_1__1_/left_grid_pin_31_ cby_1__1_/prog_clk_0_N_out sb_1__0_/prog_clk_0_N_in
+ cby_1__1_/prog_clk_0_W_in cby_1__1_/prog_clk_2_N_out cby_1__1_/prog_clk_2_S_in cby_1__1_/prog_clk_2_S_out
+ cby_1__1_/prog_clk_3_N_out cby_1__1_/prog_clk_3_S_in cby_1__1_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_6__8_ cbx_6__7_/SC_OUT_TOP grid_clb_6__8_/SC_OUT_BOT cbx_6__8_/SC_IN_BOT
+ cby_5__8_/Test_en_E_out cby_6__8_/Test_en_W_in cby_5__8_/Test_en_E_out grid_clb_6__8_/Test_en_W_out
+ VGND VPWR cbx_6__7_/REGIN_FEEDTHROUGH grid_clb_6__8_/bottom_width_0_height_0__pin_51_
+ cby_5__8_/ccff_tail cby_6__8_/ccff_head cbx_6__7_/clk_1_N_out cbx_6__7_/clk_1_N_out
+ cby_6__8_/prog_clk_0_W_in cbx_6__7_/prog_clk_1_N_out cbx_6__8_/prog_clk_0_S_in cbx_6__7_/prog_clk_1_N_out
+ cbx_6__7_/prog_clk_0_N_in grid_clb_6__8_/prog_clk_0_W_out cby_6__8_/left_grid_pin_16_
+ cby_6__8_/left_grid_pin_17_ cby_6__8_/left_grid_pin_18_ cby_6__8_/left_grid_pin_19_
+ cby_6__8_/left_grid_pin_20_ cby_6__8_/left_grid_pin_21_ cby_6__8_/left_grid_pin_22_
+ cby_6__8_/left_grid_pin_23_ cby_6__8_/left_grid_pin_24_ cby_6__8_/left_grid_pin_25_
+ cby_6__8_/left_grid_pin_26_ cby_6__8_/left_grid_pin_27_ cby_6__8_/left_grid_pin_28_
+ cby_6__8_/left_grid_pin_29_ cby_6__8_/left_grid_pin_30_ cby_6__8_/left_grid_pin_31_
+ sb_6__7_/top_left_grid_pin_42_ sb_6__8_/bottom_left_grid_pin_42_ sb_6__7_/top_left_grid_pin_43_
+ sb_6__8_/bottom_left_grid_pin_43_ sb_6__7_/top_left_grid_pin_44_ sb_6__8_/bottom_left_grid_pin_44_
+ sb_6__7_/top_left_grid_pin_45_ sb_6__8_/bottom_left_grid_pin_45_ sb_6__7_/top_left_grid_pin_46_
+ sb_6__8_/bottom_left_grid_pin_46_ sb_6__7_/top_left_grid_pin_47_ sb_6__8_/bottom_left_grid_pin_47_
+ sb_6__7_/top_left_grid_pin_48_ sb_6__8_/bottom_left_grid_pin_48_ sb_6__7_/top_left_grid_pin_49_
+ sb_6__8_/bottom_left_grid_pin_49_ cbx_6__8_/bottom_grid_pin_0_ cbx_6__8_/bottom_grid_pin_10_
+ cbx_6__8_/bottom_grid_pin_11_ cbx_6__8_/bottom_grid_pin_12_ cbx_6__8_/bottom_grid_pin_13_
+ cbx_6__8_/bottom_grid_pin_14_ cbx_6__8_/bottom_grid_pin_15_ cbx_6__8_/bottom_grid_pin_1_
+ cbx_6__8_/bottom_grid_pin_2_ tie_array/x[5] grid_clb_6__8_/top_width_0_height_0__pin_33_
+ sb_6__8_/left_bottom_grid_pin_34_ sb_5__8_/right_bottom_grid_pin_34_ sb_6__8_/left_bottom_grid_pin_35_
+ sb_5__8_/right_bottom_grid_pin_35_ sb_6__8_/left_bottom_grid_pin_36_ sb_5__8_/right_bottom_grid_pin_36_
+ sb_6__8_/left_bottom_grid_pin_37_ sb_5__8_/right_bottom_grid_pin_37_ sb_6__8_/left_bottom_grid_pin_38_
+ sb_5__8_/right_bottom_grid_pin_38_ sb_6__8_/left_bottom_grid_pin_39_ sb_5__8_/right_bottom_grid_pin_39_
+ cbx_6__8_/bottom_grid_pin_3_ sb_6__8_/left_bottom_grid_pin_40_ sb_5__8_/right_bottom_grid_pin_40_
+ sb_6__8_/left_bottom_grid_pin_41_ sb_5__8_/right_bottom_grid_pin_41_ cbx_6__8_/bottom_grid_pin_4_
+ cbx_6__8_/bottom_grid_pin_5_ cbx_6__8_/bottom_grid_pin_6_ cbx_6__8_/bottom_grid_pin_7_
+ cbx_6__8_/bottom_grid_pin_8_ cbx_6__8_/bottom_grid_pin_9_ grid_clb
Xcbx_4__5_ cbx_4__5_/REGIN_FEEDTHROUGH cbx_4__5_/REGOUT_FEEDTHROUGH cbx_4__5_/SC_IN_BOT
+ cbx_4__5_/SC_IN_TOP cbx_4__5_/SC_OUT_BOT cbx_4__5_/SC_OUT_TOP VGND VPWR cbx_4__5_/bottom_grid_pin_0_
+ cbx_4__5_/bottom_grid_pin_10_ cbx_4__5_/bottom_grid_pin_11_ cbx_4__5_/bottom_grid_pin_12_
+ cbx_4__5_/bottom_grid_pin_13_ cbx_4__5_/bottom_grid_pin_14_ cbx_4__5_/bottom_grid_pin_15_
+ cbx_4__5_/bottom_grid_pin_1_ cbx_4__5_/bottom_grid_pin_2_ cbx_4__5_/bottom_grid_pin_3_
+ cbx_4__5_/bottom_grid_pin_4_ cbx_4__5_/bottom_grid_pin_5_ cbx_4__5_/bottom_grid_pin_6_
+ cbx_4__5_/bottom_grid_pin_7_ cbx_4__5_/bottom_grid_pin_8_ cbx_4__5_/bottom_grid_pin_9_
+ sb_4__5_/ccff_tail sb_3__5_/ccff_head cbx_4__5_/chanx_left_in[0] cbx_4__5_/chanx_left_in[10]
+ cbx_4__5_/chanx_left_in[11] cbx_4__5_/chanx_left_in[12] cbx_4__5_/chanx_left_in[13]
+ cbx_4__5_/chanx_left_in[14] cbx_4__5_/chanx_left_in[15] cbx_4__5_/chanx_left_in[16]
+ cbx_4__5_/chanx_left_in[17] cbx_4__5_/chanx_left_in[18] cbx_4__5_/chanx_left_in[19]
+ cbx_4__5_/chanx_left_in[1] cbx_4__5_/chanx_left_in[2] cbx_4__5_/chanx_left_in[3]
+ cbx_4__5_/chanx_left_in[4] cbx_4__5_/chanx_left_in[5] cbx_4__5_/chanx_left_in[6]
+ cbx_4__5_/chanx_left_in[7] cbx_4__5_/chanx_left_in[8] cbx_4__5_/chanx_left_in[9]
+ sb_3__5_/chanx_right_in[0] sb_3__5_/chanx_right_in[10] sb_3__5_/chanx_right_in[11]
+ sb_3__5_/chanx_right_in[12] sb_3__5_/chanx_right_in[13] sb_3__5_/chanx_right_in[14]
+ sb_3__5_/chanx_right_in[15] sb_3__5_/chanx_right_in[16] sb_3__5_/chanx_right_in[17]
+ sb_3__5_/chanx_right_in[18] sb_3__5_/chanx_right_in[19] sb_3__5_/chanx_right_in[1]
+ sb_3__5_/chanx_right_in[2] sb_3__5_/chanx_right_in[3] sb_3__5_/chanx_right_in[4]
+ sb_3__5_/chanx_right_in[5] sb_3__5_/chanx_right_in[6] sb_3__5_/chanx_right_in[7]
+ sb_3__5_/chanx_right_in[8] sb_3__5_/chanx_right_in[9] sb_4__5_/chanx_left_out[0]
+ sb_4__5_/chanx_left_out[10] sb_4__5_/chanx_left_out[11] sb_4__5_/chanx_left_out[12]
+ sb_4__5_/chanx_left_out[13] sb_4__5_/chanx_left_out[14] sb_4__5_/chanx_left_out[15]
+ sb_4__5_/chanx_left_out[16] sb_4__5_/chanx_left_out[17] sb_4__5_/chanx_left_out[18]
+ sb_4__5_/chanx_left_out[19] sb_4__5_/chanx_left_out[1] sb_4__5_/chanx_left_out[2]
+ sb_4__5_/chanx_left_out[3] sb_4__5_/chanx_left_out[4] sb_4__5_/chanx_left_out[5]
+ sb_4__5_/chanx_left_out[6] sb_4__5_/chanx_left_out[7] sb_4__5_/chanx_left_out[8]
+ sb_4__5_/chanx_left_out[9] sb_4__5_/chanx_left_in[0] sb_4__5_/chanx_left_in[10]
+ sb_4__5_/chanx_left_in[11] sb_4__5_/chanx_left_in[12] sb_4__5_/chanx_left_in[13]
+ sb_4__5_/chanx_left_in[14] sb_4__5_/chanx_left_in[15] sb_4__5_/chanx_left_in[16]
+ sb_4__5_/chanx_left_in[17] sb_4__5_/chanx_left_in[18] sb_4__5_/chanx_left_in[19]
+ sb_4__5_/chanx_left_in[1] sb_4__5_/chanx_left_in[2] sb_4__5_/chanx_left_in[3] sb_4__5_/chanx_left_in[4]
+ sb_4__5_/chanx_left_in[5] sb_4__5_/chanx_left_in[6] sb_4__5_/chanx_left_in[7] sb_4__5_/chanx_left_in[8]
+ sb_4__5_/chanx_left_in[9] cbx_4__5_/clk_1_N_out cbx_4__5_/clk_1_S_out sb_3__5_/clk_1_E_out
+ cbx_4__5_/clk_2_E_out cbx_4__5_/clk_2_W_in cbx_4__5_/clk_2_W_out cbx_4__5_/clk_3_E_out
+ cbx_4__5_/clk_3_W_in cbx_4__5_/clk_3_W_out cbx_4__5_/prog_clk_0_N_in cbx_4__5_/prog_clk_0_W_out
+ cbx_4__5_/prog_clk_1_N_out cbx_4__5_/prog_clk_1_S_out sb_3__5_/prog_clk_1_E_out
+ cbx_4__5_/prog_clk_2_E_out cbx_4__5_/prog_clk_2_W_in cbx_4__5_/prog_clk_2_W_out
+ cbx_4__5_/prog_clk_3_E_out cbx_4__5_/prog_clk_3_W_in cbx_4__5_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_3__5_ cbx_3__5_/SC_OUT_BOT cbx_3__4_/SC_IN_TOP grid_clb_3__5_/SC_OUT_TOP
+ cby_3__5_/Test_en_W_out grid_clb_3__5_/Test_en_E_out cby_3__5_/Test_en_W_out cby_2__5_/Test_en_W_in
+ VGND VPWR cbx_3__4_/REGIN_FEEDTHROUGH grid_clb_3__5_/bottom_width_0_height_0__pin_51_
+ cby_2__5_/ccff_tail cby_3__5_/ccff_head cbx_3__5_/clk_1_S_out cbx_3__5_/clk_1_S_out
+ cby_3__5_/prog_clk_0_W_in cbx_3__5_/prog_clk_1_S_out grid_clb_3__5_/prog_clk_0_N_out
+ cbx_3__5_/prog_clk_1_S_out cbx_3__4_/prog_clk_0_N_in grid_clb_3__5_/prog_clk_0_W_out
+ cby_3__5_/left_grid_pin_16_ cby_3__5_/left_grid_pin_17_ cby_3__5_/left_grid_pin_18_
+ cby_3__5_/left_grid_pin_19_ cby_3__5_/left_grid_pin_20_ cby_3__5_/left_grid_pin_21_
+ cby_3__5_/left_grid_pin_22_ cby_3__5_/left_grid_pin_23_ cby_3__5_/left_grid_pin_24_
+ cby_3__5_/left_grid_pin_25_ cby_3__5_/left_grid_pin_26_ cby_3__5_/left_grid_pin_27_
+ cby_3__5_/left_grid_pin_28_ cby_3__5_/left_grid_pin_29_ cby_3__5_/left_grid_pin_30_
+ cby_3__5_/left_grid_pin_31_ sb_3__4_/top_left_grid_pin_42_ sb_3__5_/bottom_left_grid_pin_42_
+ sb_3__4_/top_left_grid_pin_43_ sb_3__5_/bottom_left_grid_pin_43_ sb_3__4_/top_left_grid_pin_44_
+ sb_3__5_/bottom_left_grid_pin_44_ sb_3__4_/top_left_grid_pin_45_ sb_3__5_/bottom_left_grid_pin_45_
+ sb_3__4_/top_left_grid_pin_46_ sb_3__5_/bottom_left_grid_pin_46_ sb_3__4_/top_left_grid_pin_47_
+ sb_3__5_/bottom_left_grid_pin_47_ sb_3__4_/top_left_grid_pin_48_ sb_3__5_/bottom_left_grid_pin_48_
+ sb_3__4_/top_left_grid_pin_49_ sb_3__5_/bottom_left_grid_pin_49_ cbx_3__5_/bottom_grid_pin_0_
+ cbx_3__5_/bottom_grid_pin_10_ cbx_3__5_/bottom_grid_pin_11_ cbx_3__5_/bottom_grid_pin_12_
+ cbx_3__5_/bottom_grid_pin_13_ cbx_3__5_/bottom_grid_pin_14_ cbx_3__5_/bottom_grid_pin_15_
+ cbx_3__5_/bottom_grid_pin_1_ cbx_3__5_/bottom_grid_pin_2_ cbx_3__5_/REGOUT_FEEDTHROUGH
+ grid_clb_3__5_/top_width_0_height_0__pin_33_ sb_3__5_/left_bottom_grid_pin_34_ sb_2__5_/right_bottom_grid_pin_34_
+ sb_3__5_/left_bottom_grid_pin_35_ sb_2__5_/right_bottom_grid_pin_35_ sb_3__5_/left_bottom_grid_pin_36_
+ sb_2__5_/right_bottom_grid_pin_36_ sb_3__5_/left_bottom_grid_pin_37_ sb_2__5_/right_bottom_grid_pin_37_
+ sb_3__5_/left_bottom_grid_pin_38_ sb_2__5_/right_bottom_grid_pin_38_ sb_3__5_/left_bottom_grid_pin_39_
+ sb_2__5_/right_bottom_grid_pin_39_ cbx_3__5_/bottom_grid_pin_3_ sb_3__5_/left_bottom_grid_pin_40_
+ sb_2__5_/right_bottom_grid_pin_40_ sb_3__5_/left_bottom_grid_pin_41_ sb_2__5_/right_bottom_grid_pin_41_
+ cbx_3__5_/bottom_grid_pin_4_ cbx_3__5_/bottom_grid_pin_5_ cbx_3__5_/bottom_grid_pin_6_
+ cbx_3__5_/bottom_grid_pin_7_ cbx_3__5_/bottom_grid_pin_8_ cbx_3__5_/bottom_grid_pin_9_
+ grid_clb
Xcbx_1__2_ cbx_1__2_/REGIN_FEEDTHROUGH cbx_1__2_/REGOUT_FEEDTHROUGH cbx_1__2_/SC_IN_BOT
+ cbx_1__2_/SC_IN_TOP cbx_1__2_/SC_OUT_BOT cbx_1__2_/SC_OUT_TOP VGND VPWR cbx_1__2_/bottom_grid_pin_0_
+ cbx_1__2_/bottom_grid_pin_10_ cbx_1__2_/bottom_grid_pin_11_ cbx_1__2_/bottom_grid_pin_12_
+ cbx_1__2_/bottom_grid_pin_13_ cbx_1__2_/bottom_grid_pin_14_ cbx_1__2_/bottom_grid_pin_15_
+ cbx_1__2_/bottom_grid_pin_1_ cbx_1__2_/bottom_grid_pin_2_ cbx_1__2_/bottom_grid_pin_3_
+ cbx_1__2_/bottom_grid_pin_4_ cbx_1__2_/bottom_grid_pin_5_ cbx_1__2_/bottom_grid_pin_6_
+ cbx_1__2_/bottom_grid_pin_7_ cbx_1__2_/bottom_grid_pin_8_ cbx_1__2_/bottom_grid_pin_9_
+ sb_1__2_/ccff_tail sb_0__2_/ccff_head cbx_1__2_/chanx_left_in[0] cbx_1__2_/chanx_left_in[10]
+ cbx_1__2_/chanx_left_in[11] cbx_1__2_/chanx_left_in[12] cbx_1__2_/chanx_left_in[13]
+ cbx_1__2_/chanx_left_in[14] cbx_1__2_/chanx_left_in[15] cbx_1__2_/chanx_left_in[16]
+ cbx_1__2_/chanx_left_in[17] cbx_1__2_/chanx_left_in[18] cbx_1__2_/chanx_left_in[19]
+ cbx_1__2_/chanx_left_in[1] cbx_1__2_/chanx_left_in[2] cbx_1__2_/chanx_left_in[3]
+ cbx_1__2_/chanx_left_in[4] cbx_1__2_/chanx_left_in[5] cbx_1__2_/chanx_left_in[6]
+ cbx_1__2_/chanx_left_in[7] cbx_1__2_/chanx_left_in[8] cbx_1__2_/chanx_left_in[9]
+ sb_0__2_/chanx_right_in[0] sb_0__2_/chanx_right_in[10] sb_0__2_/chanx_right_in[11]
+ sb_0__2_/chanx_right_in[12] sb_0__2_/chanx_right_in[13] sb_0__2_/chanx_right_in[14]
+ sb_0__2_/chanx_right_in[15] sb_0__2_/chanx_right_in[16] sb_0__2_/chanx_right_in[17]
+ sb_0__2_/chanx_right_in[18] sb_0__2_/chanx_right_in[19] sb_0__2_/chanx_right_in[1]
+ sb_0__2_/chanx_right_in[2] sb_0__2_/chanx_right_in[3] sb_0__2_/chanx_right_in[4]
+ sb_0__2_/chanx_right_in[5] sb_0__2_/chanx_right_in[6] sb_0__2_/chanx_right_in[7]
+ sb_0__2_/chanx_right_in[8] sb_0__2_/chanx_right_in[9] sb_1__2_/chanx_left_out[0]
+ sb_1__2_/chanx_left_out[10] sb_1__2_/chanx_left_out[11] sb_1__2_/chanx_left_out[12]
+ sb_1__2_/chanx_left_out[13] sb_1__2_/chanx_left_out[14] sb_1__2_/chanx_left_out[15]
+ sb_1__2_/chanx_left_out[16] sb_1__2_/chanx_left_out[17] sb_1__2_/chanx_left_out[18]
+ sb_1__2_/chanx_left_out[19] sb_1__2_/chanx_left_out[1] sb_1__2_/chanx_left_out[2]
+ sb_1__2_/chanx_left_out[3] sb_1__2_/chanx_left_out[4] sb_1__2_/chanx_left_out[5]
+ sb_1__2_/chanx_left_out[6] sb_1__2_/chanx_left_out[7] sb_1__2_/chanx_left_out[8]
+ sb_1__2_/chanx_left_out[9] sb_1__2_/chanx_left_in[0] sb_1__2_/chanx_left_in[10]
+ sb_1__2_/chanx_left_in[11] sb_1__2_/chanx_left_in[12] sb_1__2_/chanx_left_in[13]
+ sb_1__2_/chanx_left_in[14] sb_1__2_/chanx_left_in[15] sb_1__2_/chanx_left_in[16]
+ sb_1__2_/chanx_left_in[17] sb_1__2_/chanx_left_in[18] sb_1__2_/chanx_left_in[19]
+ sb_1__2_/chanx_left_in[1] sb_1__2_/chanx_left_in[2] sb_1__2_/chanx_left_in[3] sb_1__2_/chanx_left_in[4]
+ sb_1__2_/chanx_left_in[5] sb_1__2_/chanx_left_in[6] sb_1__2_/chanx_left_in[7] sb_1__2_/chanx_left_in[8]
+ sb_1__2_/chanx_left_in[9] cbx_1__2_/clk_1_N_out cbx_1__2_/clk_1_S_out cbx_1__2_/clk_1_W_in
+ cbx_1__2_/clk_2_E_out cbx_1__2_/clk_2_W_in cbx_1__2_/clk_2_W_out cbx_1__2_/clk_3_E_out
+ cbx_1__2_/clk_3_W_in cbx_1__2_/clk_3_W_out cbx_1__2_/prog_clk_0_N_in sb_0__2_/prog_clk_0_E_in
+ cbx_1__2_/prog_clk_1_N_out cbx_1__2_/prog_clk_1_S_out cbx_1__2_/prog_clk_1_W_in
+ cbx_1__2_/prog_clk_2_E_out cbx_1__2_/prog_clk_2_W_in cbx_1__2_/prog_clk_2_W_out
+ cbx_1__2_/prog_clk_3_E_out cbx_1__2_/prog_clk_3_W_in cbx_1__2_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_8__2_ VGND VPWR sb_8__2_/bottom_left_grid_pin_42_ sb_8__2_/bottom_left_grid_pin_43_
+ sb_8__2_/bottom_left_grid_pin_44_ sb_8__2_/bottom_left_grid_pin_45_ sb_8__2_/bottom_left_grid_pin_46_
+ sb_8__2_/bottom_left_grid_pin_47_ sb_8__2_/bottom_left_grid_pin_48_ sb_8__2_/bottom_left_grid_pin_49_
+ sb_8__2_/bottom_right_grid_pin_1_ sb_8__2_/ccff_head sb_8__2_/ccff_tail sb_8__2_/chanx_left_in[0]
+ sb_8__2_/chanx_left_in[10] sb_8__2_/chanx_left_in[11] sb_8__2_/chanx_left_in[12]
+ sb_8__2_/chanx_left_in[13] sb_8__2_/chanx_left_in[14] sb_8__2_/chanx_left_in[15]
+ sb_8__2_/chanx_left_in[16] sb_8__2_/chanx_left_in[17] sb_8__2_/chanx_left_in[18]
+ sb_8__2_/chanx_left_in[19] sb_8__2_/chanx_left_in[1] sb_8__2_/chanx_left_in[2] sb_8__2_/chanx_left_in[3]
+ sb_8__2_/chanx_left_in[4] sb_8__2_/chanx_left_in[5] sb_8__2_/chanx_left_in[6] sb_8__2_/chanx_left_in[7]
+ sb_8__2_/chanx_left_in[8] sb_8__2_/chanx_left_in[9] sb_8__2_/chanx_left_out[0] sb_8__2_/chanx_left_out[10]
+ sb_8__2_/chanx_left_out[11] sb_8__2_/chanx_left_out[12] sb_8__2_/chanx_left_out[13]
+ sb_8__2_/chanx_left_out[14] sb_8__2_/chanx_left_out[15] sb_8__2_/chanx_left_out[16]
+ sb_8__2_/chanx_left_out[17] sb_8__2_/chanx_left_out[18] sb_8__2_/chanx_left_out[19]
+ sb_8__2_/chanx_left_out[1] sb_8__2_/chanx_left_out[2] sb_8__2_/chanx_left_out[3]
+ sb_8__2_/chanx_left_out[4] sb_8__2_/chanx_left_out[5] sb_8__2_/chanx_left_out[6]
+ sb_8__2_/chanx_left_out[7] sb_8__2_/chanx_left_out[8] sb_8__2_/chanx_left_out[9]
+ cby_8__2_/chany_top_out[0] cby_8__2_/chany_top_out[10] cby_8__2_/chany_top_out[11]
+ cby_8__2_/chany_top_out[12] cby_8__2_/chany_top_out[13] cby_8__2_/chany_top_out[14]
+ cby_8__2_/chany_top_out[15] cby_8__2_/chany_top_out[16] cby_8__2_/chany_top_out[17]
+ cby_8__2_/chany_top_out[18] cby_8__2_/chany_top_out[19] cby_8__2_/chany_top_out[1]
+ cby_8__2_/chany_top_out[2] cby_8__2_/chany_top_out[3] cby_8__2_/chany_top_out[4]
+ cby_8__2_/chany_top_out[5] cby_8__2_/chany_top_out[6] cby_8__2_/chany_top_out[7]
+ cby_8__2_/chany_top_out[8] cby_8__2_/chany_top_out[9] cby_8__2_/chany_top_in[0]
+ cby_8__2_/chany_top_in[10] cby_8__2_/chany_top_in[11] cby_8__2_/chany_top_in[12]
+ cby_8__2_/chany_top_in[13] cby_8__2_/chany_top_in[14] cby_8__2_/chany_top_in[15]
+ cby_8__2_/chany_top_in[16] cby_8__2_/chany_top_in[17] cby_8__2_/chany_top_in[18]
+ cby_8__2_/chany_top_in[19] cby_8__2_/chany_top_in[1] cby_8__2_/chany_top_in[2] cby_8__2_/chany_top_in[3]
+ cby_8__2_/chany_top_in[4] cby_8__2_/chany_top_in[5] cby_8__2_/chany_top_in[6] cby_8__2_/chany_top_in[7]
+ cby_8__2_/chany_top_in[8] cby_8__2_/chany_top_in[9] sb_8__2_/chany_top_in[0] sb_8__2_/chany_top_in[10]
+ sb_8__2_/chany_top_in[11] sb_8__2_/chany_top_in[12] sb_8__2_/chany_top_in[13] sb_8__2_/chany_top_in[14]
+ sb_8__2_/chany_top_in[15] sb_8__2_/chany_top_in[16] sb_8__2_/chany_top_in[17] sb_8__2_/chany_top_in[18]
+ sb_8__2_/chany_top_in[19] sb_8__2_/chany_top_in[1] sb_8__2_/chany_top_in[2] sb_8__2_/chany_top_in[3]
+ sb_8__2_/chany_top_in[4] sb_8__2_/chany_top_in[5] sb_8__2_/chany_top_in[6] sb_8__2_/chany_top_in[7]
+ sb_8__2_/chany_top_in[8] sb_8__2_/chany_top_in[9] sb_8__2_/chany_top_out[0] sb_8__2_/chany_top_out[10]
+ sb_8__2_/chany_top_out[11] sb_8__2_/chany_top_out[12] sb_8__2_/chany_top_out[13]
+ sb_8__2_/chany_top_out[14] sb_8__2_/chany_top_out[15] sb_8__2_/chany_top_out[16]
+ sb_8__2_/chany_top_out[17] sb_8__2_/chany_top_out[18] sb_8__2_/chany_top_out[19]
+ sb_8__2_/chany_top_out[1] sb_8__2_/chany_top_out[2] sb_8__2_/chany_top_out[3] sb_8__2_/chany_top_out[4]
+ sb_8__2_/chany_top_out[5] sb_8__2_/chany_top_out[6] sb_8__2_/chany_top_out[7] sb_8__2_/chany_top_out[8]
+ sb_8__2_/chany_top_out[9] sb_8__2_/left_bottom_grid_pin_34_ sb_8__2_/left_bottom_grid_pin_35_
+ sb_8__2_/left_bottom_grid_pin_36_ sb_8__2_/left_bottom_grid_pin_37_ sb_8__2_/left_bottom_grid_pin_38_
+ sb_8__2_/left_bottom_grid_pin_39_ sb_8__2_/left_bottom_grid_pin_40_ sb_8__2_/left_bottom_grid_pin_41_
+ sb_8__2_/prog_clk_0_N_in sb_8__2_/top_left_grid_pin_42_ sb_8__2_/top_left_grid_pin_43_
+ sb_8__2_/top_left_grid_pin_44_ sb_8__2_/top_left_grid_pin_45_ sb_8__2_/top_left_grid_pin_46_
+ sb_8__2_/top_left_grid_pin_47_ sb_8__2_/top_left_grid_pin_48_ sb_8__2_/top_left_grid_pin_49_
+ sb_8__2_/top_right_grid_pin_1_ sb_2__1_
Xsb_1__7_ sb_1__7_/Test_en_N_out sb_1__7_/Test_en_S_in VGND VPWR sb_1__7_/bottom_left_grid_pin_42_
+ sb_1__7_/bottom_left_grid_pin_43_ sb_1__7_/bottom_left_grid_pin_44_ sb_1__7_/bottom_left_grid_pin_45_
+ sb_1__7_/bottom_left_grid_pin_46_ sb_1__7_/bottom_left_grid_pin_47_ sb_1__7_/bottom_left_grid_pin_48_
+ sb_1__7_/bottom_left_grid_pin_49_ sb_1__7_/ccff_head sb_1__7_/ccff_tail sb_1__7_/chanx_left_in[0]
+ sb_1__7_/chanx_left_in[10] sb_1__7_/chanx_left_in[11] sb_1__7_/chanx_left_in[12]
+ sb_1__7_/chanx_left_in[13] sb_1__7_/chanx_left_in[14] sb_1__7_/chanx_left_in[15]
+ sb_1__7_/chanx_left_in[16] sb_1__7_/chanx_left_in[17] sb_1__7_/chanx_left_in[18]
+ sb_1__7_/chanx_left_in[19] sb_1__7_/chanx_left_in[1] sb_1__7_/chanx_left_in[2] sb_1__7_/chanx_left_in[3]
+ sb_1__7_/chanx_left_in[4] sb_1__7_/chanx_left_in[5] sb_1__7_/chanx_left_in[6] sb_1__7_/chanx_left_in[7]
+ sb_1__7_/chanx_left_in[8] sb_1__7_/chanx_left_in[9] sb_1__7_/chanx_left_out[0] sb_1__7_/chanx_left_out[10]
+ sb_1__7_/chanx_left_out[11] sb_1__7_/chanx_left_out[12] sb_1__7_/chanx_left_out[13]
+ sb_1__7_/chanx_left_out[14] sb_1__7_/chanx_left_out[15] sb_1__7_/chanx_left_out[16]
+ sb_1__7_/chanx_left_out[17] sb_1__7_/chanx_left_out[18] sb_1__7_/chanx_left_out[19]
+ sb_1__7_/chanx_left_out[1] sb_1__7_/chanx_left_out[2] sb_1__7_/chanx_left_out[3]
+ sb_1__7_/chanx_left_out[4] sb_1__7_/chanx_left_out[5] sb_1__7_/chanx_left_out[6]
+ sb_1__7_/chanx_left_out[7] sb_1__7_/chanx_left_out[8] sb_1__7_/chanx_left_out[9]
+ sb_1__7_/chanx_right_in[0] sb_1__7_/chanx_right_in[10] sb_1__7_/chanx_right_in[11]
+ sb_1__7_/chanx_right_in[12] sb_1__7_/chanx_right_in[13] sb_1__7_/chanx_right_in[14]
+ sb_1__7_/chanx_right_in[15] sb_1__7_/chanx_right_in[16] sb_1__7_/chanx_right_in[17]
+ sb_1__7_/chanx_right_in[18] sb_1__7_/chanx_right_in[19] sb_1__7_/chanx_right_in[1]
+ sb_1__7_/chanx_right_in[2] sb_1__7_/chanx_right_in[3] sb_1__7_/chanx_right_in[4]
+ sb_1__7_/chanx_right_in[5] sb_1__7_/chanx_right_in[6] sb_1__7_/chanx_right_in[7]
+ sb_1__7_/chanx_right_in[8] sb_1__7_/chanx_right_in[9] cbx_2__7_/chanx_left_in[0]
+ cbx_2__7_/chanx_left_in[10] cbx_2__7_/chanx_left_in[11] cbx_2__7_/chanx_left_in[12]
+ cbx_2__7_/chanx_left_in[13] cbx_2__7_/chanx_left_in[14] cbx_2__7_/chanx_left_in[15]
+ cbx_2__7_/chanx_left_in[16] cbx_2__7_/chanx_left_in[17] cbx_2__7_/chanx_left_in[18]
+ cbx_2__7_/chanx_left_in[19] cbx_2__7_/chanx_left_in[1] cbx_2__7_/chanx_left_in[2]
+ cbx_2__7_/chanx_left_in[3] cbx_2__7_/chanx_left_in[4] cbx_2__7_/chanx_left_in[5]
+ cbx_2__7_/chanx_left_in[6] cbx_2__7_/chanx_left_in[7] cbx_2__7_/chanx_left_in[8]
+ cbx_2__7_/chanx_left_in[9] cby_1__7_/chany_top_out[0] cby_1__7_/chany_top_out[10]
+ cby_1__7_/chany_top_out[11] cby_1__7_/chany_top_out[12] cby_1__7_/chany_top_out[13]
+ cby_1__7_/chany_top_out[14] cby_1__7_/chany_top_out[15] cby_1__7_/chany_top_out[16]
+ cby_1__7_/chany_top_out[17] cby_1__7_/chany_top_out[18] cby_1__7_/chany_top_out[19]
+ cby_1__7_/chany_top_out[1] cby_1__7_/chany_top_out[2] cby_1__7_/chany_top_out[3]
+ cby_1__7_/chany_top_out[4] cby_1__7_/chany_top_out[5] cby_1__7_/chany_top_out[6]
+ cby_1__7_/chany_top_out[7] cby_1__7_/chany_top_out[8] cby_1__7_/chany_top_out[9]
+ cby_1__7_/chany_top_in[0] cby_1__7_/chany_top_in[10] cby_1__7_/chany_top_in[11]
+ cby_1__7_/chany_top_in[12] cby_1__7_/chany_top_in[13] cby_1__7_/chany_top_in[14]
+ cby_1__7_/chany_top_in[15] cby_1__7_/chany_top_in[16] cby_1__7_/chany_top_in[17]
+ cby_1__7_/chany_top_in[18] cby_1__7_/chany_top_in[19] cby_1__7_/chany_top_in[1]
+ cby_1__7_/chany_top_in[2] cby_1__7_/chany_top_in[3] cby_1__7_/chany_top_in[4] cby_1__7_/chany_top_in[5]
+ cby_1__7_/chany_top_in[6] cby_1__7_/chany_top_in[7] cby_1__7_/chany_top_in[8] cby_1__7_/chany_top_in[9]
+ sb_1__7_/chany_top_in[0] sb_1__7_/chany_top_in[10] sb_1__7_/chany_top_in[11] sb_1__7_/chany_top_in[12]
+ sb_1__7_/chany_top_in[13] sb_1__7_/chany_top_in[14] sb_1__7_/chany_top_in[15] sb_1__7_/chany_top_in[16]
+ sb_1__7_/chany_top_in[17] sb_1__7_/chany_top_in[18] sb_1__7_/chany_top_in[19] sb_1__7_/chany_top_in[1]
+ sb_1__7_/chany_top_in[2] sb_1__7_/chany_top_in[3] sb_1__7_/chany_top_in[4] sb_1__7_/chany_top_in[5]
+ sb_1__7_/chany_top_in[6] sb_1__7_/chany_top_in[7] sb_1__7_/chany_top_in[8] sb_1__7_/chany_top_in[9]
+ sb_1__7_/chany_top_out[0] sb_1__7_/chany_top_out[10] sb_1__7_/chany_top_out[11]
+ sb_1__7_/chany_top_out[12] sb_1__7_/chany_top_out[13] sb_1__7_/chany_top_out[14]
+ sb_1__7_/chany_top_out[15] sb_1__7_/chany_top_out[16] sb_1__7_/chany_top_out[17]
+ sb_1__7_/chany_top_out[18] sb_1__7_/chany_top_out[19] sb_1__7_/chany_top_out[1]
+ sb_1__7_/chany_top_out[2] sb_1__7_/chany_top_out[3] sb_1__7_/chany_top_out[4] sb_1__7_/chany_top_out[5]
+ sb_1__7_/chany_top_out[6] sb_1__7_/chany_top_out[7] sb_1__7_/chany_top_out[8] sb_1__7_/chany_top_out[9]
+ sb_1__7_/clk_1_E_out sb_1__7_/clk_1_N_in sb_1__7_/clk_1_W_out sb_1__7_/clk_2_E_out
+ sb_1__7_/clk_2_N_in sb_1__7_/clk_2_N_out sb_1__7_/clk_2_S_out sb_1__7_/clk_2_W_out
+ sb_1__7_/clk_3_E_out sb_1__7_/clk_3_N_in sb_1__7_/clk_3_N_out sb_1__7_/clk_3_S_out
+ sb_1__7_/clk_3_W_out sb_1__7_/left_bottom_grid_pin_34_ sb_1__7_/left_bottom_grid_pin_35_
+ sb_1__7_/left_bottom_grid_pin_36_ sb_1__7_/left_bottom_grid_pin_37_ sb_1__7_/left_bottom_grid_pin_38_
+ sb_1__7_/left_bottom_grid_pin_39_ sb_1__7_/left_bottom_grid_pin_40_ sb_1__7_/left_bottom_grid_pin_41_
+ sb_1__7_/prog_clk_0_N_in sb_1__7_/prog_clk_1_E_out sb_1__7_/prog_clk_1_N_in sb_1__7_/prog_clk_1_W_out
+ sb_1__7_/prog_clk_2_E_out sb_1__7_/prog_clk_2_N_in sb_1__7_/prog_clk_2_N_out sb_1__7_/prog_clk_2_S_out
+ sb_1__7_/prog_clk_2_W_out sb_1__7_/prog_clk_3_E_out sb_1__7_/prog_clk_3_N_in sb_1__7_/prog_clk_3_N_out
+ sb_1__7_/prog_clk_3_S_out sb_1__7_/prog_clk_3_W_out sb_1__7_/right_bottom_grid_pin_34_
+ sb_1__7_/right_bottom_grid_pin_35_ sb_1__7_/right_bottom_grid_pin_36_ sb_1__7_/right_bottom_grid_pin_37_
+ sb_1__7_/right_bottom_grid_pin_38_ sb_1__7_/right_bottom_grid_pin_39_ sb_1__7_/right_bottom_grid_pin_40_
+ sb_1__7_/right_bottom_grid_pin_41_ sb_1__7_/top_left_grid_pin_42_ sb_1__7_/top_left_grid_pin_43_
+ sb_1__7_/top_left_grid_pin_44_ sb_1__7_/top_left_grid_pin_45_ sb_1__7_/top_left_grid_pin_46_
+ sb_1__7_/top_left_grid_pin_47_ sb_1__7_/top_left_grid_pin_48_ sb_1__7_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_7__6_ cby_7__6_/Test_en_W_in cby_7__6_/Test_en_E_out cby_7__6_/Test_en_N_out
+ cby_7__6_/Test_en_W_in cby_7__6_/Test_en_W_in cby_7__6_/Test_en_W_out VGND VPWR
+ cby_7__6_/ccff_head cby_7__6_/ccff_tail sb_7__5_/chany_top_out[0] sb_7__5_/chany_top_out[10]
+ sb_7__5_/chany_top_out[11] sb_7__5_/chany_top_out[12] sb_7__5_/chany_top_out[13]
+ sb_7__5_/chany_top_out[14] sb_7__5_/chany_top_out[15] sb_7__5_/chany_top_out[16]
+ sb_7__5_/chany_top_out[17] sb_7__5_/chany_top_out[18] sb_7__5_/chany_top_out[19]
+ sb_7__5_/chany_top_out[1] sb_7__5_/chany_top_out[2] sb_7__5_/chany_top_out[3] sb_7__5_/chany_top_out[4]
+ sb_7__5_/chany_top_out[5] sb_7__5_/chany_top_out[6] sb_7__5_/chany_top_out[7] sb_7__5_/chany_top_out[8]
+ sb_7__5_/chany_top_out[9] sb_7__5_/chany_top_in[0] sb_7__5_/chany_top_in[10] sb_7__5_/chany_top_in[11]
+ sb_7__5_/chany_top_in[12] sb_7__5_/chany_top_in[13] sb_7__5_/chany_top_in[14] sb_7__5_/chany_top_in[15]
+ sb_7__5_/chany_top_in[16] sb_7__5_/chany_top_in[17] sb_7__5_/chany_top_in[18] sb_7__5_/chany_top_in[19]
+ sb_7__5_/chany_top_in[1] sb_7__5_/chany_top_in[2] sb_7__5_/chany_top_in[3] sb_7__5_/chany_top_in[4]
+ sb_7__5_/chany_top_in[5] sb_7__5_/chany_top_in[6] sb_7__5_/chany_top_in[7] sb_7__5_/chany_top_in[8]
+ sb_7__5_/chany_top_in[9] cby_7__6_/chany_top_in[0] cby_7__6_/chany_top_in[10] cby_7__6_/chany_top_in[11]
+ cby_7__6_/chany_top_in[12] cby_7__6_/chany_top_in[13] cby_7__6_/chany_top_in[14]
+ cby_7__6_/chany_top_in[15] cby_7__6_/chany_top_in[16] cby_7__6_/chany_top_in[17]
+ cby_7__6_/chany_top_in[18] cby_7__6_/chany_top_in[19] cby_7__6_/chany_top_in[1]
+ cby_7__6_/chany_top_in[2] cby_7__6_/chany_top_in[3] cby_7__6_/chany_top_in[4] cby_7__6_/chany_top_in[5]
+ cby_7__6_/chany_top_in[6] cby_7__6_/chany_top_in[7] cby_7__6_/chany_top_in[8] cby_7__6_/chany_top_in[9]
+ cby_7__6_/chany_top_out[0] cby_7__6_/chany_top_out[10] cby_7__6_/chany_top_out[11]
+ cby_7__6_/chany_top_out[12] cby_7__6_/chany_top_out[13] cby_7__6_/chany_top_out[14]
+ cby_7__6_/chany_top_out[15] cby_7__6_/chany_top_out[16] cby_7__6_/chany_top_out[17]
+ cby_7__6_/chany_top_out[18] cby_7__6_/chany_top_out[19] cby_7__6_/chany_top_out[1]
+ cby_7__6_/chany_top_out[2] cby_7__6_/chany_top_out[3] cby_7__6_/chany_top_out[4]
+ cby_7__6_/chany_top_out[5] cby_7__6_/chany_top_out[6] cby_7__6_/chany_top_out[7]
+ cby_7__6_/chany_top_out[8] cby_7__6_/chany_top_out[9] cby_7__6_/clk_2_N_out sb_7__6_/clk_2_S_out
+ sb_7__5_/clk_1_N_in cby_7__6_/clk_3_N_out cby_7__6_/clk_3_S_in cby_7__6_/clk_3_S_out
+ cby_7__6_/left_grid_pin_16_ cby_7__6_/left_grid_pin_17_ cby_7__6_/left_grid_pin_18_
+ cby_7__6_/left_grid_pin_19_ cby_7__6_/left_grid_pin_20_ cby_7__6_/left_grid_pin_21_
+ cby_7__6_/left_grid_pin_22_ cby_7__6_/left_grid_pin_23_ cby_7__6_/left_grid_pin_24_
+ cby_7__6_/left_grid_pin_25_ cby_7__6_/left_grid_pin_26_ cby_7__6_/left_grid_pin_27_
+ cby_7__6_/left_grid_pin_28_ cby_7__6_/left_grid_pin_29_ cby_7__6_/left_grid_pin_30_
+ cby_7__6_/left_grid_pin_31_ cby_7__6_/prog_clk_0_N_out sb_7__5_/prog_clk_0_N_in
+ cby_7__6_/prog_clk_0_W_in cby_7__6_/prog_clk_2_N_out sb_7__6_/prog_clk_2_S_out sb_7__5_/prog_clk_1_N_in
+ cby_7__6_/prog_clk_3_N_out cby_7__6_/prog_clk_3_S_in cby_7__6_/prog_clk_3_S_out
+ cby_1__1_
Xcby_4__3_ sb_4__2_/Test_en_N_out cby_4__3_/Test_en_E_out sb_4__3_/Test_en_S_in sb_4__2_/Test_en_N_out
+ sb_4__2_/Test_en_N_out cby_4__3_/Test_en_W_out VGND VPWR cby_4__3_/ccff_head cby_4__3_/ccff_tail
+ sb_4__2_/chany_top_out[0] sb_4__2_/chany_top_out[10] sb_4__2_/chany_top_out[11]
+ sb_4__2_/chany_top_out[12] sb_4__2_/chany_top_out[13] sb_4__2_/chany_top_out[14]
+ sb_4__2_/chany_top_out[15] sb_4__2_/chany_top_out[16] sb_4__2_/chany_top_out[17]
+ sb_4__2_/chany_top_out[18] sb_4__2_/chany_top_out[19] sb_4__2_/chany_top_out[1]
+ sb_4__2_/chany_top_out[2] sb_4__2_/chany_top_out[3] sb_4__2_/chany_top_out[4] sb_4__2_/chany_top_out[5]
+ sb_4__2_/chany_top_out[6] sb_4__2_/chany_top_out[7] sb_4__2_/chany_top_out[8] sb_4__2_/chany_top_out[9]
+ sb_4__2_/chany_top_in[0] sb_4__2_/chany_top_in[10] sb_4__2_/chany_top_in[11] sb_4__2_/chany_top_in[12]
+ sb_4__2_/chany_top_in[13] sb_4__2_/chany_top_in[14] sb_4__2_/chany_top_in[15] sb_4__2_/chany_top_in[16]
+ sb_4__2_/chany_top_in[17] sb_4__2_/chany_top_in[18] sb_4__2_/chany_top_in[19] sb_4__2_/chany_top_in[1]
+ sb_4__2_/chany_top_in[2] sb_4__2_/chany_top_in[3] sb_4__2_/chany_top_in[4] sb_4__2_/chany_top_in[5]
+ sb_4__2_/chany_top_in[6] sb_4__2_/chany_top_in[7] sb_4__2_/chany_top_in[8] sb_4__2_/chany_top_in[9]
+ cby_4__3_/chany_top_in[0] cby_4__3_/chany_top_in[10] cby_4__3_/chany_top_in[11]
+ cby_4__3_/chany_top_in[12] cby_4__3_/chany_top_in[13] cby_4__3_/chany_top_in[14]
+ cby_4__3_/chany_top_in[15] cby_4__3_/chany_top_in[16] cby_4__3_/chany_top_in[17]
+ cby_4__3_/chany_top_in[18] cby_4__3_/chany_top_in[19] cby_4__3_/chany_top_in[1]
+ cby_4__3_/chany_top_in[2] cby_4__3_/chany_top_in[3] cby_4__3_/chany_top_in[4] cby_4__3_/chany_top_in[5]
+ cby_4__3_/chany_top_in[6] cby_4__3_/chany_top_in[7] cby_4__3_/chany_top_in[8] cby_4__3_/chany_top_in[9]
+ cby_4__3_/chany_top_out[0] cby_4__3_/chany_top_out[10] cby_4__3_/chany_top_out[11]
+ cby_4__3_/chany_top_out[12] cby_4__3_/chany_top_out[13] cby_4__3_/chany_top_out[14]
+ cby_4__3_/chany_top_out[15] cby_4__3_/chany_top_out[16] cby_4__3_/chany_top_out[17]
+ cby_4__3_/chany_top_out[18] cby_4__3_/chany_top_out[19] cby_4__3_/chany_top_out[1]
+ cby_4__3_/chany_top_out[2] cby_4__3_/chany_top_out[3] cby_4__3_/chany_top_out[4]
+ cby_4__3_/chany_top_out[5] cby_4__3_/chany_top_out[6] cby_4__3_/chany_top_out[7]
+ cby_4__3_/chany_top_out[8] cby_4__3_/chany_top_out[9] cby_4__3_/clk_2_N_out cby_4__3_/clk_2_S_in
+ cby_4__3_/clk_2_S_out sb_4__3_/clk_3_N_in sb_4__2_/clk_3_N_out cby_4__3_/clk_3_S_out
+ cby_4__3_/left_grid_pin_16_ cby_4__3_/left_grid_pin_17_ cby_4__3_/left_grid_pin_18_
+ cby_4__3_/left_grid_pin_19_ cby_4__3_/left_grid_pin_20_ cby_4__3_/left_grid_pin_21_
+ cby_4__3_/left_grid_pin_22_ cby_4__3_/left_grid_pin_23_ cby_4__3_/left_grid_pin_24_
+ cby_4__3_/left_grid_pin_25_ cby_4__3_/left_grid_pin_26_ cby_4__3_/left_grid_pin_27_
+ cby_4__3_/left_grid_pin_28_ cby_4__3_/left_grid_pin_29_ cby_4__3_/left_grid_pin_30_
+ cby_4__3_/left_grid_pin_31_ cby_4__3_/prog_clk_0_N_out sb_4__2_/prog_clk_0_N_in
+ cby_4__3_/prog_clk_0_W_in cby_4__3_/prog_clk_2_N_out cby_4__3_/prog_clk_2_S_in cby_4__3_/prog_clk_2_S_out
+ sb_4__3_/prog_clk_3_N_in sb_4__2_/prog_clk_3_N_out cby_4__3_/prog_clk_3_S_out cby_1__1_
Xcbx_7__7_ cbx_7__7_/REGIN_FEEDTHROUGH cbx_7__7_/REGOUT_FEEDTHROUGH cbx_7__7_/SC_IN_BOT
+ cbx_7__7_/SC_IN_TOP cbx_7__7_/SC_OUT_BOT cbx_7__7_/SC_OUT_TOP VGND VPWR cbx_7__7_/bottom_grid_pin_0_
+ cbx_7__7_/bottom_grid_pin_10_ cbx_7__7_/bottom_grid_pin_11_ cbx_7__7_/bottom_grid_pin_12_
+ cbx_7__7_/bottom_grid_pin_13_ cbx_7__7_/bottom_grid_pin_14_ cbx_7__7_/bottom_grid_pin_15_
+ cbx_7__7_/bottom_grid_pin_1_ cbx_7__7_/bottom_grid_pin_2_ cbx_7__7_/bottom_grid_pin_3_
+ cbx_7__7_/bottom_grid_pin_4_ cbx_7__7_/bottom_grid_pin_5_ cbx_7__7_/bottom_grid_pin_6_
+ cbx_7__7_/bottom_grid_pin_7_ cbx_7__7_/bottom_grid_pin_8_ cbx_7__7_/bottom_grid_pin_9_
+ sb_7__7_/ccff_tail sb_6__7_/ccff_head cbx_7__7_/chanx_left_in[0] cbx_7__7_/chanx_left_in[10]
+ cbx_7__7_/chanx_left_in[11] cbx_7__7_/chanx_left_in[12] cbx_7__7_/chanx_left_in[13]
+ cbx_7__7_/chanx_left_in[14] cbx_7__7_/chanx_left_in[15] cbx_7__7_/chanx_left_in[16]
+ cbx_7__7_/chanx_left_in[17] cbx_7__7_/chanx_left_in[18] cbx_7__7_/chanx_left_in[19]
+ cbx_7__7_/chanx_left_in[1] cbx_7__7_/chanx_left_in[2] cbx_7__7_/chanx_left_in[3]
+ cbx_7__7_/chanx_left_in[4] cbx_7__7_/chanx_left_in[5] cbx_7__7_/chanx_left_in[6]
+ cbx_7__7_/chanx_left_in[7] cbx_7__7_/chanx_left_in[8] cbx_7__7_/chanx_left_in[9]
+ sb_6__7_/chanx_right_in[0] sb_6__7_/chanx_right_in[10] sb_6__7_/chanx_right_in[11]
+ sb_6__7_/chanx_right_in[12] sb_6__7_/chanx_right_in[13] sb_6__7_/chanx_right_in[14]
+ sb_6__7_/chanx_right_in[15] sb_6__7_/chanx_right_in[16] sb_6__7_/chanx_right_in[17]
+ sb_6__7_/chanx_right_in[18] sb_6__7_/chanx_right_in[19] sb_6__7_/chanx_right_in[1]
+ sb_6__7_/chanx_right_in[2] sb_6__7_/chanx_right_in[3] sb_6__7_/chanx_right_in[4]
+ sb_6__7_/chanx_right_in[5] sb_6__7_/chanx_right_in[6] sb_6__7_/chanx_right_in[7]
+ sb_6__7_/chanx_right_in[8] sb_6__7_/chanx_right_in[9] sb_7__7_/chanx_left_out[0]
+ sb_7__7_/chanx_left_out[10] sb_7__7_/chanx_left_out[11] sb_7__7_/chanx_left_out[12]
+ sb_7__7_/chanx_left_out[13] sb_7__7_/chanx_left_out[14] sb_7__7_/chanx_left_out[15]
+ sb_7__7_/chanx_left_out[16] sb_7__7_/chanx_left_out[17] sb_7__7_/chanx_left_out[18]
+ sb_7__7_/chanx_left_out[19] sb_7__7_/chanx_left_out[1] sb_7__7_/chanx_left_out[2]
+ sb_7__7_/chanx_left_out[3] sb_7__7_/chanx_left_out[4] sb_7__7_/chanx_left_out[5]
+ sb_7__7_/chanx_left_out[6] sb_7__7_/chanx_left_out[7] sb_7__7_/chanx_left_out[8]
+ sb_7__7_/chanx_left_out[9] sb_7__7_/chanx_left_in[0] sb_7__7_/chanx_left_in[10]
+ sb_7__7_/chanx_left_in[11] sb_7__7_/chanx_left_in[12] sb_7__7_/chanx_left_in[13]
+ sb_7__7_/chanx_left_in[14] sb_7__7_/chanx_left_in[15] sb_7__7_/chanx_left_in[16]
+ sb_7__7_/chanx_left_in[17] sb_7__7_/chanx_left_in[18] sb_7__7_/chanx_left_in[19]
+ sb_7__7_/chanx_left_in[1] sb_7__7_/chanx_left_in[2] sb_7__7_/chanx_left_in[3] sb_7__7_/chanx_left_in[4]
+ sb_7__7_/chanx_left_in[5] sb_7__7_/chanx_left_in[6] sb_7__7_/chanx_left_in[7] sb_7__7_/chanx_left_in[8]
+ sb_7__7_/chanx_left_in[9] cbx_7__7_/clk_1_N_out cbx_7__7_/clk_1_S_out sb_7__7_/clk_1_W_out
+ cbx_7__7_/clk_2_E_out cbx_7__7_/clk_2_W_in cbx_7__7_/clk_2_W_out cbx_7__7_/clk_3_E_out
+ cbx_7__7_/clk_3_W_in cbx_7__7_/clk_3_W_out cbx_7__7_/prog_clk_0_N_in cbx_7__7_/prog_clk_0_W_out
+ cbx_7__7_/prog_clk_1_N_out cbx_7__7_/prog_clk_1_S_out sb_7__7_/prog_clk_1_W_out
+ cbx_7__7_/prog_clk_2_E_out cbx_7__7_/prog_clk_2_W_in cbx_7__7_/prog_clk_2_W_out
+ cbx_7__7_/prog_clk_3_E_out cbx_7__7_/prog_clk_3_W_in cbx_7__7_/prog_clk_3_W_out
+ cbx_1__1_
Xcbx_4__4_ cbx_4__4_/REGIN_FEEDTHROUGH cbx_4__4_/REGOUT_FEEDTHROUGH cbx_4__4_/SC_IN_BOT
+ cbx_4__4_/SC_IN_TOP cbx_4__4_/SC_OUT_BOT cbx_4__4_/SC_OUT_TOP VGND VPWR cbx_4__4_/bottom_grid_pin_0_
+ cbx_4__4_/bottom_grid_pin_10_ cbx_4__4_/bottom_grid_pin_11_ cbx_4__4_/bottom_grid_pin_12_
+ cbx_4__4_/bottom_grid_pin_13_ cbx_4__4_/bottom_grid_pin_14_ cbx_4__4_/bottom_grid_pin_15_
+ cbx_4__4_/bottom_grid_pin_1_ cbx_4__4_/bottom_grid_pin_2_ cbx_4__4_/bottom_grid_pin_3_
+ cbx_4__4_/bottom_grid_pin_4_ cbx_4__4_/bottom_grid_pin_5_ cbx_4__4_/bottom_grid_pin_6_
+ cbx_4__4_/bottom_grid_pin_7_ cbx_4__4_/bottom_grid_pin_8_ cbx_4__4_/bottom_grid_pin_9_
+ sb_4__4_/ccff_tail sb_3__4_/ccff_head cbx_4__4_/chanx_left_in[0] cbx_4__4_/chanx_left_in[10]
+ cbx_4__4_/chanx_left_in[11] cbx_4__4_/chanx_left_in[12] cbx_4__4_/chanx_left_in[13]
+ cbx_4__4_/chanx_left_in[14] cbx_4__4_/chanx_left_in[15] cbx_4__4_/chanx_left_in[16]
+ cbx_4__4_/chanx_left_in[17] cbx_4__4_/chanx_left_in[18] cbx_4__4_/chanx_left_in[19]
+ cbx_4__4_/chanx_left_in[1] cbx_4__4_/chanx_left_in[2] cbx_4__4_/chanx_left_in[3]
+ cbx_4__4_/chanx_left_in[4] cbx_4__4_/chanx_left_in[5] cbx_4__4_/chanx_left_in[6]
+ cbx_4__4_/chanx_left_in[7] cbx_4__4_/chanx_left_in[8] cbx_4__4_/chanx_left_in[9]
+ sb_3__4_/chanx_right_in[0] sb_3__4_/chanx_right_in[10] sb_3__4_/chanx_right_in[11]
+ sb_3__4_/chanx_right_in[12] sb_3__4_/chanx_right_in[13] sb_3__4_/chanx_right_in[14]
+ sb_3__4_/chanx_right_in[15] sb_3__4_/chanx_right_in[16] sb_3__4_/chanx_right_in[17]
+ sb_3__4_/chanx_right_in[18] sb_3__4_/chanx_right_in[19] sb_3__4_/chanx_right_in[1]
+ sb_3__4_/chanx_right_in[2] sb_3__4_/chanx_right_in[3] sb_3__4_/chanx_right_in[4]
+ sb_3__4_/chanx_right_in[5] sb_3__4_/chanx_right_in[6] sb_3__4_/chanx_right_in[7]
+ sb_3__4_/chanx_right_in[8] sb_3__4_/chanx_right_in[9] sb_4__4_/chanx_left_out[0]
+ sb_4__4_/chanx_left_out[10] sb_4__4_/chanx_left_out[11] sb_4__4_/chanx_left_out[12]
+ sb_4__4_/chanx_left_out[13] sb_4__4_/chanx_left_out[14] sb_4__4_/chanx_left_out[15]
+ sb_4__4_/chanx_left_out[16] sb_4__4_/chanx_left_out[17] sb_4__4_/chanx_left_out[18]
+ sb_4__4_/chanx_left_out[19] sb_4__4_/chanx_left_out[1] sb_4__4_/chanx_left_out[2]
+ sb_4__4_/chanx_left_out[3] sb_4__4_/chanx_left_out[4] sb_4__4_/chanx_left_out[5]
+ sb_4__4_/chanx_left_out[6] sb_4__4_/chanx_left_out[7] sb_4__4_/chanx_left_out[8]
+ sb_4__4_/chanx_left_out[9] sb_4__4_/chanx_left_in[0] sb_4__4_/chanx_left_in[10]
+ sb_4__4_/chanx_left_in[11] sb_4__4_/chanx_left_in[12] sb_4__4_/chanx_left_in[13]
+ sb_4__4_/chanx_left_in[14] sb_4__4_/chanx_left_in[15] sb_4__4_/chanx_left_in[16]
+ sb_4__4_/chanx_left_in[17] sb_4__4_/chanx_left_in[18] sb_4__4_/chanx_left_in[19]
+ sb_4__4_/chanx_left_in[1] sb_4__4_/chanx_left_in[2] sb_4__4_/chanx_left_in[3] sb_4__4_/chanx_left_in[4]
+ sb_4__4_/chanx_left_in[5] sb_4__4_/chanx_left_in[6] sb_4__4_/chanx_left_in[7] sb_4__4_/chanx_left_in[8]
+ sb_4__4_/chanx_left_in[9] cbx_4__4_/clk_1_N_out cbx_4__4_/clk_1_S_out cbx_4__4_/clk_1_W_in
+ cbx_4__4_/clk_2_E_out cbx_4__4_/clk_2_W_in cbx_4__4_/clk_2_W_out cbx_4__4_/clk_3_E_out
+ sb_4__4_/clk_3_W_out sb_3__4_/clk_3_N_in cbx_4__4_/prog_clk_0_N_in cbx_4__4_/prog_clk_0_W_out
+ cbx_4__4_/prog_clk_1_N_out cbx_4__4_/prog_clk_1_S_out cbx_4__4_/prog_clk_1_W_in
+ cbx_4__4_/prog_clk_2_E_out cbx_4__4_/prog_clk_2_W_in cbx_4__4_/prog_clk_2_W_out
+ cbx_4__4_/prog_clk_3_E_out sb_4__4_/prog_clk_3_W_out sb_3__4_/prog_clk_3_N_in cbx_1__1_
Xgrid_clb_6__7_ cbx_6__6_/SC_OUT_TOP grid_clb_6__7_/SC_OUT_BOT cbx_6__7_/SC_IN_BOT
+ cby_5__7_/Test_en_E_out cby_6__7_/Test_en_W_in cby_5__7_/Test_en_E_out grid_clb_6__7_/Test_en_W_out
+ VGND VPWR cbx_6__6_/REGIN_FEEDTHROUGH grid_clb_6__7_/bottom_width_0_height_0__pin_51_
+ cby_5__7_/ccff_tail cby_6__7_/ccff_head cbx_6__7_/clk_1_S_out cbx_6__7_/clk_1_S_out
+ cby_6__7_/prog_clk_0_W_in cbx_6__7_/prog_clk_1_S_out grid_clb_6__7_/prog_clk_0_N_out
+ cbx_6__7_/prog_clk_1_S_out cbx_6__6_/prog_clk_0_N_in grid_clb_6__7_/prog_clk_0_W_out
+ cby_6__7_/left_grid_pin_16_ cby_6__7_/left_grid_pin_17_ cby_6__7_/left_grid_pin_18_
+ cby_6__7_/left_grid_pin_19_ cby_6__7_/left_grid_pin_20_ cby_6__7_/left_grid_pin_21_
+ cby_6__7_/left_grid_pin_22_ cby_6__7_/left_grid_pin_23_ cby_6__7_/left_grid_pin_24_
+ cby_6__7_/left_grid_pin_25_ cby_6__7_/left_grid_pin_26_ cby_6__7_/left_grid_pin_27_
+ cby_6__7_/left_grid_pin_28_ cby_6__7_/left_grid_pin_29_ cby_6__7_/left_grid_pin_30_
+ cby_6__7_/left_grid_pin_31_ sb_6__6_/top_left_grid_pin_42_ sb_6__7_/bottom_left_grid_pin_42_
+ sb_6__6_/top_left_grid_pin_43_ sb_6__7_/bottom_left_grid_pin_43_ sb_6__6_/top_left_grid_pin_44_
+ sb_6__7_/bottom_left_grid_pin_44_ sb_6__6_/top_left_grid_pin_45_ sb_6__7_/bottom_left_grid_pin_45_
+ sb_6__6_/top_left_grid_pin_46_ sb_6__7_/bottom_left_grid_pin_46_ sb_6__6_/top_left_grid_pin_47_
+ sb_6__7_/bottom_left_grid_pin_47_ sb_6__6_/top_left_grid_pin_48_ sb_6__7_/bottom_left_grid_pin_48_
+ sb_6__6_/top_left_grid_pin_49_ sb_6__7_/bottom_left_grid_pin_49_ cbx_6__7_/bottom_grid_pin_0_
+ cbx_6__7_/bottom_grid_pin_10_ cbx_6__7_/bottom_grid_pin_11_ cbx_6__7_/bottom_grid_pin_12_
+ cbx_6__7_/bottom_grid_pin_13_ cbx_6__7_/bottom_grid_pin_14_ cbx_6__7_/bottom_grid_pin_15_
+ cbx_6__7_/bottom_grid_pin_1_ cbx_6__7_/bottom_grid_pin_2_ cbx_6__7_/REGOUT_FEEDTHROUGH
+ grid_clb_6__7_/top_width_0_height_0__pin_33_ sb_6__7_/left_bottom_grid_pin_34_ sb_5__7_/right_bottom_grid_pin_34_
+ sb_6__7_/left_bottom_grid_pin_35_ sb_5__7_/right_bottom_grid_pin_35_ sb_6__7_/left_bottom_grid_pin_36_
+ sb_5__7_/right_bottom_grid_pin_36_ sb_6__7_/left_bottom_grid_pin_37_ sb_5__7_/right_bottom_grid_pin_37_
+ sb_6__7_/left_bottom_grid_pin_38_ sb_5__7_/right_bottom_grid_pin_38_ sb_6__7_/left_bottom_grid_pin_39_
+ sb_5__7_/right_bottom_grid_pin_39_ cbx_6__7_/bottom_grid_pin_3_ sb_6__7_/left_bottom_grid_pin_40_
+ sb_5__7_/right_bottom_grid_pin_40_ sb_6__7_/left_bottom_grid_pin_41_ sb_5__7_/right_bottom_grid_pin_41_
+ cbx_6__7_/bottom_grid_pin_4_ cbx_6__7_/bottom_grid_pin_5_ cbx_6__7_/bottom_grid_pin_6_
+ cbx_6__7_/bottom_grid_pin_7_ cbx_6__7_/bottom_grid_pin_8_ cbx_6__7_/bottom_grid_pin_9_
+ grid_clb
Xgrid_clb_3__4_ cbx_3__4_/SC_OUT_BOT cbx_3__3_/SC_IN_TOP grid_clb_3__4_/SC_OUT_TOP
+ cby_3__4_/Test_en_W_out grid_clb_3__4_/Test_en_E_out cby_3__4_/Test_en_W_out cby_2__4_/Test_en_W_in
+ VGND VPWR cbx_3__3_/REGIN_FEEDTHROUGH grid_clb_3__4_/bottom_width_0_height_0__pin_51_
+ cby_2__4_/ccff_tail cby_3__4_/ccff_head cbx_3__3_/clk_1_N_out cbx_3__3_/clk_1_N_out
+ cby_3__4_/prog_clk_0_W_in cbx_3__3_/prog_clk_1_N_out grid_clb_3__4_/prog_clk_0_N_out
+ cbx_3__3_/prog_clk_1_N_out cbx_3__3_/prog_clk_0_N_in grid_clb_3__4_/prog_clk_0_W_out
+ cby_3__4_/left_grid_pin_16_ cby_3__4_/left_grid_pin_17_ cby_3__4_/left_grid_pin_18_
+ cby_3__4_/left_grid_pin_19_ cby_3__4_/left_grid_pin_20_ cby_3__4_/left_grid_pin_21_
+ cby_3__4_/left_grid_pin_22_ cby_3__4_/left_grid_pin_23_ cby_3__4_/left_grid_pin_24_
+ cby_3__4_/left_grid_pin_25_ cby_3__4_/left_grid_pin_26_ cby_3__4_/left_grid_pin_27_
+ cby_3__4_/left_grid_pin_28_ cby_3__4_/left_grid_pin_29_ cby_3__4_/left_grid_pin_30_
+ cby_3__4_/left_grid_pin_31_ sb_3__3_/top_left_grid_pin_42_ sb_3__4_/bottom_left_grid_pin_42_
+ sb_3__3_/top_left_grid_pin_43_ sb_3__4_/bottom_left_grid_pin_43_ sb_3__3_/top_left_grid_pin_44_
+ sb_3__4_/bottom_left_grid_pin_44_ sb_3__3_/top_left_grid_pin_45_ sb_3__4_/bottom_left_grid_pin_45_
+ sb_3__3_/top_left_grid_pin_46_ sb_3__4_/bottom_left_grid_pin_46_ sb_3__3_/top_left_grid_pin_47_
+ sb_3__4_/bottom_left_grid_pin_47_ sb_3__3_/top_left_grid_pin_48_ sb_3__4_/bottom_left_grid_pin_48_
+ sb_3__3_/top_left_grid_pin_49_ sb_3__4_/bottom_left_grid_pin_49_ cbx_3__4_/bottom_grid_pin_0_
+ cbx_3__4_/bottom_grid_pin_10_ cbx_3__4_/bottom_grid_pin_11_ cbx_3__4_/bottom_grid_pin_12_
+ cbx_3__4_/bottom_grid_pin_13_ cbx_3__4_/bottom_grid_pin_14_ cbx_3__4_/bottom_grid_pin_15_
+ cbx_3__4_/bottom_grid_pin_1_ cbx_3__4_/bottom_grid_pin_2_ cbx_3__4_/REGOUT_FEEDTHROUGH
+ grid_clb_3__4_/top_width_0_height_0__pin_33_ sb_3__4_/left_bottom_grid_pin_34_ sb_2__4_/right_bottom_grid_pin_34_
+ sb_3__4_/left_bottom_grid_pin_35_ sb_2__4_/right_bottom_grid_pin_35_ sb_3__4_/left_bottom_grid_pin_36_
+ sb_2__4_/right_bottom_grid_pin_36_ sb_3__4_/left_bottom_grid_pin_37_ sb_2__4_/right_bottom_grid_pin_37_
+ sb_3__4_/left_bottom_grid_pin_38_ sb_2__4_/right_bottom_grid_pin_38_ sb_3__4_/left_bottom_grid_pin_39_
+ sb_2__4_/right_bottom_grid_pin_39_ cbx_3__4_/bottom_grid_pin_3_ sb_3__4_/left_bottom_grid_pin_40_
+ sb_2__4_/right_bottom_grid_pin_40_ sb_3__4_/left_bottom_grid_pin_41_ sb_2__4_/right_bottom_grid_pin_41_
+ cbx_3__4_/bottom_grid_pin_4_ cbx_3__4_/bottom_grid_pin_5_ cbx_3__4_/bottom_grid_pin_6_
+ cbx_3__4_/bottom_grid_pin_7_ cbx_3__4_/bottom_grid_pin_8_ cbx_3__4_/bottom_grid_pin_9_
+ grid_clb
Xcbx_1__1_ cbx_1__1_/REGIN_FEEDTHROUGH cbx_1__1_/REGOUT_FEEDTHROUGH cbx_1__1_/SC_IN_BOT
+ cbx_1__1_/SC_IN_TOP cbx_1__1_/SC_OUT_BOT cbx_1__1_/SC_OUT_TOP VGND VPWR cbx_1__1_/bottom_grid_pin_0_
+ cbx_1__1_/bottom_grid_pin_10_ cbx_1__1_/bottom_grid_pin_11_ cbx_1__1_/bottom_grid_pin_12_
+ cbx_1__1_/bottom_grid_pin_13_ cbx_1__1_/bottom_grid_pin_14_ cbx_1__1_/bottom_grid_pin_15_
+ cbx_1__1_/bottom_grid_pin_1_ cbx_1__1_/bottom_grid_pin_2_ cbx_1__1_/bottom_grid_pin_3_
+ cbx_1__1_/bottom_grid_pin_4_ cbx_1__1_/bottom_grid_pin_5_ cbx_1__1_/bottom_grid_pin_6_
+ cbx_1__1_/bottom_grid_pin_7_ cbx_1__1_/bottom_grid_pin_8_ cbx_1__1_/bottom_grid_pin_9_
+ sb_1__1_/ccff_tail sb_0__1_/ccff_head cbx_1__1_/chanx_left_in[0] cbx_1__1_/chanx_left_in[10]
+ cbx_1__1_/chanx_left_in[11] cbx_1__1_/chanx_left_in[12] cbx_1__1_/chanx_left_in[13]
+ cbx_1__1_/chanx_left_in[14] cbx_1__1_/chanx_left_in[15] cbx_1__1_/chanx_left_in[16]
+ cbx_1__1_/chanx_left_in[17] cbx_1__1_/chanx_left_in[18] cbx_1__1_/chanx_left_in[19]
+ cbx_1__1_/chanx_left_in[1] cbx_1__1_/chanx_left_in[2] cbx_1__1_/chanx_left_in[3]
+ cbx_1__1_/chanx_left_in[4] cbx_1__1_/chanx_left_in[5] cbx_1__1_/chanx_left_in[6]
+ cbx_1__1_/chanx_left_in[7] cbx_1__1_/chanx_left_in[8] cbx_1__1_/chanx_left_in[9]
+ sb_0__1_/chanx_right_in[0] sb_0__1_/chanx_right_in[10] sb_0__1_/chanx_right_in[11]
+ sb_0__1_/chanx_right_in[12] sb_0__1_/chanx_right_in[13] sb_0__1_/chanx_right_in[14]
+ sb_0__1_/chanx_right_in[15] sb_0__1_/chanx_right_in[16] sb_0__1_/chanx_right_in[17]
+ sb_0__1_/chanx_right_in[18] sb_0__1_/chanx_right_in[19] sb_0__1_/chanx_right_in[1]
+ sb_0__1_/chanx_right_in[2] sb_0__1_/chanx_right_in[3] sb_0__1_/chanx_right_in[4]
+ sb_0__1_/chanx_right_in[5] sb_0__1_/chanx_right_in[6] sb_0__1_/chanx_right_in[7]
+ sb_0__1_/chanx_right_in[8] sb_0__1_/chanx_right_in[9] sb_1__1_/chanx_left_out[0]
+ sb_1__1_/chanx_left_out[10] sb_1__1_/chanx_left_out[11] sb_1__1_/chanx_left_out[12]
+ sb_1__1_/chanx_left_out[13] sb_1__1_/chanx_left_out[14] sb_1__1_/chanx_left_out[15]
+ sb_1__1_/chanx_left_out[16] sb_1__1_/chanx_left_out[17] sb_1__1_/chanx_left_out[18]
+ sb_1__1_/chanx_left_out[19] sb_1__1_/chanx_left_out[1] sb_1__1_/chanx_left_out[2]
+ sb_1__1_/chanx_left_out[3] sb_1__1_/chanx_left_out[4] sb_1__1_/chanx_left_out[5]
+ sb_1__1_/chanx_left_out[6] sb_1__1_/chanx_left_out[7] sb_1__1_/chanx_left_out[8]
+ sb_1__1_/chanx_left_out[9] sb_1__1_/chanx_left_in[0] sb_1__1_/chanx_left_in[10]
+ sb_1__1_/chanx_left_in[11] sb_1__1_/chanx_left_in[12] sb_1__1_/chanx_left_in[13]
+ sb_1__1_/chanx_left_in[14] sb_1__1_/chanx_left_in[15] sb_1__1_/chanx_left_in[16]
+ sb_1__1_/chanx_left_in[17] sb_1__1_/chanx_left_in[18] sb_1__1_/chanx_left_in[19]
+ sb_1__1_/chanx_left_in[1] sb_1__1_/chanx_left_in[2] sb_1__1_/chanx_left_in[3] sb_1__1_/chanx_left_in[4]
+ sb_1__1_/chanx_left_in[5] sb_1__1_/chanx_left_in[6] sb_1__1_/chanx_left_in[7] sb_1__1_/chanx_left_in[8]
+ sb_1__1_/chanx_left_in[9] cbx_1__1_/clk_1_N_out cbx_1__1_/clk_1_S_out sb_1__1_/clk_1_W_out
+ cbx_1__1_/clk_2_E_out cbx_1__1_/clk_2_W_in cbx_1__1_/clk_2_W_out cbx_1__1_/clk_3_E_out
+ cbx_1__1_/clk_3_W_in cbx_1__1_/clk_3_W_out cbx_1__1_/prog_clk_0_N_in sb_0__1_/prog_clk_0_E_in
+ cbx_1__1_/prog_clk_1_N_out cbx_1__1_/prog_clk_1_S_out sb_1__1_/prog_clk_1_W_out
+ cbx_1__1_/prog_clk_2_E_out cbx_1__1_/prog_clk_2_W_in cbx_1__1_/prog_clk_2_W_out
+ cbx_1__1_/prog_clk_3_E_out cbx_1__1_/prog_clk_3_W_in cbx_1__1_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_8__1_ VGND VPWR sb_8__1_/bottom_left_grid_pin_42_ sb_8__1_/bottom_left_grid_pin_43_
+ sb_8__1_/bottom_left_grid_pin_44_ sb_8__1_/bottom_left_grid_pin_45_ sb_8__1_/bottom_left_grid_pin_46_
+ sb_8__1_/bottom_left_grid_pin_47_ sb_8__1_/bottom_left_grid_pin_48_ sb_8__1_/bottom_left_grid_pin_49_
+ sb_8__1_/bottom_right_grid_pin_1_ sb_8__1_/ccff_head sb_8__1_/ccff_tail sb_8__1_/chanx_left_in[0]
+ sb_8__1_/chanx_left_in[10] sb_8__1_/chanx_left_in[11] sb_8__1_/chanx_left_in[12]
+ sb_8__1_/chanx_left_in[13] sb_8__1_/chanx_left_in[14] sb_8__1_/chanx_left_in[15]
+ sb_8__1_/chanx_left_in[16] sb_8__1_/chanx_left_in[17] sb_8__1_/chanx_left_in[18]
+ sb_8__1_/chanx_left_in[19] sb_8__1_/chanx_left_in[1] sb_8__1_/chanx_left_in[2] sb_8__1_/chanx_left_in[3]
+ sb_8__1_/chanx_left_in[4] sb_8__1_/chanx_left_in[5] sb_8__1_/chanx_left_in[6] sb_8__1_/chanx_left_in[7]
+ sb_8__1_/chanx_left_in[8] sb_8__1_/chanx_left_in[9] sb_8__1_/chanx_left_out[0] sb_8__1_/chanx_left_out[10]
+ sb_8__1_/chanx_left_out[11] sb_8__1_/chanx_left_out[12] sb_8__1_/chanx_left_out[13]
+ sb_8__1_/chanx_left_out[14] sb_8__1_/chanx_left_out[15] sb_8__1_/chanx_left_out[16]
+ sb_8__1_/chanx_left_out[17] sb_8__1_/chanx_left_out[18] sb_8__1_/chanx_left_out[19]
+ sb_8__1_/chanx_left_out[1] sb_8__1_/chanx_left_out[2] sb_8__1_/chanx_left_out[3]
+ sb_8__1_/chanx_left_out[4] sb_8__1_/chanx_left_out[5] sb_8__1_/chanx_left_out[6]
+ sb_8__1_/chanx_left_out[7] sb_8__1_/chanx_left_out[8] sb_8__1_/chanx_left_out[9]
+ cby_8__1_/chany_top_out[0] cby_8__1_/chany_top_out[10] cby_8__1_/chany_top_out[11]
+ cby_8__1_/chany_top_out[12] cby_8__1_/chany_top_out[13] cby_8__1_/chany_top_out[14]
+ cby_8__1_/chany_top_out[15] cby_8__1_/chany_top_out[16] cby_8__1_/chany_top_out[17]
+ cby_8__1_/chany_top_out[18] cby_8__1_/chany_top_out[19] cby_8__1_/chany_top_out[1]
+ cby_8__1_/chany_top_out[2] cby_8__1_/chany_top_out[3] cby_8__1_/chany_top_out[4]
+ cby_8__1_/chany_top_out[5] cby_8__1_/chany_top_out[6] cby_8__1_/chany_top_out[7]
+ cby_8__1_/chany_top_out[8] cby_8__1_/chany_top_out[9] cby_8__1_/chany_top_in[0]
+ cby_8__1_/chany_top_in[10] cby_8__1_/chany_top_in[11] cby_8__1_/chany_top_in[12]
+ cby_8__1_/chany_top_in[13] cby_8__1_/chany_top_in[14] cby_8__1_/chany_top_in[15]
+ cby_8__1_/chany_top_in[16] cby_8__1_/chany_top_in[17] cby_8__1_/chany_top_in[18]
+ cby_8__1_/chany_top_in[19] cby_8__1_/chany_top_in[1] cby_8__1_/chany_top_in[2] cby_8__1_/chany_top_in[3]
+ cby_8__1_/chany_top_in[4] cby_8__1_/chany_top_in[5] cby_8__1_/chany_top_in[6] cby_8__1_/chany_top_in[7]
+ cby_8__1_/chany_top_in[8] cby_8__1_/chany_top_in[9] sb_8__1_/chany_top_in[0] sb_8__1_/chany_top_in[10]
+ sb_8__1_/chany_top_in[11] sb_8__1_/chany_top_in[12] sb_8__1_/chany_top_in[13] sb_8__1_/chany_top_in[14]
+ sb_8__1_/chany_top_in[15] sb_8__1_/chany_top_in[16] sb_8__1_/chany_top_in[17] sb_8__1_/chany_top_in[18]
+ sb_8__1_/chany_top_in[19] sb_8__1_/chany_top_in[1] sb_8__1_/chany_top_in[2] sb_8__1_/chany_top_in[3]
+ sb_8__1_/chany_top_in[4] sb_8__1_/chany_top_in[5] sb_8__1_/chany_top_in[6] sb_8__1_/chany_top_in[7]
+ sb_8__1_/chany_top_in[8] sb_8__1_/chany_top_in[9] sb_8__1_/chany_top_out[0] sb_8__1_/chany_top_out[10]
+ sb_8__1_/chany_top_out[11] sb_8__1_/chany_top_out[12] sb_8__1_/chany_top_out[13]
+ sb_8__1_/chany_top_out[14] sb_8__1_/chany_top_out[15] sb_8__1_/chany_top_out[16]
+ sb_8__1_/chany_top_out[17] sb_8__1_/chany_top_out[18] sb_8__1_/chany_top_out[19]
+ sb_8__1_/chany_top_out[1] sb_8__1_/chany_top_out[2] sb_8__1_/chany_top_out[3] sb_8__1_/chany_top_out[4]
+ sb_8__1_/chany_top_out[5] sb_8__1_/chany_top_out[6] sb_8__1_/chany_top_out[7] sb_8__1_/chany_top_out[8]
+ sb_8__1_/chany_top_out[9] sb_8__1_/left_bottom_grid_pin_34_ sb_8__1_/left_bottom_grid_pin_35_
+ sb_8__1_/left_bottom_grid_pin_36_ sb_8__1_/left_bottom_grid_pin_37_ sb_8__1_/left_bottom_grid_pin_38_
+ sb_8__1_/left_bottom_grid_pin_39_ sb_8__1_/left_bottom_grid_pin_40_ sb_8__1_/left_bottom_grid_pin_41_
+ sb_8__1_/prog_clk_0_N_in sb_8__1_/top_left_grid_pin_42_ sb_8__1_/top_left_grid_pin_43_
+ sb_8__1_/top_left_grid_pin_44_ sb_8__1_/top_left_grid_pin_45_ sb_8__1_/top_left_grid_pin_46_
+ sb_8__1_/top_left_grid_pin_47_ sb_8__1_/top_left_grid_pin_48_ sb_8__1_/top_left_grid_pin_49_
+ sb_8__1_/top_right_grid_pin_1_ sb_2__1_
Xsb_1__6_ sb_1__6_/Test_en_N_out sb_1__6_/Test_en_S_in VGND VPWR sb_1__6_/bottom_left_grid_pin_42_
+ sb_1__6_/bottom_left_grid_pin_43_ sb_1__6_/bottom_left_grid_pin_44_ sb_1__6_/bottom_left_grid_pin_45_
+ sb_1__6_/bottom_left_grid_pin_46_ sb_1__6_/bottom_left_grid_pin_47_ sb_1__6_/bottom_left_grid_pin_48_
+ sb_1__6_/bottom_left_grid_pin_49_ sb_1__6_/ccff_head sb_1__6_/ccff_tail sb_1__6_/chanx_left_in[0]
+ sb_1__6_/chanx_left_in[10] sb_1__6_/chanx_left_in[11] sb_1__6_/chanx_left_in[12]
+ sb_1__6_/chanx_left_in[13] sb_1__6_/chanx_left_in[14] sb_1__6_/chanx_left_in[15]
+ sb_1__6_/chanx_left_in[16] sb_1__6_/chanx_left_in[17] sb_1__6_/chanx_left_in[18]
+ sb_1__6_/chanx_left_in[19] sb_1__6_/chanx_left_in[1] sb_1__6_/chanx_left_in[2] sb_1__6_/chanx_left_in[3]
+ sb_1__6_/chanx_left_in[4] sb_1__6_/chanx_left_in[5] sb_1__6_/chanx_left_in[6] sb_1__6_/chanx_left_in[7]
+ sb_1__6_/chanx_left_in[8] sb_1__6_/chanx_left_in[9] sb_1__6_/chanx_left_out[0] sb_1__6_/chanx_left_out[10]
+ sb_1__6_/chanx_left_out[11] sb_1__6_/chanx_left_out[12] sb_1__6_/chanx_left_out[13]
+ sb_1__6_/chanx_left_out[14] sb_1__6_/chanx_left_out[15] sb_1__6_/chanx_left_out[16]
+ sb_1__6_/chanx_left_out[17] sb_1__6_/chanx_left_out[18] sb_1__6_/chanx_left_out[19]
+ sb_1__6_/chanx_left_out[1] sb_1__6_/chanx_left_out[2] sb_1__6_/chanx_left_out[3]
+ sb_1__6_/chanx_left_out[4] sb_1__6_/chanx_left_out[5] sb_1__6_/chanx_left_out[6]
+ sb_1__6_/chanx_left_out[7] sb_1__6_/chanx_left_out[8] sb_1__6_/chanx_left_out[9]
+ sb_1__6_/chanx_right_in[0] sb_1__6_/chanx_right_in[10] sb_1__6_/chanx_right_in[11]
+ sb_1__6_/chanx_right_in[12] sb_1__6_/chanx_right_in[13] sb_1__6_/chanx_right_in[14]
+ sb_1__6_/chanx_right_in[15] sb_1__6_/chanx_right_in[16] sb_1__6_/chanx_right_in[17]
+ sb_1__6_/chanx_right_in[18] sb_1__6_/chanx_right_in[19] sb_1__6_/chanx_right_in[1]
+ sb_1__6_/chanx_right_in[2] sb_1__6_/chanx_right_in[3] sb_1__6_/chanx_right_in[4]
+ sb_1__6_/chanx_right_in[5] sb_1__6_/chanx_right_in[6] sb_1__6_/chanx_right_in[7]
+ sb_1__6_/chanx_right_in[8] sb_1__6_/chanx_right_in[9] cbx_2__6_/chanx_left_in[0]
+ cbx_2__6_/chanx_left_in[10] cbx_2__6_/chanx_left_in[11] cbx_2__6_/chanx_left_in[12]
+ cbx_2__6_/chanx_left_in[13] cbx_2__6_/chanx_left_in[14] cbx_2__6_/chanx_left_in[15]
+ cbx_2__6_/chanx_left_in[16] cbx_2__6_/chanx_left_in[17] cbx_2__6_/chanx_left_in[18]
+ cbx_2__6_/chanx_left_in[19] cbx_2__6_/chanx_left_in[1] cbx_2__6_/chanx_left_in[2]
+ cbx_2__6_/chanx_left_in[3] cbx_2__6_/chanx_left_in[4] cbx_2__6_/chanx_left_in[5]
+ cbx_2__6_/chanx_left_in[6] cbx_2__6_/chanx_left_in[7] cbx_2__6_/chanx_left_in[8]
+ cbx_2__6_/chanx_left_in[9] cby_1__6_/chany_top_out[0] cby_1__6_/chany_top_out[10]
+ cby_1__6_/chany_top_out[11] cby_1__6_/chany_top_out[12] cby_1__6_/chany_top_out[13]
+ cby_1__6_/chany_top_out[14] cby_1__6_/chany_top_out[15] cby_1__6_/chany_top_out[16]
+ cby_1__6_/chany_top_out[17] cby_1__6_/chany_top_out[18] cby_1__6_/chany_top_out[19]
+ cby_1__6_/chany_top_out[1] cby_1__6_/chany_top_out[2] cby_1__6_/chany_top_out[3]
+ cby_1__6_/chany_top_out[4] cby_1__6_/chany_top_out[5] cby_1__6_/chany_top_out[6]
+ cby_1__6_/chany_top_out[7] cby_1__6_/chany_top_out[8] cby_1__6_/chany_top_out[9]
+ cby_1__6_/chany_top_in[0] cby_1__6_/chany_top_in[10] cby_1__6_/chany_top_in[11]
+ cby_1__6_/chany_top_in[12] cby_1__6_/chany_top_in[13] cby_1__6_/chany_top_in[14]
+ cby_1__6_/chany_top_in[15] cby_1__6_/chany_top_in[16] cby_1__6_/chany_top_in[17]
+ cby_1__6_/chany_top_in[18] cby_1__6_/chany_top_in[19] cby_1__6_/chany_top_in[1]
+ cby_1__6_/chany_top_in[2] cby_1__6_/chany_top_in[3] cby_1__6_/chany_top_in[4] cby_1__6_/chany_top_in[5]
+ cby_1__6_/chany_top_in[6] cby_1__6_/chany_top_in[7] cby_1__6_/chany_top_in[8] cby_1__6_/chany_top_in[9]
+ sb_1__6_/chany_top_in[0] sb_1__6_/chany_top_in[10] sb_1__6_/chany_top_in[11] sb_1__6_/chany_top_in[12]
+ sb_1__6_/chany_top_in[13] sb_1__6_/chany_top_in[14] sb_1__6_/chany_top_in[15] sb_1__6_/chany_top_in[16]
+ sb_1__6_/chany_top_in[17] sb_1__6_/chany_top_in[18] sb_1__6_/chany_top_in[19] sb_1__6_/chany_top_in[1]
+ sb_1__6_/chany_top_in[2] sb_1__6_/chany_top_in[3] sb_1__6_/chany_top_in[4] sb_1__6_/chany_top_in[5]
+ sb_1__6_/chany_top_in[6] sb_1__6_/chany_top_in[7] sb_1__6_/chany_top_in[8] sb_1__6_/chany_top_in[9]
+ sb_1__6_/chany_top_out[0] sb_1__6_/chany_top_out[10] sb_1__6_/chany_top_out[11]
+ sb_1__6_/chany_top_out[12] sb_1__6_/chany_top_out[13] sb_1__6_/chany_top_out[14]
+ sb_1__6_/chany_top_out[15] sb_1__6_/chany_top_out[16] sb_1__6_/chany_top_out[17]
+ sb_1__6_/chany_top_out[18] sb_1__6_/chany_top_out[19] sb_1__6_/chany_top_out[1]
+ sb_1__6_/chany_top_out[2] sb_1__6_/chany_top_out[3] sb_1__6_/chany_top_out[4] sb_1__6_/chany_top_out[5]
+ sb_1__6_/chany_top_out[6] sb_1__6_/chany_top_out[7] sb_1__6_/chany_top_out[8] sb_1__6_/chany_top_out[9]
+ sb_1__6_/clk_1_E_out sb_1__6_/clk_1_N_in sb_1__6_/clk_1_W_out sb_1__6_/clk_2_E_out
+ sb_1__6_/clk_2_N_in sb_1__6_/clk_2_N_out sb_1__6_/clk_2_S_out sb_1__6_/clk_2_W_out
+ sb_1__6_/clk_3_E_out sb_1__6_/clk_3_N_in sb_1__6_/clk_3_N_out sb_1__6_/clk_3_S_out
+ sb_1__6_/clk_3_W_out sb_1__6_/left_bottom_grid_pin_34_ sb_1__6_/left_bottom_grid_pin_35_
+ sb_1__6_/left_bottom_grid_pin_36_ sb_1__6_/left_bottom_grid_pin_37_ sb_1__6_/left_bottom_grid_pin_38_
+ sb_1__6_/left_bottom_grid_pin_39_ sb_1__6_/left_bottom_grid_pin_40_ sb_1__6_/left_bottom_grid_pin_41_
+ sb_1__6_/prog_clk_0_N_in sb_1__6_/prog_clk_1_E_out sb_1__6_/prog_clk_1_N_in sb_1__6_/prog_clk_1_W_out
+ sb_1__6_/prog_clk_2_E_out sb_1__6_/prog_clk_2_N_in sb_1__6_/prog_clk_2_N_out sb_1__6_/prog_clk_2_S_out
+ sb_1__6_/prog_clk_2_W_out sb_1__6_/prog_clk_3_E_out sb_1__6_/prog_clk_3_N_in sb_1__6_/prog_clk_3_N_out
+ sb_1__6_/prog_clk_3_S_out sb_1__6_/prog_clk_3_W_out sb_1__6_/right_bottom_grid_pin_34_
+ sb_1__6_/right_bottom_grid_pin_35_ sb_1__6_/right_bottom_grid_pin_36_ sb_1__6_/right_bottom_grid_pin_37_
+ sb_1__6_/right_bottom_grid_pin_38_ sb_1__6_/right_bottom_grid_pin_39_ sb_1__6_/right_bottom_grid_pin_40_
+ sb_1__6_/right_bottom_grid_pin_41_ sb_1__6_/top_left_grid_pin_42_ sb_1__6_/top_left_grid_pin_43_
+ sb_1__6_/top_left_grid_pin_44_ sb_1__6_/top_left_grid_pin_45_ sb_1__6_/top_left_grid_pin_46_
+ sb_1__6_/top_left_grid_pin_47_ sb_1__6_/top_left_grid_pin_48_ sb_1__6_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_7__5_ cby_7__5_/Test_en_W_in cby_7__5_/Test_en_E_out cby_7__5_/Test_en_N_out
+ cby_7__5_/Test_en_W_in cby_7__5_/Test_en_W_in cby_7__5_/Test_en_W_out VGND VPWR
+ cby_7__5_/ccff_head cby_7__5_/ccff_tail sb_7__4_/chany_top_out[0] sb_7__4_/chany_top_out[10]
+ sb_7__4_/chany_top_out[11] sb_7__4_/chany_top_out[12] sb_7__4_/chany_top_out[13]
+ sb_7__4_/chany_top_out[14] sb_7__4_/chany_top_out[15] sb_7__4_/chany_top_out[16]
+ sb_7__4_/chany_top_out[17] sb_7__4_/chany_top_out[18] sb_7__4_/chany_top_out[19]
+ sb_7__4_/chany_top_out[1] sb_7__4_/chany_top_out[2] sb_7__4_/chany_top_out[3] sb_7__4_/chany_top_out[4]
+ sb_7__4_/chany_top_out[5] sb_7__4_/chany_top_out[6] sb_7__4_/chany_top_out[7] sb_7__4_/chany_top_out[8]
+ sb_7__4_/chany_top_out[9] sb_7__4_/chany_top_in[0] sb_7__4_/chany_top_in[10] sb_7__4_/chany_top_in[11]
+ sb_7__4_/chany_top_in[12] sb_7__4_/chany_top_in[13] sb_7__4_/chany_top_in[14] sb_7__4_/chany_top_in[15]
+ sb_7__4_/chany_top_in[16] sb_7__4_/chany_top_in[17] sb_7__4_/chany_top_in[18] sb_7__4_/chany_top_in[19]
+ sb_7__4_/chany_top_in[1] sb_7__4_/chany_top_in[2] sb_7__4_/chany_top_in[3] sb_7__4_/chany_top_in[4]
+ sb_7__4_/chany_top_in[5] sb_7__4_/chany_top_in[6] sb_7__4_/chany_top_in[7] sb_7__4_/chany_top_in[8]
+ sb_7__4_/chany_top_in[9] cby_7__5_/chany_top_in[0] cby_7__5_/chany_top_in[10] cby_7__5_/chany_top_in[11]
+ cby_7__5_/chany_top_in[12] cby_7__5_/chany_top_in[13] cby_7__5_/chany_top_in[14]
+ cby_7__5_/chany_top_in[15] cby_7__5_/chany_top_in[16] cby_7__5_/chany_top_in[17]
+ cby_7__5_/chany_top_in[18] cby_7__5_/chany_top_in[19] cby_7__5_/chany_top_in[1]
+ cby_7__5_/chany_top_in[2] cby_7__5_/chany_top_in[3] cby_7__5_/chany_top_in[4] cby_7__5_/chany_top_in[5]
+ cby_7__5_/chany_top_in[6] cby_7__5_/chany_top_in[7] cby_7__5_/chany_top_in[8] cby_7__5_/chany_top_in[9]
+ cby_7__5_/chany_top_out[0] cby_7__5_/chany_top_out[10] cby_7__5_/chany_top_out[11]
+ cby_7__5_/chany_top_out[12] cby_7__5_/chany_top_out[13] cby_7__5_/chany_top_out[14]
+ cby_7__5_/chany_top_out[15] cby_7__5_/chany_top_out[16] cby_7__5_/chany_top_out[17]
+ cby_7__5_/chany_top_out[18] cby_7__5_/chany_top_out[19] cby_7__5_/chany_top_out[1]
+ cby_7__5_/chany_top_out[2] cby_7__5_/chany_top_out[3] cby_7__5_/chany_top_out[4]
+ cby_7__5_/chany_top_out[5] cby_7__5_/chany_top_out[6] cby_7__5_/chany_top_out[7]
+ cby_7__5_/chany_top_out[8] cby_7__5_/chany_top_out[9] cby_7__5_/clk_2_N_out cby_7__5_/clk_2_S_in
+ cby_7__5_/clk_2_S_out cby_7__5_/clk_3_N_out cby_7__5_/clk_3_S_in cby_7__5_/clk_3_S_out
+ cby_7__5_/left_grid_pin_16_ cby_7__5_/left_grid_pin_17_ cby_7__5_/left_grid_pin_18_
+ cby_7__5_/left_grid_pin_19_ cby_7__5_/left_grid_pin_20_ cby_7__5_/left_grid_pin_21_
+ cby_7__5_/left_grid_pin_22_ cby_7__5_/left_grid_pin_23_ cby_7__5_/left_grid_pin_24_
+ cby_7__5_/left_grid_pin_25_ cby_7__5_/left_grid_pin_26_ cby_7__5_/left_grid_pin_27_
+ cby_7__5_/left_grid_pin_28_ cby_7__5_/left_grid_pin_29_ cby_7__5_/left_grid_pin_30_
+ cby_7__5_/left_grid_pin_31_ cby_7__5_/prog_clk_0_N_out sb_7__4_/prog_clk_0_N_in
+ cby_7__5_/prog_clk_0_W_in cby_7__5_/prog_clk_2_N_out cby_7__5_/prog_clk_2_S_in cby_7__5_/prog_clk_2_S_out
+ cby_7__5_/prog_clk_3_N_out cby_7__5_/prog_clk_3_S_in cby_7__5_/prog_clk_3_S_out
+ cby_1__1_
Xcby_4__2_ sb_4__1_/Test_en_N_out cby_4__2_/Test_en_E_out sb_4__2_/Test_en_S_in sb_4__1_/Test_en_N_out
+ sb_4__1_/Test_en_N_out cby_4__2_/Test_en_W_out VGND VPWR cby_4__2_/ccff_head cby_4__2_/ccff_tail
+ sb_4__1_/chany_top_out[0] sb_4__1_/chany_top_out[10] sb_4__1_/chany_top_out[11]
+ sb_4__1_/chany_top_out[12] sb_4__1_/chany_top_out[13] sb_4__1_/chany_top_out[14]
+ sb_4__1_/chany_top_out[15] sb_4__1_/chany_top_out[16] sb_4__1_/chany_top_out[17]
+ sb_4__1_/chany_top_out[18] sb_4__1_/chany_top_out[19] sb_4__1_/chany_top_out[1]
+ sb_4__1_/chany_top_out[2] sb_4__1_/chany_top_out[3] sb_4__1_/chany_top_out[4] sb_4__1_/chany_top_out[5]
+ sb_4__1_/chany_top_out[6] sb_4__1_/chany_top_out[7] sb_4__1_/chany_top_out[8] sb_4__1_/chany_top_out[9]
+ sb_4__1_/chany_top_in[0] sb_4__1_/chany_top_in[10] sb_4__1_/chany_top_in[11] sb_4__1_/chany_top_in[12]
+ sb_4__1_/chany_top_in[13] sb_4__1_/chany_top_in[14] sb_4__1_/chany_top_in[15] sb_4__1_/chany_top_in[16]
+ sb_4__1_/chany_top_in[17] sb_4__1_/chany_top_in[18] sb_4__1_/chany_top_in[19] sb_4__1_/chany_top_in[1]
+ sb_4__1_/chany_top_in[2] sb_4__1_/chany_top_in[3] sb_4__1_/chany_top_in[4] sb_4__1_/chany_top_in[5]
+ sb_4__1_/chany_top_in[6] sb_4__1_/chany_top_in[7] sb_4__1_/chany_top_in[8] sb_4__1_/chany_top_in[9]
+ cby_4__2_/chany_top_in[0] cby_4__2_/chany_top_in[10] cby_4__2_/chany_top_in[11]
+ cby_4__2_/chany_top_in[12] cby_4__2_/chany_top_in[13] cby_4__2_/chany_top_in[14]
+ cby_4__2_/chany_top_in[15] cby_4__2_/chany_top_in[16] cby_4__2_/chany_top_in[17]
+ cby_4__2_/chany_top_in[18] cby_4__2_/chany_top_in[19] cby_4__2_/chany_top_in[1]
+ cby_4__2_/chany_top_in[2] cby_4__2_/chany_top_in[3] cby_4__2_/chany_top_in[4] cby_4__2_/chany_top_in[5]
+ cby_4__2_/chany_top_in[6] cby_4__2_/chany_top_in[7] cby_4__2_/chany_top_in[8] cby_4__2_/chany_top_in[9]
+ cby_4__2_/chany_top_out[0] cby_4__2_/chany_top_out[10] cby_4__2_/chany_top_out[11]
+ cby_4__2_/chany_top_out[12] cby_4__2_/chany_top_out[13] cby_4__2_/chany_top_out[14]
+ cby_4__2_/chany_top_out[15] cby_4__2_/chany_top_out[16] cby_4__2_/chany_top_out[17]
+ cby_4__2_/chany_top_out[18] cby_4__2_/chany_top_out[19] cby_4__2_/chany_top_out[1]
+ cby_4__2_/chany_top_out[2] cby_4__2_/chany_top_out[3] cby_4__2_/chany_top_out[4]
+ cby_4__2_/chany_top_out[5] cby_4__2_/chany_top_out[6] cby_4__2_/chany_top_out[7]
+ cby_4__2_/chany_top_out[8] cby_4__2_/chany_top_out[9] cby_4__2_/clk_2_N_out cby_4__2_/clk_2_S_in
+ cby_4__2_/clk_2_S_out sb_4__2_/clk_3_N_in sb_4__1_/clk_3_N_out cby_4__2_/clk_3_S_out
+ cby_4__2_/left_grid_pin_16_ cby_4__2_/left_grid_pin_17_ cby_4__2_/left_grid_pin_18_
+ cby_4__2_/left_grid_pin_19_ cby_4__2_/left_grid_pin_20_ cby_4__2_/left_grid_pin_21_
+ cby_4__2_/left_grid_pin_22_ cby_4__2_/left_grid_pin_23_ cby_4__2_/left_grid_pin_24_
+ cby_4__2_/left_grid_pin_25_ cby_4__2_/left_grid_pin_26_ cby_4__2_/left_grid_pin_27_
+ cby_4__2_/left_grid_pin_28_ cby_4__2_/left_grid_pin_29_ cby_4__2_/left_grid_pin_30_
+ cby_4__2_/left_grid_pin_31_ cby_4__2_/prog_clk_0_N_out sb_4__1_/prog_clk_0_N_in
+ cby_4__2_/prog_clk_0_W_in cby_4__2_/prog_clk_2_N_out cby_4__2_/prog_clk_2_S_in cby_4__2_/prog_clk_2_S_out
+ sb_4__2_/prog_clk_3_N_in sb_4__1_/prog_clk_3_N_out cby_4__2_/prog_clk_3_S_out cby_1__1_
Xcbx_7__6_ cbx_7__6_/REGIN_FEEDTHROUGH cbx_7__6_/REGOUT_FEEDTHROUGH cbx_7__6_/SC_IN_BOT
+ cbx_7__6_/SC_IN_TOP cbx_7__6_/SC_OUT_BOT cbx_7__6_/SC_OUT_TOP VGND VPWR cbx_7__6_/bottom_grid_pin_0_
+ cbx_7__6_/bottom_grid_pin_10_ cbx_7__6_/bottom_grid_pin_11_ cbx_7__6_/bottom_grid_pin_12_
+ cbx_7__6_/bottom_grid_pin_13_ cbx_7__6_/bottom_grid_pin_14_ cbx_7__6_/bottom_grid_pin_15_
+ cbx_7__6_/bottom_grid_pin_1_ cbx_7__6_/bottom_grid_pin_2_ cbx_7__6_/bottom_grid_pin_3_
+ cbx_7__6_/bottom_grid_pin_4_ cbx_7__6_/bottom_grid_pin_5_ cbx_7__6_/bottom_grid_pin_6_
+ cbx_7__6_/bottom_grid_pin_7_ cbx_7__6_/bottom_grid_pin_8_ cbx_7__6_/bottom_grid_pin_9_
+ sb_7__6_/ccff_tail sb_6__6_/ccff_head cbx_7__6_/chanx_left_in[0] cbx_7__6_/chanx_left_in[10]
+ cbx_7__6_/chanx_left_in[11] cbx_7__6_/chanx_left_in[12] cbx_7__6_/chanx_left_in[13]
+ cbx_7__6_/chanx_left_in[14] cbx_7__6_/chanx_left_in[15] cbx_7__6_/chanx_left_in[16]
+ cbx_7__6_/chanx_left_in[17] cbx_7__6_/chanx_left_in[18] cbx_7__6_/chanx_left_in[19]
+ cbx_7__6_/chanx_left_in[1] cbx_7__6_/chanx_left_in[2] cbx_7__6_/chanx_left_in[3]
+ cbx_7__6_/chanx_left_in[4] cbx_7__6_/chanx_left_in[5] cbx_7__6_/chanx_left_in[6]
+ cbx_7__6_/chanx_left_in[7] cbx_7__6_/chanx_left_in[8] cbx_7__6_/chanx_left_in[9]
+ sb_6__6_/chanx_right_in[0] sb_6__6_/chanx_right_in[10] sb_6__6_/chanx_right_in[11]
+ sb_6__6_/chanx_right_in[12] sb_6__6_/chanx_right_in[13] sb_6__6_/chanx_right_in[14]
+ sb_6__6_/chanx_right_in[15] sb_6__6_/chanx_right_in[16] sb_6__6_/chanx_right_in[17]
+ sb_6__6_/chanx_right_in[18] sb_6__6_/chanx_right_in[19] sb_6__6_/chanx_right_in[1]
+ sb_6__6_/chanx_right_in[2] sb_6__6_/chanx_right_in[3] sb_6__6_/chanx_right_in[4]
+ sb_6__6_/chanx_right_in[5] sb_6__6_/chanx_right_in[6] sb_6__6_/chanx_right_in[7]
+ sb_6__6_/chanx_right_in[8] sb_6__6_/chanx_right_in[9] sb_7__6_/chanx_left_out[0]
+ sb_7__6_/chanx_left_out[10] sb_7__6_/chanx_left_out[11] sb_7__6_/chanx_left_out[12]
+ sb_7__6_/chanx_left_out[13] sb_7__6_/chanx_left_out[14] sb_7__6_/chanx_left_out[15]
+ sb_7__6_/chanx_left_out[16] sb_7__6_/chanx_left_out[17] sb_7__6_/chanx_left_out[18]
+ sb_7__6_/chanx_left_out[19] sb_7__6_/chanx_left_out[1] sb_7__6_/chanx_left_out[2]
+ sb_7__6_/chanx_left_out[3] sb_7__6_/chanx_left_out[4] sb_7__6_/chanx_left_out[5]
+ sb_7__6_/chanx_left_out[6] sb_7__6_/chanx_left_out[7] sb_7__6_/chanx_left_out[8]
+ sb_7__6_/chanx_left_out[9] sb_7__6_/chanx_left_in[0] sb_7__6_/chanx_left_in[10]
+ sb_7__6_/chanx_left_in[11] sb_7__6_/chanx_left_in[12] sb_7__6_/chanx_left_in[13]
+ sb_7__6_/chanx_left_in[14] sb_7__6_/chanx_left_in[15] sb_7__6_/chanx_left_in[16]
+ sb_7__6_/chanx_left_in[17] sb_7__6_/chanx_left_in[18] sb_7__6_/chanx_left_in[19]
+ sb_7__6_/chanx_left_in[1] sb_7__6_/chanx_left_in[2] sb_7__6_/chanx_left_in[3] sb_7__6_/chanx_left_in[4]
+ sb_7__6_/chanx_left_in[5] sb_7__6_/chanx_left_in[6] sb_7__6_/chanx_left_in[7] sb_7__6_/chanx_left_in[8]
+ sb_7__6_/chanx_left_in[9] cbx_7__6_/clk_1_N_out cbx_7__6_/clk_1_S_out cbx_7__6_/clk_1_W_in
+ sb_7__6_/clk_2_N_in sb_6__6_/clk_2_E_out cbx_7__6_/clk_2_W_out cbx_7__6_/clk_3_E_out
+ cbx_7__6_/clk_3_W_in cbx_7__6_/clk_3_W_out cbx_7__6_/prog_clk_0_N_in cbx_7__6_/prog_clk_0_W_out
+ cbx_7__6_/prog_clk_1_N_out cbx_7__6_/prog_clk_1_S_out cbx_7__6_/prog_clk_1_W_in
+ sb_7__6_/prog_clk_2_N_in sb_6__6_/prog_clk_2_E_out cbx_7__6_/prog_clk_2_W_out cbx_7__6_/prog_clk_3_E_out
+ cbx_7__6_/prog_clk_3_W_in cbx_7__6_/prog_clk_3_W_out cbx_1__1_
Xgrid_clb_6__6_ cbx_6__5_/SC_OUT_TOP grid_clb_6__6_/SC_OUT_BOT cbx_6__6_/SC_IN_BOT
+ cby_5__6_/Test_en_E_out cby_6__6_/Test_en_W_in cby_5__6_/Test_en_E_out grid_clb_6__6_/Test_en_W_out
+ VGND VPWR cbx_6__5_/REGIN_FEEDTHROUGH grid_clb_6__6_/bottom_width_0_height_0__pin_51_
+ cby_5__6_/ccff_tail cby_6__6_/ccff_head cbx_6__5_/clk_1_N_out cbx_6__5_/clk_1_N_out
+ cby_6__6_/prog_clk_0_W_in cbx_6__5_/prog_clk_1_N_out grid_clb_6__6_/prog_clk_0_N_out
+ cbx_6__5_/prog_clk_1_N_out cbx_6__5_/prog_clk_0_N_in grid_clb_6__6_/prog_clk_0_W_out
+ cby_6__6_/left_grid_pin_16_ cby_6__6_/left_grid_pin_17_ cby_6__6_/left_grid_pin_18_
+ cby_6__6_/left_grid_pin_19_ cby_6__6_/left_grid_pin_20_ cby_6__6_/left_grid_pin_21_
+ cby_6__6_/left_grid_pin_22_ cby_6__6_/left_grid_pin_23_ cby_6__6_/left_grid_pin_24_
+ cby_6__6_/left_grid_pin_25_ cby_6__6_/left_grid_pin_26_ cby_6__6_/left_grid_pin_27_
+ cby_6__6_/left_grid_pin_28_ cby_6__6_/left_grid_pin_29_ cby_6__6_/left_grid_pin_30_
+ cby_6__6_/left_grid_pin_31_ sb_6__5_/top_left_grid_pin_42_ sb_6__6_/bottom_left_grid_pin_42_
+ sb_6__5_/top_left_grid_pin_43_ sb_6__6_/bottom_left_grid_pin_43_ sb_6__5_/top_left_grid_pin_44_
+ sb_6__6_/bottom_left_grid_pin_44_ sb_6__5_/top_left_grid_pin_45_ sb_6__6_/bottom_left_grid_pin_45_
+ sb_6__5_/top_left_grid_pin_46_ sb_6__6_/bottom_left_grid_pin_46_ sb_6__5_/top_left_grid_pin_47_
+ sb_6__6_/bottom_left_grid_pin_47_ sb_6__5_/top_left_grid_pin_48_ sb_6__6_/bottom_left_grid_pin_48_
+ sb_6__5_/top_left_grid_pin_49_ sb_6__6_/bottom_left_grid_pin_49_ cbx_6__6_/bottom_grid_pin_0_
+ cbx_6__6_/bottom_grid_pin_10_ cbx_6__6_/bottom_grid_pin_11_ cbx_6__6_/bottom_grid_pin_12_
+ cbx_6__6_/bottom_grid_pin_13_ cbx_6__6_/bottom_grid_pin_14_ cbx_6__6_/bottom_grid_pin_15_
+ cbx_6__6_/bottom_grid_pin_1_ cbx_6__6_/bottom_grid_pin_2_ cbx_6__6_/REGOUT_FEEDTHROUGH
+ grid_clb_6__6_/top_width_0_height_0__pin_33_ sb_6__6_/left_bottom_grid_pin_34_ sb_5__6_/right_bottom_grid_pin_34_
+ sb_6__6_/left_bottom_grid_pin_35_ sb_5__6_/right_bottom_grid_pin_35_ sb_6__6_/left_bottom_grid_pin_36_
+ sb_5__6_/right_bottom_grid_pin_36_ sb_6__6_/left_bottom_grid_pin_37_ sb_5__6_/right_bottom_grid_pin_37_
+ sb_6__6_/left_bottom_grid_pin_38_ sb_5__6_/right_bottom_grid_pin_38_ sb_6__6_/left_bottom_grid_pin_39_
+ sb_5__6_/right_bottom_grid_pin_39_ cbx_6__6_/bottom_grid_pin_3_ sb_6__6_/left_bottom_grid_pin_40_
+ sb_5__6_/right_bottom_grid_pin_40_ sb_6__6_/left_bottom_grid_pin_41_ sb_5__6_/right_bottom_grid_pin_41_
+ cbx_6__6_/bottom_grid_pin_4_ cbx_6__6_/bottom_grid_pin_5_ cbx_6__6_/bottom_grid_pin_6_
+ cbx_6__6_/bottom_grid_pin_7_ cbx_6__6_/bottom_grid_pin_8_ cbx_6__6_/bottom_grid_pin_9_
+ grid_clb
Xcbx_4__3_ cbx_4__3_/REGIN_FEEDTHROUGH cbx_4__3_/REGOUT_FEEDTHROUGH cbx_4__3_/SC_IN_BOT
+ cbx_4__3_/SC_IN_TOP cbx_4__3_/SC_OUT_BOT cbx_4__3_/SC_OUT_TOP VGND VPWR cbx_4__3_/bottom_grid_pin_0_
+ cbx_4__3_/bottom_grid_pin_10_ cbx_4__3_/bottom_grid_pin_11_ cbx_4__3_/bottom_grid_pin_12_
+ cbx_4__3_/bottom_grid_pin_13_ cbx_4__3_/bottom_grid_pin_14_ cbx_4__3_/bottom_grid_pin_15_
+ cbx_4__3_/bottom_grid_pin_1_ cbx_4__3_/bottom_grid_pin_2_ cbx_4__3_/bottom_grid_pin_3_
+ cbx_4__3_/bottom_grid_pin_4_ cbx_4__3_/bottom_grid_pin_5_ cbx_4__3_/bottom_grid_pin_6_
+ cbx_4__3_/bottom_grid_pin_7_ cbx_4__3_/bottom_grid_pin_8_ cbx_4__3_/bottom_grid_pin_9_
+ sb_4__3_/ccff_tail sb_3__3_/ccff_head cbx_4__3_/chanx_left_in[0] cbx_4__3_/chanx_left_in[10]
+ cbx_4__3_/chanx_left_in[11] cbx_4__3_/chanx_left_in[12] cbx_4__3_/chanx_left_in[13]
+ cbx_4__3_/chanx_left_in[14] cbx_4__3_/chanx_left_in[15] cbx_4__3_/chanx_left_in[16]
+ cbx_4__3_/chanx_left_in[17] cbx_4__3_/chanx_left_in[18] cbx_4__3_/chanx_left_in[19]
+ cbx_4__3_/chanx_left_in[1] cbx_4__3_/chanx_left_in[2] cbx_4__3_/chanx_left_in[3]
+ cbx_4__3_/chanx_left_in[4] cbx_4__3_/chanx_left_in[5] cbx_4__3_/chanx_left_in[6]
+ cbx_4__3_/chanx_left_in[7] cbx_4__3_/chanx_left_in[8] cbx_4__3_/chanx_left_in[9]
+ sb_3__3_/chanx_right_in[0] sb_3__3_/chanx_right_in[10] sb_3__3_/chanx_right_in[11]
+ sb_3__3_/chanx_right_in[12] sb_3__3_/chanx_right_in[13] sb_3__3_/chanx_right_in[14]
+ sb_3__3_/chanx_right_in[15] sb_3__3_/chanx_right_in[16] sb_3__3_/chanx_right_in[17]
+ sb_3__3_/chanx_right_in[18] sb_3__3_/chanx_right_in[19] sb_3__3_/chanx_right_in[1]
+ sb_3__3_/chanx_right_in[2] sb_3__3_/chanx_right_in[3] sb_3__3_/chanx_right_in[4]
+ sb_3__3_/chanx_right_in[5] sb_3__3_/chanx_right_in[6] sb_3__3_/chanx_right_in[7]
+ sb_3__3_/chanx_right_in[8] sb_3__3_/chanx_right_in[9] sb_4__3_/chanx_left_out[0]
+ sb_4__3_/chanx_left_out[10] sb_4__3_/chanx_left_out[11] sb_4__3_/chanx_left_out[12]
+ sb_4__3_/chanx_left_out[13] sb_4__3_/chanx_left_out[14] sb_4__3_/chanx_left_out[15]
+ sb_4__3_/chanx_left_out[16] sb_4__3_/chanx_left_out[17] sb_4__3_/chanx_left_out[18]
+ sb_4__3_/chanx_left_out[19] sb_4__3_/chanx_left_out[1] sb_4__3_/chanx_left_out[2]
+ sb_4__3_/chanx_left_out[3] sb_4__3_/chanx_left_out[4] sb_4__3_/chanx_left_out[5]
+ sb_4__3_/chanx_left_out[6] sb_4__3_/chanx_left_out[7] sb_4__3_/chanx_left_out[8]
+ sb_4__3_/chanx_left_out[9] sb_4__3_/chanx_left_in[0] sb_4__3_/chanx_left_in[10]
+ sb_4__3_/chanx_left_in[11] sb_4__3_/chanx_left_in[12] sb_4__3_/chanx_left_in[13]
+ sb_4__3_/chanx_left_in[14] sb_4__3_/chanx_left_in[15] sb_4__3_/chanx_left_in[16]
+ sb_4__3_/chanx_left_in[17] sb_4__3_/chanx_left_in[18] sb_4__3_/chanx_left_in[19]
+ sb_4__3_/chanx_left_in[1] sb_4__3_/chanx_left_in[2] sb_4__3_/chanx_left_in[3] sb_4__3_/chanx_left_in[4]
+ sb_4__3_/chanx_left_in[5] sb_4__3_/chanx_left_in[6] sb_4__3_/chanx_left_in[7] sb_4__3_/chanx_left_in[8]
+ sb_4__3_/chanx_left_in[9] cbx_4__3_/clk_1_N_out cbx_4__3_/clk_1_S_out sb_3__3_/clk_1_E_out
+ cbx_4__3_/clk_2_E_out cbx_4__3_/clk_2_W_in cbx_4__3_/clk_2_W_out cbx_4__3_/clk_3_E_out
+ cbx_4__3_/clk_3_W_in cbx_4__3_/clk_3_W_out cbx_4__3_/prog_clk_0_N_in cbx_4__3_/prog_clk_0_W_out
+ cbx_4__3_/prog_clk_1_N_out cbx_4__3_/prog_clk_1_S_out sb_3__3_/prog_clk_1_E_out
+ cbx_4__3_/prog_clk_2_E_out cbx_4__3_/prog_clk_2_W_in cbx_4__3_/prog_clk_2_W_out
+ cbx_4__3_/prog_clk_3_E_out cbx_4__3_/prog_clk_3_W_in cbx_4__3_/prog_clk_3_W_out
+ cbx_1__1_
Xcbx_1__0_ IO_ISOL_N cbx_1__0_/SC_IN_BOT cbx_1__0_/SC_IN_TOP sb_1__0_/SC_IN_TOP cbx_1__0_/SC_OUT_TOP
+ VGND VPWR cbx_1__0_/bottom_grid_pin_0_ cbx_1__0_/bottom_grid_pin_10_ cbx_1__0_/bottom_grid_pin_12_
+ cbx_1__0_/bottom_grid_pin_14_ cbx_1__0_/bottom_grid_pin_16_ cbx_1__0_/bottom_grid_pin_2_
+ cbx_1__0_/bottom_grid_pin_4_ cbx_1__0_/bottom_grid_pin_6_ cbx_1__0_/bottom_grid_pin_8_
+ sb_1__0_/ccff_tail sb_0__0_/ccff_head cbx_1__0_/chanx_left_in[0] cbx_1__0_/chanx_left_in[10]
+ cbx_1__0_/chanx_left_in[11] cbx_1__0_/chanx_left_in[12] cbx_1__0_/chanx_left_in[13]
+ cbx_1__0_/chanx_left_in[14] cbx_1__0_/chanx_left_in[15] cbx_1__0_/chanx_left_in[16]
+ cbx_1__0_/chanx_left_in[17] cbx_1__0_/chanx_left_in[18] cbx_1__0_/chanx_left_in[19]
+ cbx_1__0_/chanx_left_in[1] cbx_1__0_/chanx_left_in[2] cbx_1__0_/chanx_left_in[3]
+ cbx_1__0_/chanx_left_in[4] cbx_1__0_/chanx_left_in[5] cbx_1__0_/chanx_left_in[6]
+ cbx_1__0_/chanx_left_in[7] cbx_1__0_/chanx_left_in[8] cbx_1__0_/chanx_left_in[9]
+ sb_0__0_/chanx_right_in[0] sb_0__0_/chanx_right_in[10] sb_0__0_/chanx_right_in[11]
+ sb_0__0_/chanx_right_in[12] sb_0__0_/chanx_right_in[13] sb_0__0_/chanx_right_in[14]
+ sb_0__0_/chanx_right_in[15] sb_0__0_/chanx_right_in[16] sb_0__0_/chanx_right_in[17]
+ sb_0__0_/chanx_right_in[18] sb_0__0_/chanx_right_in[19] sb_0__0_/chanx_right_in[1]
+ sb_0__0_/chanx_right_in[2] sb_0__0_/chanx_right_in[3] sb_0__0_/chanx_right_in[4]
+ sb_0__0_/chanx_right_in[5] sb_0__0_/chanx_right_in[6] sb_0__0_/chanx_right_in[7]
+ sb_0__0_/chanx_right_in[8] sb_0__0_/chanx_right_in[9] sb_1__0_/chanx_left_out[0]
+ sb_1__0_/chanx_left_out[10] sb_1__0_/chanx_left_out[11] sb_1__0_/chanx_left_out[12]
+ sb_1__0_/chanx_left_out[13] sb_1__0_/chanx_left_out[14] sb_1__0_/chanx_left_out[15]
+ sb_1__0_/chanx_left_out[16] sb_1__0_/chanx_left_out[17] sb_1__0_/chanx_left_out[18]
+ sb_1__0_/chanx_left_out[19] sb_1__0_/chanx_left_out[1] sb_1__0_/chanx_left_out[2]
+ sb_1__0_/chanx_left_out[3] sb_1__0_/chanx_left_out[4] sb_1__0_/chanx_left_out[5]
+ sb_1__0_/chanx_left_out[6] sb_1__0_/chanx_left_out[7] sb_1__0_/chanx_left_out[8]
+ sb_1__0_/chanx_left_out[9] sb_1__0_/chanx_left_in[0] sb_1__0_/chanx_left_in[10]
+ sb_1__0_/chanx_left_in[11] sb_1__0_/chanx_left_in[12] sb_1__0_/chanx_left_in[13]
+ sb_1__0_/chanx_left_in[14] sb_1__0_/chanx_left_in[15] sb_1__0_/chanx_left_in[16]
+ sb_1__0_/chanx_left_in[17] sb_1__0_/chanx_left_in[18] sb_1__0_/chanx_left_in[19]
+ sb_1__0_/chanx_left_in[1] sb_1__0_/chanx_left_in[2] sb_1__0_/chanx_left_in[3] sb_1__0_/chanx_left_in[4]
+ sb_1__0_/chanx_left_in[5] sb_1__0_/chanx_left_in[6] sb_1__0_/chanx_left_in[7] sb_1__0_/chanx_left_in[8]
+ sb_1__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87] cbx_1__0_/prog_clk_0_N_in sb_0__0_/prog_clk_0_E_in
+ cbx_1__0_/bottom_grid_pin_0_ cbx_1__0_/bottom_grid_pin_10_ sb_1__0_/left_bottom_grid_pin_11_
+ sb_0__0_/right_bottom_grid_pin_11_ cbx_1__0_/bottom_grid_pin_12_ sb_1__0_/left_bottom_grid_pin_13_
+ sb_0__0_/right_bottom_grid_pin_13_ cbx_1__0_/bottom_grid_pin_14_ sb_1__0_/left_bottom_grid_pin_15_
+ sb_0__0_/right_bottom_grid_pin_15_ cbx_1__0_/bottom_grid_pin_16_ sb_1__0_/left_bottom_grid_pin_17_
+ sb_0__0_/right_bottom_grid_pin_17_ sb_1__0_/left_bottom_grid_pin_1_ sb_0__0_/right_bottom_grid_pin_1_
+ cbx_1__0_/bottom_grid_pin_2_ sb_1__0_/left_bottom_grid_pin_3_ sb_0__0_/right_bottom_grid_pin_3_
+ cbx_1__0_/bottom_grid_pin_4_ sb_1__0_/left_bottom_grid_pin_5_ sb_0__0_/right_bottom_grid_pin_5_
+ cbx_1__0_/bottom_grid_pin_6_ sb_1__0_/left_bottom_grid_pin_7_ sb_0__0_/right_bottom_grid_pin_7_
+ cbx_1__0_/bottom_grid_pin_8_ sb_1__0_/left_bottom_grid_pin_9_ sb_0__0_/right_bottom_grid_pin_9_
+ cbx_1__0_
Xsb_8__0_ VGND VPWR sb_8__0_/ccff_head sb_8__0_/ccff_tail sb_8__0_/chanx_left_in[0]
+ sb_8__0_/chanx_left_in[10] sb_8__0_/chanx_left_in[11] sb_8__0_/chanx_left_in[12]
+ sb_8__0_/chanx_left_in[13] sb_8__0_/chanx_left_in[14] sb_8__0_/chanx_left_in[15]
+ sb_8__0_/chanx_left_in[16] sb_8__0_/chanx_left_in[17] sb_8__0_/chanx_left_in[18]
+ sb_8__0_/chanx_left_in[19] sb_8__0_/chanx_left_in[1] sb_8__0_/chanx_left_in[2] sb_8__0_/chanx_left_in[3]
+ sb_8__0_/chanx_left_in[4] sb_8__0_/chanx_left_in[5] sb_8__0_/chanx_left_in[6] sb_8__0_/chanx_left_in[7]
+ sb_8__0_/chanx_left_in[8] sb_8__0_/chanx_left_in[9] sb_8__0_/chanx_left_out[0] sb_8__0_/chanx_left_out[10]
+ sb_8__0_/chanx_left_out[11] sb_8__0_/chanx_left_out[12] sb_8__0_/chanx_left_out[13]
+ sb_8__0_/chanx_left_out[14] sb_8__0_/chanx_left_out[15] sb_8__0_/chanx_left_out[16]
+ sb_8__0_/chanx_left_out[17] sb_8__0_/chanx_left_out[18] sb_8__0_/chanx_left_out[19]
+ sb_8__0_/chanx_left_out[1] sb_8__0_/chanx_left_out[2] sb_8__0_/chanx_left_out[3]
+ sb_8__0_/chanx_left_out[4] sb_8__0_/chanx_left_out[5] sb_8__0_/chanx_left_out[6]
+ sb_8__0_/chanx_left_out[7] sb_8__0_/chanx_left_out[8] sb_8__0_/chanx_left_out[9]
+ sb_8__0_/chany_top_in[0] sb_8__0_/chany_top_in[10] sb_8__0_/chany_top_in[11] sb_8__0_/chany_top_in[12]
+ sb_8__0_/chany_top_in[13] sb_8__0_/chany_top_in[14] sb_8__0_/chany_top_in[15] sb_8__0_/chany_top_in[16]
+ sb_8__0_/chany_top_in[17] sb_8__0_/chany_top_in[18] sb_8__0_/chany_top_in[19] sb_8__0_/chany_top_in[1]
+ sb_8__0_/chany_top_in[2] sb_8__0_/chany_top_in[3] sb_8__0_/chany_top_in[4] sb_8__0_/chany_top_in[5]
+ sb_8__0_/chany_top_in[6] sb_8__0_/chany_top_in[7] sb_8__0_/chany_top_in[8] sb_8__0_/chany_top_in[9]
+ sb_8__0_/chany_top_out[0] sb_8__0_/chany_top_out[10] sb_8__0_/chany_top_out[11]
+ sb_8__0_/chany_top_out[12] sb_8__0_/chany_top_out[13] sb_8__0_/chany_top_out[14]
+ sb_8__0_/chany_top_out[15] sb_8__0_/chany_top_out[16] sb_8__0_/chany_top_out[17]
+ sb_8__0_/chany_top_out[18] sb_8__0_/chany_top_out[19] sb_8__0_/chany_top_out[1]
+ sb_8__0_/chany_top_out[2] sb_8__0_/chany_top_out[3] sb_8__0_/chany_top_out[4] sb_8__0_/chany_top_out[5]
+ sb_8__0_/chany_top_out[6] sb_8__0_/chany_top_out[7] sb_8__0_/chany_top_out[8] sb_8__0_/chany_top_out[9]
+ sb_8__0_/left_bottom_grid_pin_11_ sb_8__0_/left_bottom_grid_pin_13_ sb_8__0_/left_bottom_grid_pin_15_
+ sb_8__0_/left_bottom_grid_pin_17_ sb_8__0_/left_bottom_grid_pin_1_ sb_8__0_/left_bottom_grid_pin_3_
+ sb_8__0_/left_bottom_grid_pin_5_ sb_8__0_/left_bottom_grid_pin_7_ sb_8__0_/left_bottom_grid_pin_9_
+ sb_8__0_/prog_clk_0_N_in sb_8__0_/top_left_grid_pin_42_ sb_8__0_/top_left_grid_pin_43_
+ sb_8__0_/top_left_grid_pin_44_ sb_8__0_/top_left_grid_pin_45_ sb_8__0_/top_left_grid_pin_46_
+ sb_8__0_/top_left_grid_pin_47_ sb_8__0_/top_left_grid_pin_48_ sb_8__0_/top_left_grid_pin_49_
+ sb_8__0_/top_right_grid_pin_1_ sb_2__0_
Xsb_4__8_ sb_4__8_/SC_IN_BOT sb_4__8_/SC_OUT_BOT VGND VPWR sb_4__8_/bottom_left_grid_pin_42_
+ sb_4__8_/bottom_left_grid_pin_43_ sb_4__8_/bottom_left_grid_pin_44_ sb_4__8_/bottom_left_grid_pin_45_
+ sb_4__8_/bottom_left_grid_pin_46_ sb_4__8_/bottom_left_grid_pin_47_ sb_4__8_/bottom_left_grid_pin_48_
+ sb_4__8_/bottom_left_grid_pin_49_ sb_4__8_/ccff_head sb_4__8_/ccff_tail sb_4__8_/chanx_left_in[0]
+ sb_4__8_/chanx_left_in[10] sb_4__8_/chanx_left_in[11] sb_4__8_/chanx_left_in[12]
+ sb_4__8_/chanx_left_in[13] sb_4__8_/chanx_left_in[14] sb_4__8_/chanx_left_in[15]
+ sb_4__8_/chanx_left_in[16] sb_4__8_/chanx_left_in[17] sb_4__8_/chanx_left_in[18]
+ sb_4__8_/chanx_left_in[19] sb_4__8_/chanx_left_in[1] sb_4__8_/chanx_left_in[2] sb_4__8_/chanx_left_in[3]
+ sb_4__8_/chanx_left_in[4] sb_4__8_/chanx_left_in[5] sb_4__8_/chanx_left_in[6] sb_4__8_/chanx_left_in[7]
+ sb_4__8_/chanx_left_in[8] sb_4__8_/chanx_left_in[9] sb_4__8_/chanx_left_out[0] sb_4__8_/chanx_left_out[10]
+ sb_4__8_/chanx_left_out[11] sb_4__8_/chanx_left_out[12] sb_4__8_/chanx_left_out[13]
+ sb_4__8_/chanx_left_out[14] sb_4__8_/chanx_left_out[15] sb_4__8_/chanx_left_out[16]
+ sb_4__8_/chanx_left_out[17] sb_4__8_/chanx_left_out[18] sb_4__8_/chanx_left_out[19]
+ sb_4__8_/chanx_left_out[1] sb_4__8_/chanx_left_out[2] sb_4__8_/chanx_left_out[3]
+ sb_4__8_/chanx_left_out[4] sb_4__8_/chanx_left_out[5] sb_4__8_/chanx_left_out[6]
+ sb_4__8_/chanx_left_out[7] sb_4__8_/chanx_left_out[8] sb_4__8_/chanx_left_out[9]
+ sb_4__8_/chanx_right_in[0] sb_4__8_/chanx_right_in[10] sb_4__8_/chanx_right_in[11]
+ sb_4__8_/chanx_right_in[12] sb_4__8_/chanx_right_in[13] sb_4__8_/chanx_right_in[14]
+ sb_4__8_/chanx_right_in[15] sb_4__8_/chanx_right_in[16] sb_4__8_/chanx_right_in[17]
+ sb_4__8_/chanx_right_in[18] sb_4__8_/chanx_right_in[19] sb_4__8_/chanx_right_in[1]
+ sb_4__8_/chanx_right_in[2] sb_4__8_/chanx_right_in[3] sb_4__8_/chanx_right_in[4]
+ sb_4__8_/chanx_right_in[5] sb_4__8_/chanx_right_in[6] sb_4__8_/chanx_right_in[7]
+ sb_4__8_/chanx_right_in[8] sb_4__8_/chanx_right_in[9] cbx_5__8_/chanx_left_in[0]
+ cbx_5__8_/chanx_left_in[10] cbx_5__8_/chanx_left_in[11] cbx_5__8_/chanx_left_in[12]
+ cbx_5__8_/chanx_left_in[13] cbx_5__8_/chanx_left_in[14] cbx_5__8_/chanx_left_in[15]
+ cbx_5__8_/chanx_left_in[16] cbx_5__8_/chanx_left_in[17] cbx_5__8_/chanx_left_in[18]
+ cbx_5__8_/chanx_left_in[19] cbx_5__8_/chanx_left_in[1] cbx_5__8_/chanx_left_in[2]
+ cbx_5__8_/chanx_left_in[3] cbx_5__8_/chanx_left_in[4] cbx_5__8_/chanx_left_in[5]
+ cbx_5__8_/chanx_left_in[6] cbx_5__8_/chanx_left_in[7] cbx_5__8_/chanx_left_in[8]
+ cbx_5__8_/chanx_left_in[9] cby_4__8_/chany_top_out[0] cby_4__8_/chany_top_out[10]
+ cby_4__8_/chany_top_out[11] cby_4__8_/chany_top_out[12] cby_4__8_/chany_top_out[13]
+ cby_4__8_/chany_top_out[14] cby_4__8_/chany_top_out[15] cby_4__8_/chany_top_out[16]
+ cby_4__8_/chany_top_out[17] cby_4__8_/chany_top_out[18] cby_4__8_/chany_top_out[19]
+ cby_4__8_/chany_top_out[1] cby_4__8_/chany_top_out[2] cby_4__8_/chany_top_out[3]
+ cby_4__8_/chany_top_out[4] cby_4__8_/chany_top_out[5] cby_4__8_/chany_top_out[6]
+ cby_4__8_/chany_top_out[7] cby_4__8_/chany_top_out[8] cby_4__8_/chany_top_out[9]
+ cby_4__8_/chany_top_in[0] cby_4__8_/chany_top_in[10] cby_4__8_/chany_top_in[11]
+ cby_4__8_/chany_top_in[12] cby_4__8_/chany_top_in[13] cby_4__8_/chany_top_in[14]
+ cby_4__8_/chany_top_in[15] cby_4__8_/chany_top_in[16] cby_4__8_/chany_top_in[17]
+ cby_4__8_/chany_top_in[18] cby_4__8_/chany_top_in[19] cby_4__8_/chany_top_in[1]
+ cby_4__8_/chany_top_in[2] cby_4__8_/chany_top_in[3] cby_4__8_/chany_top_in[4] cby_4__8_/chany_top_in[5]
+ cby_4__8_/chany_top_in[6] cby_4__8_/chany_top_in[7] cby_4__8_/chany_top_in[8] cby_4__8_/chany_top_in[9]
+ sb_4__8_/left_bottom_grid_pin_34_ sb_4__8_/left_bottom_grid_pin_35_ sb_4__8_/left_bottom_grid_pin_36_
+ sb_4__8_/left_bottom_grid_pin_37_ sb_4__8_/left_bottom_grid_pin_38_ sb_4__8_/left_bottom_grid_pin_39_
+ sb_4__8_/left_bottom_grid_pin_40_ sb_4__8_/left_bottom_grid_pin_41_ sb_4__8_/left_top_grid_pin_1_
+ sb_4__8_/prog_clk_0_S_in sb_4__8_/right_bottom_grid_pin_34_ sb_4__8_/right_bottom_grid_pin_35_
+ sb_4__8_/right_bottom_grid_pin_36_ sb_4__8_/right_bottom_grid_pin_37_ sb_4__8_/right_bottom_grid_pin_38_
+ sb_4__8_/right_bottom_grid_pin_39_ sb_4__8_/right_bottom_grid_pin_40_ sb_4__8_/right_bottom_grid_pin_41_
+ sb_4__8_/right_top_grid_pin_1_ sb_1__2_
Xsb_1__5_ sb_1__5_/Test_en_N_out sb_1__5_/Test_en_S_in VGND VPWR sb_1__5_/bottom_left_grid_pin_42_
+ sb_1__5_/bottom_left_grid_pin_43_ sb_1__5_/bottom_left_grid_pin_44_ sb_1__5_/bottom_left_grid_pin_45_
+ sb_1__5_/bottom_left_grid_pin_46_ sb_1__5_/bottom_left_grid_pin_47_ sb_1__5_/bottom_left_grid_pin_48_
+ sb_1__5_/bottom_left_grid_pin_49_ sb_1__5_/ccff_head sb_1__5_/ccff_tail sb_1__5_/chanx_left_in[0]
+ sb_1__5_/chanx_left_in[10] sb_1__5_/chanx_left_in[11] sb_1__5_/chanx_left_in[12]
+ sb_1__5_/chanx_left_in[13] sb_1__5_/chanx_left_in[14] sb_1__5_/chanx_left_in[15]
+ sb_1__5_/chanx_left_in[16] sb_1__5_/chanx_left_in[17] sb_1__5_/chanx_left_in[18]
+ sb_1__5_/chanx_left_in[19] sb_1__5_/chanx_left_in[1] sb_1__5_/chanx_left_in[2] sb_1__5_/chanx_left_in[3]
+ sb_1__5_/chanx_left_in[4] sb_1__5_/chanx_left_in[5] sb_1__5_/chanx_left_in[6] sb_1__5_/chanx_left_in[7]
+ sb_1__5_/chanx_left_in[8] sb_1__5_/chanx_left_in[9] sb_1__5_/chanx_left_out[0] sb_1__5_/chanx_left_out[10]
+ sb_1__5_/chanx_left_out[11] sb_1__5_/chanx_left_out[12] sb_1__5_/chanx_left_out[13]
+ sb_1__5_/chanx_left_out[14] sb_1__5_/chanx_left_out[15] sb_1__5_/chanx_left_out[16]
+ sb_1__5_/chanx_left_out[17] sb_1__5_/chanx_left_out[18] sb_1__5_/chanx_left_out[19]
+ sb_1__5_/chanx_left_out[1] sb_1__5_/chanx_left_out[2] sb_1__5_/chanx_left_out[3]
+ sb_1__5_/chanx_left_out[4] sb_1__5_/chanx_left_out[5] sb_1__5_/chanx_left_out[6]
+ sb_1__5_/chanx_left_out[7] sb_1__5_/chanx_left_out[8] sb_1__5_/chanx_left_out[9]
+ sb_1__5_/chanx_right_in[0] sb_1__5_/chanx_right_in[10] sb_1__5_/chanx_right_in[11]
+ sb_1__5_/chanx_right_in[12] sb_1__5_/chanx_right_in[13] sb_1__5_/chanx_right_in[14]
+ sb_1__5_/chanx_right_in[15] sb_1__5_/chanx_right_in[16] sb_1__5_/chanx_right_in[17]
+ sb_1__5_/chanx_right_in[18] sb_1__5_/chanx_right_in[19] sb_1__5_/chanx_right_in[1]
+ sb_1__5_/chanx_right_in[2] sb_1__5_/chanx_right_in[3] sb_1__5_/chanx_right_in[4]
+ sb_1__5_/chanx_right_in[5] sb_1__5_/chanx_right_in[6] sb_1__5_/chanx_right_in[7]
+ sb_1__5_/chanx_right_in[8] sb_1__5_/chanx_right_in[9] cbx_2__5_/chanx_left_in[0]
+ cbx_2__5_/chanx_left_in[10] cbx_2__5_/chanx_left_in[11] cbx_2__5_/chanx_left_in[12]
+ cbx_2__5_/chanx_left_in[13] cbx_2__5_/chanx_left_in[14] cbx_2__5_/chanx_left_in[15]
+ cbx_2__5_/chanx_left_in[16] cbx_2__5_/chanx_left_in[17] cbx_2__5_/chanx_left_in[18]
+ cbx_2__5_/chanx_left_in[19] cbx_2__5_/chanx_left_in[1] cbx_2__5_/chanx_left_in[2]
+ cbx_2__5_/chanx_left_in[3] cbx_2__5_/chanx_left_in[4] cbx_2__5_/chanx_left_in[5]
+ cbx_2__5_/chanx_left_in[6] cbx_2__5_/chanx_left_in[7] cbx_2__5_/chanx_left_in[8]
+ cbx_2__5_/chanx_left_in[9] cby_1__5_/chany_top_out[0] cby_1__5_/chany_top_out[10]
+ cby_1__5_/chany_top_out[11] cby_1__5_/chany_top_out[12] cby_1__5_/chany_top_out[13]
+ cby_1__5_/chany_top_out[14] cby_1__5_/chany_top_out[15] cby_1__5_/chany_top_out[16]
+ cby_1__5_/chany_top_out[17] cby_1__5_/chany_top_out[18] cby_1__5_/chany_top_out[19]
+ cby_1__5_/chany_top_out[1] cby_1__5_/chany_top_out[2] cby_1__5_/chany_top_out[3]
+ cby_1__5_/chany_top_out[4] cby_1__5_/chany_top_out[5] cby_1__5_/chany_top_out[6]
+ cby_1__5_/chany_top_out[7] cby_1__5_/chany_top_out[8] cby_1__5_/chany_top_out[9]
+ cby_1__5_/chany_top_in[0] cby_1__5_/chany_top_in[10] cby_1__5_/chany_top_in[11]
+ cby_1__5_/chany_top_in[12] cby_1__5_/chany_top_in[13] cby_1__5_/chany_top_in[14]
+ cby_1__5_/chany_top_in[15] cby_1__5_/chany_top_in[16] cby_1__5_/chany_top_in[17]
+ cby_1__5_/chany_top_in[18] cby_1__5_/chany_top_in[19] cby_1__5_/chany_top_in[1]
+ cby_1__5_/chany_top_in[2] cby_1__5_/chany_top_in[3] cby_1__5_/chany_top_in[4] cby_1__5_/chany_top_in[5]
+ cby_1__5_/chany_top_in[6] cby_1__5_/chany_top_in[7] cby_1__5_/chany_top_in[8] cby_1__5_/chany_top_in[9]
+ sb_1__5_/chany_top_in[0] sb_1__5_/chany_top_in[10] sb_1__5_/chany_top_in[11] sb_1__5_/chany_top_in[12]
+ sb_1__5_/chany_top_in[13] sb_1__5_/chany_top_in[14] sb_1__5_/chany_top_in[15] sb_1__5_/chany_top_in[16]
+ sb_1__5_/chany_top_in[17] sb_1__5_/chany_top_in[18] sb_1__5_/chany_top_in[19] sb_1__5_/chany_top_in[1]
+ sb_1__5_/chany_top_in[2] sb_1__5_/chany_top_in[3] sb_1__5_/chany_top_in[4] sb_1__5_/chany_top_in[5]
+ sb_1__5_/chany_top_in[6] sb_1__5_/chany_top_in[7] sb_1__5_/chany_top_in[8] sb_1__5_/chany_top_in[9]
+ sb_1__5_/chany_top_out[0] sb_1__5_/chany_top_out[10] sb_1__5_/chany_top_out[11]
+ sb_1__5_/chany_top_out[12] sb_1__5_/chany_top_out[13] sb_1__5_/chany_top_out[14]
+ sb_1__5_/chany_top_out[15] sb_1__5_/chany_top_out[16] sb_1__5_/chany_top_out[17]
+ sb_1__5_/chany_top_out[18] sb_1__5_/chany_top_out[19] sb_1__5_/chany_top_out[1]
+ sb_1__5_/chany_top_out[2] sb_1__5_/chany_top_out[3] sb_1__5_/chany_top_out[4] sb_1__5_/chany_top_out[5]
+ sb_1__5_/chany_top_out[6] sb_1__5_/chany_top_out[7] sb_1__5_/chany_top_out[8] sb_1__5_/chany_top_out[9]
+ sb_1__5_/clk_1_E_out sb_1__5_/clk_1_N_in sb_1__5_/clk_1_W_out sb_1__5_/clk_2_E_out
+ sb_1__5_/clk_2_N_in sb_1__5_/clk_2_N_out sb_1__5_/clk_2_S_out sb_1__5_/clk_2_W_out
+ sb_1__5_/clk_3_E_out sb_1__5_/clk_3_N_in sb_1__5_/clk_3_N_out sb_1__5_/clk_3_S_out
+ sb_1__5_/clk_3_W_out sb_1__5_/left_bottom_grid_pin_34_ sb_1__5_/left_bottom_grid_pin_35_
+ sb_1__5_/left_bottom_grid_pin_36_ sb_1__5_/left_bottom_grid_pin_37_ sb_1__5_/left_bottom_grid_pin_38_
+ sb_1__5_/left_bottom_grid_pin_39_ sb_1__5_/left_bottom_grid_pin_40_ sb_1__5_/left_bottom_grid_pin_41_
+ sb_1__5_/prog_clk_0_N_in sb_1__5_/prog_clk_1_E_out sb_1__5_/prog_clk_1_N_in sb_1__5_/prog_clk_1_W_out
+ sb_1__5_/prog_clk_2_E_out sb_1__5_/prog_clk_2_N_in sb_1__5_/prog_clk_2_N_out sb_1__5_/prog_clk_2_S_out
+ sb_1__5_/prog_clk_2_W_out sb_1__5_/prog_clk_3_E_out sb_1__5_/prog_clk_3_N_in sb_1__5_/prog_clk_3_N_out
+ sb_1__5_/prog_clk_3_S_out sb_1__5_/prog_clk_3_W_out sb_1__5_/right_bottom_grid_pin_34_
+ sb_1__5_/right_bottom_grid_pin_35_ sb_1__5_/right_bottom_grid_pin_36_ sb_1__5_/right_bottom_grid_pin_37_
+ sb_1__5_/right_bottom_grid_pin_38_ sb_1__5_/right_bottom_grid_pin_39_ sb_1__5_/right_bottom_grid_pin_40_
+ sb_1__5_/right_bottom_grid_pin_41_ sb_1__5_/top_left_grid_pin_42_ sb_1__5_/top_left_grid_pin_43_
+ sb_1__5_/top_left_grid_pin_44_ sb_1__5_/top_left_grid_pin_45_ sb_1__5_/top_left_grid_pin_46_
+ sb_1__5_/top_left_grid_pin_47_ sb_1__5_/top_left_grid_pin_48_ sb_1__5_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_3__3_ cbx_3__3_/SC_OUT_BOT cbx_3__2_/SC_IN_TOP grid_clb_3__3_/SC_OUT_TOP
+ cby_3__3_/Test_en_W_out grid_clb_3__3_/Test_en_E_out cby_3__3_/Test_en_W_out cby_2__3_/Test_en_W_in
+ VGND VPWR cbx_3__2_/REGIN_FEEDTHROUGH grid_clb_3__3_/bottom_width_0_height_0__pin_51_
+ cby_2__3_/ccff_tail cby_3__3_/ccff_head cbx_3__3_/clk_1_S_out cbx_3__3_/clk_1_S_out
+ cby_3__3_/prog_clk_0_W_in cbx_3__3_/prog_clk_1_S_out grid_clb_3__3_/prog_clk_0_N_out
+ cbx_3__3_/prog_clk_1_S_out cbx_3__2_/prog_clk_0_N_in grid_clb_3__3_/prog_clk_0_W_out
+ cby_3__3_/left_grid_pin_16_ cby_3__3_/left_grid_pin_17_ cby_3__3_/left_grid_pin_18_
+ cby_3__3_/left_grid_pin_19_ cby_3__3_/left_grid_pin_20_ cby_3__3_/left_grid_pin_21_
+ cby_3__3_/left_grid_pin_22_ cby_3__3_/left_grid_pin_23_ cby_3__3_/left_grid_pin_24_
+ cby_3__3_/left_grid_pin_25_ cby_3__3_/left_grid_pin_26_ cby_3__3_/left_grid_pin_27_
+ cby_3__3_/left_grid_pin_28_ cby_3__3_/left_grid_pin_29_ cby_3__3_/left_grid_pin_30_
+ cby_3__3_/left_grid_pin_31_ sb_3__2_/top_left_grid_pin_42_ sb_3__3_/bottom_left_grid_pin_42_
+ sb_3__2_/top_left_grid_pin_43_ sb_3__3_/bottom_left_grid_pin_43_ sb_3__2_/top_left_grid_pin_44_
+ sb_3__3_/bottom_left_grid_pin_44_ sb_3__2_/top_left_grid_pin_45_ sb_3__3_/bottom_left_grid_pin_45_
+ sb_3__2_/top_left_grid_pin_46_ sb_3__3_/bottom_left_grid_pin_46_ sb_3__2_/top_left_grid_pin_47_
+ sb_3__3_/bottom_left_grid_pin_47_ sb_3__2_/top_left_grid_pin_48_ sb_3__3_/bottom_left_grid_pin_48_
+ sb_3__2_/top_left_grid_pin_49_ sb_3__3_/bottom_left_grid_pin_49_ cbx_3__3_/bottom_grid_pin_0_
+ cbx_3__3_/bottom_grid_pin_10_ cbx_3__3_/bottom_grid_pin_11_ cbx_3__3_/bottom_grid_pin_12_
+ cbx_3__3_/bottom_grid_pin_13_ cbx_3__3_/bottom_grid_pin_14_ cbx_3__3_/bottom_grid_pin_15_
+ cbx_3__3_/bottom_grid_pin_1_ cbx_3__3_/bottom_grid_pin_2_ cbx_3__3_/REGOUT_FEEDTHROUGH
+ grid_clb_3__3_/top_width_0_height_0__pin_33_ sb_3__3_/left_bottom_grid_pin_34_ sb_2__3_/right_bottom_grid_pin_34_
+ sb_3__3_/left_bottom_grid_pin_35_ sb_2__3_/right_bottom_grid_pin_35_ sb_3__3_/left_bottom_grid_pin_36_
+ sb_2__3_/right_bottom_grid_pin_36_ sb_3__3_/left_bottom_grid_pin_37_ sb_2__3_/right_bottom_grid_pin_37_
+ sb_3__3_/left_bottom_grid_pin_38_ sb_2__3_/right_bottom_grid_pin_38_ sb_3__3_/left_bottom_grid_pin_39_
+ sb_2__3_/right_bottom_grid_pin_39_ cbx_3__3_/bottom_grid_pin_3_ sb_3__3_/left_bottom_grid_pin_40_
+ sb_2__3_/right_bottom_grid_pin_40_ sb_3__3_/left_bottom_grid_pin_41_ sb_2__3_/right_bottom_grid_pin_41_
+ cbx_3__3_/bottom_grid_pin_4_ cbx_3__3_/bottom_grid_pin_5_ cbx_3__3_/bottom_grid_pin_6_
+ cbx_3__3_/bottom_grid_pin_7_ cbx_3__3_/bottom_grid_pin_8_ cbx_3__3_/bottom_grid_pin_9_
+ grid_clb
Xcby_7__4_ cby_7__4_/Test_en_W_in cby_7__4_/Test_en_E_out cby_7__4_/Test_en_N_out
+ cby_7__4_/Test_en_W_in cby_7__4_/Test_en_W_in cby_7__4_/Test_en_W_out VGND VPWR
+ cby_7__4_/ccff_head cby_7__4_/ccff_tail sb_7__3_/chany_top_out[0] sb_7__3_/chany_top_out[10]
+ sb_7__3_/chany_top_out[11] sb_7__3_/chany_top_out[12] sb_7__3_/chany_top_out[13]
+ sb_7__3_/chany_top_out[14] sb_7__3_/chany_top_out[15] sb_7__3_/chany_top_out[16]
+ sb_7__3_/chany_top_out[17] sb_7__3_/chany_top_out[18] sb_7__3_/chany_top_out[19]
+ sb_7__3_/chany_top_out[1] sb_7__3_/chany_top_out[2] sb_7__3_/chany_top_out[3] sb_7__3_/chany_top_out[4]
+ sb_7__3_/chany_top_out[5] sb_7__3_/chany_top_out[6] sb_7__3_/chany_top_out[7] sb_7__3_/chany_top_out[8]
+ sb_7__3_/chany_top_out[9] sb_7__3_/chany_top_in[0] sb_7__3_/chany_top_in[10] sb_7__3_/chany_top_in[11]
+ sb_7__3_/chany_top_in[12] sb_7__3_/chany_top_in[13] sb_7__3_/chany_top_in[14] sb_7__3_/chany_top_in[15]
+ sb_7__3_/chany_top_in[16] sb_7__3_/chany_top_in[17] sb_7__3_/chany_top_in[18] sb_7__3_/chany_top_in[19]
+ sb_7__3_/chany_top_in[1] sb_7__3_/chany_top_in[2] sb_7__3_/chany_top_in[3] sb_7__3_/chany_top_in[4]
+ sb_7__3_/chany_top_in[5] sb_7__3_/chany_top_in[6] sb_7__3_/chany_top_in[7] sb_7__3_/chany_top_in[8]
+ sb_7__3_/chany_top_in[9] cby_7__4_/chany_top_in[0] cby_7__4_/chany_top_in[10] cby_7__4_/chany_top_in[11]
+ cby_7__4_/chany_top_in[12] cby_7__4_/chany_top_in[13] cby_7__4_/chany_top_in[14]
+ cby_7__4_/chany_top_in[15] cby_7__4_/chany_top_in[16] cby_7__4_/chany_top_in[17]
+ cby_7__4_/chany_top_in[18] cby_7__4_/chany_top_in[19] cby_7__4_/chany_top_in[1]
+ cby_7__4_/chany_top_in[2] cby_7__4_/chany_top_in[3] cby_7__4_/chany_top_in[4] cby_7__4_/chany_top_in[5]
+ cby_7__4_/chany_top_in[6] cby_7__4_/chany_top_in[7] cby_7__4_/chany_top_in[8] cby_7__4_/chany_top_in[9]
+ cby_7__4_/chany_top_out[0] cby_7__4_/chany_top_out[10] cby_7__4_/chany_top_out[11]
+ cby_7__4_/chany_top_out[12] cby_7__4_/chany_top_out[13] cby_7__4_/chany_top_out[14]
+ cby_7__4_/chany_top_out[15] cby_7__4_/chany_top_out[16] cby_7__4_/chany_top_out[17]
+ cby_7__4_/chany_top_out[18] cby_7__4_/chany_top_out[19] cby_7__4_/chany_top_out[1]
+ cby_7__4_/chany_top_out[2] cby_7__4_/chany_top_out[3] cby_7__4_/chany_top_out[4]
+ cby_7__4_/chany_top_out[5] cby_7__4_/chany_top_out[6] cby_7__4_/chany_top_out[7]
+ cby_7__4_/chany_top_out[8] cby_7__4_/chany_top_out[9] cby_7__4_/clk_2_N_out cby_7__4_/clk_2_S_in
+ cby_7__4_/clk_2_S_out cby_7__4_/clk_3_N_out cby_7__4_/clk_3_S_in cby_7__4_/clk_3_S_out
+ cby_7__4_/left_grid_pin_16_ cby_7__4_/left_grid_pin_17_ cby_7__4_/left_grid_pin_18_
+ cby_7__4_/left_grid_pin_19_ cby_7__4_/left_grid_pin_20_ cby_7__4_/left_grid_pin_21_
+ cby_7__4_/left_grid_pin_22_ cby_7__4_/left_grid_pin_23_ cby_7__4_/left_grid_pin_24_
+ cby_7__4_/left_grid_pin_25_ cby_7__4_/left_grid_pin_26_ cby_7__4_/left_grid_pin_27_
+ cby_7__4_/left_grid_pin_28_ cby_7__4_/left_grid_pin_29_ cby_7__4_/left_grid_pin_30_
+ cby_7__4_/left_grid_pin_31_ cby_7__4_/prog_clk_0_N_out sb_7__3_/prog_clk_0_N_in
+ cby_7__4_/prog_clk_0_W_in cby_7__4_/prog_clk_2_N_out cby_7__4_/prog_clk_2_S_in cby_7__4_/prog_clk_2_S_out
+ cby_7__4_/prog_clk_3_N_out cby_7__4_/prog_clk_3_S_in cby_7__4_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_7__5_ cbx_7__5_/REGIN_FEEDTHROUGH cbx_7__5_/REGOUT_FEEDTHROUGH cbx_7__5_/SC_IN_BOT
+ cbx_7__5_/SC_IN_TOP cbx_7__5_/SC_OUT_BOT cbx_7__5_/SC_OUT_TOP VGND VPWR cbx_7__5_/bottom_grid_pin_0_
+ cbx_7__5_/bottom_grid_pin_10_ cbx_7__5_/bottom_grid_pin_11_ cbx_7__5_/bottom_grid_pin_12_
+ cbx_7__5_/bottom_grid_pin_13_ cbx_7__5_/bottom_grid_pin_14_ cbx_7__5_/bottom_grid_pin_15_
+ cbx_7__5_/bottom_grid_pin_1_ cbx_7__5_/bottom_grid_pin_2_ cbx_7__5_/bottom_grid_pin_3_
+ cbx_7__5_/bottom_grid_pin_4_ cbx_7__5_/bottom_grid_pin_5_ cbx_7__5_/bottom_grid_pin_6_
+ cbx_7__5_/bottom_grid_pin_7_ cbx_7__5_/bottom_grid_pin_8_ cbx_7__5_/bottom_grid_pin_9_
+ sb_7__5_/ccff_tail sb_6__5_/ccff_head cbx_7__5_/chanx_left_in[0] cbx_7__5_/chanx_left_in[10]
+ cbx_7__5_/chanx_left_in[11] cbx_7__5_/chanx_left_in[12] cbx_7__5_/chanx_left_in[13]
+ cbx_7__5_/chanx_left_in[14] cbx_7__5_/chanx_left_in[15] cbx_7__5_/chanx_left_in[16]
+ cbx_7__5_/chanx_left_in[17] cbx_7__5_/chanx_left_in[18] cbx_7__5_/chanx_left_in[19]
+ cbx_7__5_/chanx_left_in[1] cbx_7__5_/chanx_left_in[2] cbx_7__5_/chanx_left_in[3]
+ cbx_7__5_/chanx_left_in[4] cbx_7__5_/chanx_left_in[5] cbx_7__5_/chanx_left_in[6]
+ cbx_7__5_/chanx_left_in[7] cbx_7__5_/chanx_left_in[8] cbx_7__5_/chanx_left_in[9]
+ sb_6__5_/chanx_right_in[0] sb_6__5_/chanx_right_in[10] sb_6__5_/chanx_right_in[11]
+ sb_6__5_/chanx_right_in[12] sb_6__5_/chanx_right_in[13] sb_6__5_/chanx_right_in[14]
+ sb_6__5_/chanx_right_in[15] sb_6__5_/chanx_right_in[16] sb_6__5_/chanx_right_in[17]
+ sb_6__5_/chanx_right_in[18] sb_6__5_/chanx_right_in[19] sb_6__5_/chanx_right_in[1]
+ sb_6__5_/chanx_right_in[2] sb_6__5_/chanx_right_in[3] sb_6__5_/chanx_right_in[4]
+ sb_6__5_/chanx_right_in[5] sb_6__5_/chanx_right_in[6] sb_6__5_/chanx_right_in[7]
+ sb_6__5_/chanx_right_in[8] sb_6__5_/chanx_right_in[9] sb_7__5_/chanx_left_out[0]
+ sb_7__5_/chanx_left_out[10] sb_7__5_/chanx_left_out[11] sb_7__5_/chanx_left_out[12]
+ sb_7__5_/chanx_left_out[13] sb_7__5_/chanx_left_out[14] sb_7__5_/chanx_left_out[15]
+ sb_7__5_/chanx_left_out[16] sb_7__5_/chanx_left_out[17] sb_7__5_/chanx_left_out[18]
+ sb_7__5_/chanx_left_out[19] sb_7__5_/chanx_left_out[1] sb_7__5_/chanx_left_out[2]
+ sb_7__5_/chanx_left_out[3] sb_7__5_/chanx_left_out[4] sb_7__5_/chanx_left_out[5]
+ sb_7__5_/chanx_left_out[6] sb_7__5_/chanx_left_out[7] sb_7__5_/chanx_left_out[8]
+ sb_7__5_/chanx_left_out[9] sb_7__5_/chanx_left_in[0] sb_7__5_/chanx_left_in[10]
+ sb_7__5_/chanx_left_in[11] sb_7__5_/chanx_left_in[12] sb_7__5_/chanx_left_in[13]
+ sb_7__5_/chanx_left_in[14] sb_7__5_/chanx_left_in[15] sb_7__5_/chanx_left_in[16]
+ sb_7__5_/chanx_left_in[17] sb_7__5_/chanx_left_in[18] sb_7__5_/chanx_left_in[19]
+ sb_7__5_/chanx_left_in[1] sb_7__5_/chanx_left_in[2] sb_7__5_/chanx_left_in[3] sb_7__5_/chanx_left_in[4]
+ sb_7__5_/chanx_left_in[5] sb_7__5_/chanx_left_in[6] sb_7__5_/chanx_left_in[7] sb_7__5_/chanx_left_in[8]
+ sb_7__5_/chanx_left_in[9] cbx_7__5_/clk_1_N_out cbx_7__5_/clk_1_S_out sb_7__5_/clk_1_W_out
+ cbx_7__5_/clk_2_E_out cbx_7__5_/clk_2_W_in cbx_7__5_/clk_2_W_out cbx_7__5_/clk_3_E_out
+ cbx_7__5_/clk_3_W_in cbx_7__5_/clk_3_W_out cbx_7__5_/prog_clk_0_N_in cbx_7__5_/prog_clk_0_W_out
+ cbx_7__5_/prog_clk_1_N_out cbx_7__5_/prog_clk_1_S_out sb_7__5_/prog_clk_1_W_out
+ cbx_7__5_/prog_clk_2_E_out cbx_7__5_/prog_clk_2_W_in cbx_7__5_/prog_clk_2_W_out
+ cbx_7__5_/prog_clk_3_E_out cbx_7__5_/prog_clk_3_W_in cbx_7__5_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_4__1_ sb_4__0_/Test_en_N_out cby_4__1_/Test_en_E_out sb_4__1_/Test_en_S_in sb_4__0_/Test_en_N_out
+ sb_4__0_/Test_en_N_out cby_4__1_/Test_en_W_out VGND VPWR cby_4__1_/ccff_head cby_4__1_/ccff_tail
+ sb_4__0_/chany_top_out[0] sb_4__0_/chany_top_out[10] sb_4__0_/chany_top_out[11]
+ sb_4__0_/chany_top_out[12] sb_4__0_/chany_top_out[13] sb_4__0_/chany_top_out[14]
+ sb_4__0_/chany_top_out[15] sb_4__0_/chany_top_out[16] sb_4__0_/chany_top_out[17]
+ sb_4__0_/chany_top_out[18] sb_4__0_/chany_top_out[19] sb_4__0_/chany_top_out[1]
+ sb_4__0_/chany_top_out[2] sb_4__0_/chany_top_out[3] sb_4__0_/chany_top_out[4] sb_4__0_/chany_top_out[5]
+ sb_4__0_/chany_top_out[6] sb_4__0_/chany_top_out[7] sb_4__0_/chany_top_out[8] sb_4__0_/chany_top_out[9]
+ sb_4__0_/chany_top_in[0] sb_4__0_/chany_top_in[10] sb_4__0_/chany_top_in[11] sb_4__0_/chany_top_in[12]
+ sb_4__0_/chany_top_in[13] sb_4__0_/chany_top_in[14] sb_4__0_/chany_top_in[15] sb_4__0_/chany_top_in[16]
+ sb_4__0_/chany_top_in[17] sb_4__0_/chany_top_in[18] sb_4__0_/chany_top_in[19] sb_4__0_/chany_top_in[1]
+ sb_4__0_/chany_top_in[2] sb_4__0_/chany_top_in[3] sb_4__0_/chany_top_in[4] sb_4__0_/chany_top_in[5]
+ sb_4__0_/chany_top_in[6] sb_4__0_/chany_top_in[7] sb_4__0_/chany_top_in[8] sb_4__0_/chany_top_in[9]
+ cby_4__1_/chany_top_in[0] cby_4__1_/chany_top_in[10] cby_4__1_/chany_top_in[11]
+ cby_4__1_/chany_top_in[12] cby_4__1_/chany_top_in[13] cby_4__1_/chany_top_in[14]
+ cby_4__1_/chany_top_in[15] cby_4__1_/chany_top_in[16] cby_4__1_/chany_top_in[17]
+ cby_4__1_/chany_top_in[18] cby_4__1_/chany_top_in[19] cby_4__1_/chany_top_in[1]
+ cby_4__1_/chany_top_in[2] cby_4__1_/chany_top_in[3] cby_4__1_/chany_top_in[4] cby_4__1_/chany_top_in[5]
+ cby_4__1_/chany_top_in[6] cby_4__1_/chany_top_in[7] cby_4__1_/chany_top_in[8] cby_4__1_/chany_top_in[9]
+ cby_4__1_/chany_top_out[0] cby_4__1_/chany_top_out[10] cby_4__1_/chany_top_out[11]
+ cby_4__1_/chany_top_out[12] cby_4__1_/chany_top_out[13] cby_4__1_/chany_top_out[14]
+ cby_4__1_/chany_top_out[15] cby_4__1_/chany_top_out[16] cby_4__1_/chany_top_out[17]
+ cby_4__1_/chany_top_out[18] cby_4__1_/chany_top_out[19] cby_4__1_/chany_top_out[1]
+ cby_4__1_/chany_top_out[2] cby_4__1_/chany_top_out[3] cby_4__1_/chany_top_out[4]
+ cby_4__1_/chany_top_out[5] cby_4__1_/chany_top_out[6] cby_4__1_/chany_top_out[7]
+ cby_4__1_/chany_top_out[8] cby_4__1_/chany_top_out[9] cby_4__1_/clk_2_N_out cby_4__1_/clk_2_S_in
+ cby_4__1_/clk_2_S_out sb_4__1_/clk_3_N_in sb_4__0_/clk_3_N_out cby_4__1_/clk_3_S_out
+ cby_4__1_/left_grid_pin_16_ cby_4__1_/left_grid_pin_17_ cby_4__1_/left_grid_pin_18_
+ cby_4__1_/left_grid_pin_19_ cby_4__1_/left_grid_pin_20_ cby_4__1_/left_grid_pin_21_
+ cby_4__1_/left_grid_pin_22_ cby_4__1_/left_grid_pin_23_ cby_4__1_/left_grid_pin_24_
+ cby_4__1_/left_grid_pin_25_ cby_4__1_/left_grid_pin_26_ cby_4__1_/left_grid_pin_27_
+ cby_4__1_/left_grid_pin_28_ cby_4__1_/left_grid_pin_29_ cby_4__1_/left_grid_pin_30_
+ cby_4__1_/left_grid_pin_31_ cby_4__1_/prog_clk_0_N_out sb_4__0_/prog_clk_0_N_in
+ cby_4__1_/prog_clk_0_W_in cby_4__1_/prog_clk_2_N_out cby_4__1_/prog_clk_2_S_in cby_4__1_/prog_clk_2_S_out
+ sb_4__1_/prog_clk_3_N_in sb_4__0_/prog_clk_3_N_out cby_4__1_/prog_clk_3_S_out cby_1__1_
Xsb_4__7_ sb_4__7_/Test_en_N_out sb_4__7_/Test_en_S_in VGND VPWR sb_4__7_/bottom_left_grid_pin_42_
+ sb_4__7_/bottom_left_grid_pin_43_ sb_4__7_/bottom_left_grid_pin_44_ sb_4__7_/bottom_left_grid_pin_45_
+ sb_4__7_/bottom_left_grid_pin_46_ sb_4__7_/bottom_left_grid_pin_47_ sb_4__7_/bottom_left_grid_pin_48_
+ sb_4__7_/bottom_left_grid_pin_49_ sb_4__7_/ccff_head sb_4__7_/ccff_tail sb_4__7_/chanx_left_in[0]
+ sb_4__7_/chanx_left_in[10] sb_4__7_/chanx_left_in[11] sb_4__7_/chanx_left_in[12]
+ sb_4__7_/chanx_left_in[13] sb_4__7_/chanx_left_in[14] sb_4__7_/chanx_left_in[15]
+ sb_4__7_/chanx_left_in[16] sb_4__7_/chanx_left_in[17] sb_4__7_/chanx_left_in[18]
+ sb_4__7_/chanx_left_in[19] sb_4__7_/chanx_left_in[1] sb_4__7_/chanx_left_in[2] sb_4__7_/chanx_left_in[3]
+ sb_4__7_/chanx_left_in[4] sb_4__7_/chanx_left_in[5] sb_4__7_/chanx_left_in[6] sb_4__7_/chanx_left_in[7]
+ sb_4__7_/chanx_left_in[8] sb_4__7_/chanx_left_in[9] sb_4__7_/chanx_left_out[0] sb_4__7_/chanx_left_out[10]
+ sb_4__7_/chanx_left_out[11] sb_4__7_/chanx_left_out[12] sb_4__7_/chanx_left_out[13]
+ sb_4__7_/chanx_left_out[14] sb_4__7_/chanx_left_out[15] sb_4__7_/chanx_left_out[16]
+ sb_4__7_/chanx_left_out[17] sb_4__7_/chanx_left_out[18] sb_4__7_/chanx_left_out[19]
+ sb_4__7_/chanx_left_out[1] sb_4__7_/chanx_left_out[2] sb_4__7_/chanx_left_out[3]
+ sb_4__7_/chanx_left_out[4] sb_4__7_/chanx_left_out[5] sb_4__7_/chanx_left_out[6]
+ sb_4__7_/chanx_left_out[7] sb_4__7_/chanx_left_out[8] sb_4__7_/chanx_left_out[9]
+ sb_4__7_/chanx_right_in[0] sb_4__7_/chanx_right_in[10] sb_4__7_/chanx_right_in[11]
+ sb_4__7_/chanx_right_in[12] sb_4__7_/chanx_right_in[13] sb_4__7_/chanx_right_in[14]
+ sb_4__7_/chanx_right_in[15] sb_4__7_/chanx_right_in[16] sb_4__7_/chanx_right_in[17]
+ sb_4__7_/chanx_right_in[18] sb_4__7_/chanx_right_in[19] sb_4__7_/chanx_right_in[1]
+ sb_4__7_/chanx_right_in[2] sb_4__7_/chanx_right_in[3] sb_4__7_/chanx_right_in[4]
+ sb_4__7_/chanx_right_in[5] sb_4__7_/chanx_right_in[6] sb_4__7_/chanx_right_in[7]
+ sb_4__7_/chanx_right_in[8] sb_4__7_/chanx_right_in[9] cbx_5__7_/chanx_left_in[0]
+ cbx_5__7_/chanx_left_in[10] cbx_5__7_/chanx_left_in[11] cbx_5__7_/chanx_left_in[12]
+ cbx_5__7_/chanx_left_in[13] cbx_5__7_/chanx_left_in[14] cbx_5__7_/chanx_left_in[15]
+ cbx_5__7_/chanx_left_in[16] cbx_5__7_/chanx_left_in[17] cbx_5__7_/chanx_left_in[18]
+ cbx_5__7_/chanx_left_in[19] cbx_5__7_/chanx_left_in[1] cbx_5__7_/chanx_left_in[2]
+ cbx_5__7_/chanx_left_in[3] cbx_5__7_/chanx_left_in[4] cbx_5__7_/chanx_left_in[5]
+ cbx_5__7_/chanx_left_in[6] cbx_5__7_/chanx_left_in[7] cbx_5__7_/chanx_left_in[8]
+ cbx_5__7_/chanx_left_in[9] cby_4__7_/chany_top_out[0] cby_4__7_/chany_top_out[10]
+ cby_4__7_/chany_top_out[11] cby_4__7_/chany_top_out[12] cby_4__7_/chany_top_out[13]
+ cby_4__7_/chany_top_out[14] cby_4__7_/chany_top_out[15] cby_4__7_/chany_top_out[16]
+ cby_4__7_/chany_top_out[17] cby_4__7_/chany_top_out[18] cby_4__7_/chany_top_out[19]
+ cby_4__7_/chany_top_out[1] cby_4__7_/chany_top_out[2] cby_4__7_/chany_top_out[3]
+ cby_4__7_/chany_top_out[4] cby_4__7_/chany_top_out[5] cby_4__7_/chany_top_out[6]
+ cby_4__7_/chany_top_out[7] cby_4__7_/chany_top_out[8] cby_4__7_/chany_top_out[9]
+ cby_4__7_/chany_top_in[0] cby_4__7_/chany_top_in[10] cby_4__7_/chany_top_in[11]
+ cby_4__7_/chany_top_in[12] cby_4__7_/chany_top_in[13] cby_4__7_/chany_top_in[14]
+ cby_4__7_/chany_top_in[15] cby_4__7_/chany_top_in[16] cby_4__7_/chany_top_in[17]
+ cby_4__7_/chany_top_in[18] cby_4__7_/chany_top_in[19] cby_4__7_/chany_top_in[1]
+ cby_4__7_/chany_top_in[2] cby_4__7_/chany_top_in[3] cby_4__7_/chany_top_in[4] cby_4__7_/chany_top_in[5]
+ cby_4__7_/chany_top_in[6] cby_4__7_/chany_top_in[7] cby_4__7_/chany_top_in[8] cby_4__7_/chany_top_in[9]
+ sb_4__7_/chany_top_in[0] sb_4__7_/chany_top_in[10] sb_4__7_/chany_top_in[11] sb_4__7_/chany_top_in[12]
+ sb_4__7_/chany_top_in[13] sb_4__7_/chany_top_in[14] sb_4__7_/chany_top_in[15] sb_4__7_/chany_top_in[16]
+ sb_4__7_/chany_top_in[17] sb_4__7_/chany_top_in[18] sb_4__7_/chany_top_in[19] sb_4__7_/chany_top_in[1]
+ sb_4__7_/chany_top_in[2] sb_4__7_/chany_top_in[3] sb_4__7_/chany_top_in[4] sb_4__7_/chany_top_in[5]
+ sb_4__7_/chany_top_in[6] sb_4__7_/chany_top_in[7] sb_4__7_/chany_top_in[8] sb_4__7_/chany_top_in[9]
+ sb_4__7_/chany_top_out[0] sb_4__7_/chany_top_out[10] sb_4__7_/chany_top_out[11]
+ sb_4__7_/chany_top_out[12] sb_4__7_/chany_top_out[13] sb_4__7_/chany_top_out[14]
+ sb_4__7_/chany_top_out[15] sb_4__7_/chany_top_out[16] sb_4__7_/chany_top_out[17]
+ sb_4__7_/chany_top_out[18] sb_4__7_/chany_top_out[19] sb_4__7_/chany_top_out[1]
+ sb_4__7_/chany_top_out[2] sb_4__7_/chany_top_out[3] sb_4__7_/chany_top_out[4] sb_4__7_/chany_top_out[5]
+ sb_4__7_/chany_top_out[6] sb_4__7_/chany_top_out[7] sb_4__7_/chany_top_out[8] sb_4__7_/chany_top_out[9]
+ sb_4__7_/clk_1_E_out sb_4__7_/clk_1_N_in sb_4__7_/clk_1_W_out sb_4__7_/clk_2_E_out
+ sb_4__7_/clk_2_N_in sb_4__7_/clk_2_N_out sb_4__7_/clk_2_S_out sb_4__7_/clk_2_W_out
+ sb_4__7_/clk_3_E_out sb_4__7_/clk_3_N_in sb_4__7_/clk_3_N_out sb_4__7_/clk_3_S_out
+ sb_4__7_/clk_3_W_out sb_4__7_/left_bottom_grid_pin_34_ sb_4__7_/left_bottom_grid_pin_35_
+ sb_4__7_/left_bottom_grid_pin_36_ sb_4__7_/left_bottom_grid_pin_37_ sb_4__7_/left_bottom_grid_pin_38_
+ sb_4__7_/left_bottom_grid_pin_39_ sb_4__7_/left_bottom_grid_pin_40_ sb_4__7_/left_bottom_grid_pin_41_
+ sb_4__7_/prog_clk_0_N_in sb_4__7_/prog_clk_1_E_out sb_4__7_/prog_clk_1_N_in sb_4__7_/prog_clk_1_W_out
+ sb_4__7_/prog_clk_2_E_out sb_4__7_/prog_clk_2_N_in sb_4__7_/prog_clk_2_N_out sb_4__7_/prog_clk_2_S_out
+ sb_4__7_/prog_clk_2_W_out sb_4__7_/prog_clk_3_E_out sb_4__7_/prog_clk_3_N_in sb_4__7_/prog_clk_3_N_out
+ sb_4__7_/prog_clk_3_S_out sb_4__7_/prog_clk_3_W_out sb_4__7_/right_bottom_grid_pin_34_
+ sb_4__7_/right_bottom_grid_pin_35_ sb_4__7_/right_bottom_grid_pin_36_ sb_4__7_/right_bottom_grid_pin_37_
+ sb_4__7_/right_bottom_grid_pin_38_ sb_4__7_/right_bottom_grid_pin_39_ sb_4__7_/right_bottom_grid_pin_40_
+ sb_4__7_/right_bottom_grid_pin_41_ sb_4__7_/top_left_grid_pin_42_ sb_4__7_/top_left_grid_pin_43_
+ sb_4__7_/top_left_grid_pin_44_ sb_4__7_/top_left_grid_pin_45_ sb_4__7_/top_left_grid_pin_46_
+ sb_4__7_/top_left_grid_pin_47_ sb_4__7_/top_left_grid_pin_48_ sb_4__7_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_6__5_ cbx_6__4_/SC_OUT_TOP grid_clb_6__5_/SC_OUT_BOT cbx_6__5_/SC_IN_BOT
+ cby_5__5_/Test_en_E_out cby_6__5_/Test_en_W_in cby_5__5_/Test_en_E_out grid_clb_6__5_/Test_en_W_out
+ VGND VPWR cbx_6__4_/REGIN_FEEDTHROUGH grid_clb_6__5_/bottom_width_0_height_0__pin_51_
+ cby_5__5_/ccff_tail cby_6__5_/ccff_head cbx_6__5_/clk_1_S_out cbx_6__5_/clk_1_S_out
+ cby_6__5_/prog_clk_0_W_in cbx_6__5_/prog_clk_1_S_out grid_clb_6__5_/prog_clk_0_N_out
+ cbx_6__5_/prog_clk_1_S_out cbx_6__4_/prog_clk_0_N_in grid_clb_6__5_/prog_clk_0_W_out
+ cby_6__5_/left_grid_pin_16_ cby_6__5_/left_grid_pin_17_ cby_6__5_/left_grid_pin_18_
+ cby_6__5_/left_grid_pin_19_ cby_6__5_/left_grid_pin_20_ cby_6__5_/left_grid_pin_21_
+ cby_6__5_/left_grid_pin_22_ cby_6__5_/left_grid_pin_23_ cby_6__5_/left_grid_pin_24_
+ cby_6__5_/left_grid_pin_25_ cby_6__5_/left_grid_pin_26_ cby_6__5_/left_grid_pin_27_
+ cby_6__5_/left_grid_pin_28_ cby_6__5_/left_grid_pin_29_ cby_6__5_/left_grid_pin_30_
+ cby_6__5_/left_grid_pin_31_ sb_6__4_/top_left_grid_pin_42_ sb_6__5_/bottom_left_grid_pin_42_
+ sb_6__4_/top_left_grid_pin_43_ sb_6__5_/bottom_left_grid_pin_43_ sb_6__4_/top_left_grid_pin_44_
+ sb_6__5_/bottom_left_grid_pin_44_ sb_6__4_/top_left_grid_pin_45_ sb_6__5_/bottom_left_grid_pin_45_
+ sb_6__4_/top_left_grid_pin_46_ sb_6__5_/bottom_left_grid_pin_46_ sb_6__4_/top_left_grid_pin_47_
+ sb_6__5_/bottom_left_grid_pin_47_ sb_6__4_/top_left_grid_pin_48_ sb_6__5_/bottom_left_grid_pin_48_
+ sb_6__4_/top_left_grid_pin_49_ sb_6__5_/bottom_left_grid_pin_49_ cbx_6__5_/bottom_grid_pin_0_
+ cbx_6__5_/bottom_grid_pin_10_ cbx_6__5_/bottom_grid_pin_11_ cbx_6__5_/bottom_grid_pin_12_
+ cbx_6__5_/bottom_grid_pin_13_ cbx_6__5_/bottom_grid_pin_14_ cbx_6__5_/bottom_grid_pin_15_
+ cbx_6__5_/bottom_grid_pin_1_ cbx_6__5_/bottom_grid_pin_2_ cbx_6__5_/REGOUT_FEEDTHROUGH
+ grid_clb_6__5_/top_width_0_height_0__pin_33_ sb_6__5_/left_bottom_grid_pin_34_ sb_5__5_/right_bottom_grid_pin_34_
+ sb_6__5_/left_bottom_grid_pin_35_ sb_5__5_/right_bottom_grid_pin_35_ sb_6__5_/left_bottom_grid_pin_36_
+ sb_5__5_/right_bottom_grid_pin_36_ sb_6__5_/left_bottom_grid_pin_37_ sb_5__5_/right_bottom_grid_pin_37_
+ sb_6__5_/left_bottom_grid_pin_38_ sb_5__5_/right_bottom_grid_pin_38_ sb_6__5_/left_bottom_grid_pin_39_
+ sb_5__5_/right_bottom_grid_pin_39_ cbx_6__5_/bottom_grid_pin_3_ sb_6__5_/left_bottom_grid_pin_40_
+ sb_5__5_/right_bottom_grid_pin_40_ sb_6__5_/left_bottom_grid_pin_41_ sb_5__5_/right_bottom_grid_pin_41_
+ cbx_6__5_/bottom_grid_pin_4_ cbx_6__5_/bottom_grid_pin_5_ cbx_6__5_/bottom_grid_pin_6_
+ cbx_6__5_/bottom_grid_pin_7_ cbx_6__5_/bottom_grid_pin_8_ cbx_6__5_/bottom_grid_pin_9_
+ grid_clb
Xgrid_clb_3__2_ cbx_3__2_/SC_OUT_BOT cbx_3__1_/SC_IN_TOP grid_clb_3__2_/SC_OUT_TOP
+ cby_3__2_/Test_en_W_out grid_clb_3__2_/Test_en_E_out cby_3__2_/Test_en_W_out cby_2__2_/Test_en_W_in
+ VGND VPWR cbx_3__1_/REGIN_FEEDTHROUGH grid_clb_3__2_/bottom_width_0_height_0__pin_51_
+ cby_2__2_/ccff_tail cby_3__2_/ccff_head cbx_3__1_/clk_1_N_out cbx_3__1_/clk_1_N_out
+ cby_3__2_/prog_clk_0_W_in cbx_3__1_/prog_clk_1_N_out grid_clb_3__2_/prog_clk_0_N_out
+ cbx_3__1_/prog_clk_1_N_out cbx_3__1_/prog_clk_0_N_in grid_clb_3__2_/prog_clk_0_W_out
+ cby_3__2_/left_grid_pin_16_ cby_3__2_/left_grid_pin_17_ cby_3__2_/left_grid_pin_18_
+ cby_3__2_/left_grid_pin_19_ cby_3__2_/left_grid_pin_20_ cby_3__2_/left_grid_pin_21_
+ cby_3__2_/left_grid_pin_22_ cby_3__2_/left_grid_pin_23_ cby_3__2_/left_grid_pin_24_
+ cby_3__2_/left_grid_pin_25_ cby_3__2_/left_grid_pin_26_ cby_3__2_/left_grid_pin_27_
+ cby_3__2_/left_grid_pin_28_ cby_3__2_/left_grid_pin_29_ cby_3__2_/left_grid_pin_30_
+ cby_3__2_/left_grid_pin_31_ sb_3__1_/top_left_grid_pin_42_ sb_3__2_/bottom_left_grid_pin_42_
+ sb_3__1_/top_left_grid_pin_43_ sb_3__2_/bottom_left_grid_pin_43_ sb_3__1_/top_left_grid_pin_44_
+ sb_3__2_/bottom_left_grid_pin_44_ sb_3__1_/top_left_grid_pin_45_ sb_3__2_/bottom_left_grid_pin_45_
+ sb_3__1_/top_left_grid_pin_46_ sb_3__2_/bottom_left_grid_pin_46_ sb_3__1_/top_left_grid_pin_47_
+ sb_3__2_/bottom_left_grid_pin_47_ sb_3__1_/top_left_grid_pin_48_ sb_3__2_/bottom_left_grid_pin_48_
+ sb_3__1_/top_left_grid_pin_49_ sb_3__2_/bottom_left_grid_pin_49_ cbx_3__2_/bottom_grid_pin_0_
+ cbx_3__2_/bottom_grid_pin_10_ cbx_3__2_/bottom_grid_pin_11_ cbx_3__2_/bottom_grid_pin_12_
+ cbx_3__2_/bottom_grid_pin_13_ cbx_3__2_/bottom_grid_pin_14_ cbx_3__2_/bottom_grid_pin_15_
+ cbx_3__2_/bottom_grid_pin_1_ cbx_3__2_/bottom_grid_pin_2_ cbx_3__2_/REGOUT_FEEDTHROUGH
+ grid_clb_3__2_/top_width_0_height_0__pin_33_ sb_3__2_/left_bottom_grid_pin_34_ sb_2__2_/right_bottom_grid_pin_34_
+ sb_3__2_/left_bottom_grid_pin_35_ sb_2__2_/right_bottom_grid_pin_35_ sb_3__2_/left_bottom_grid_pin_36_
+ sb_2__2_/right_bottom_grid_pin_36_ sb_3__2_/left_bottom_grid_pin_37_ sb_2__2_/right_bottom_grid_pin_37_
+ sb_3__2_/left_bottom_grid_pin_38_ sb_2__2_/right_bottom_grid_pin_38_ sb_3__2_/left_bottom_grid_pin_39_
+ sb_2__2_/right_bottom_grid_pin_39_ cbx_3__2_/bottom_grid_pin_3_ sb_3__2_/left_bottom_grid_pin_40_
+ sb_2__2_/right_bottom_grid_pin_40_ sb_3__2_/left_bottom_grid_pin_41_ sb_2__2_/right_bottom_grid_pin_41_
+ cbx_3__2_/bottom_grid_pin_4_ cbx_3__2_/bottom_grid_pin_5_ cbx_3__2_/bottom_grid_pin_6_
+ cbx_3__2_/bottom_grid_pin_7_ cbx_3__2_/bottom_grid_pin_8_ cbx_3__2_/bottom_grid_pin_9_
+ grid_clb
Xcbx_4__2_ cbx_4__2_/REGIN_FEEDTHROUGH cbx_4__2_/REGOUT_FEEDTHROUGH cbx_4__2_/SC_IN_BOT
+ cbx_4__2_/SC_IN_TOP cbx_4__2_/SC_OUT_BOT cbx_4__2_/SC_OUT_TOP VGND VPWR cbx_4__2_/bottom_grid_pin_0_
+ cbx_4__2_/bottom_grid_pin_10_ cbx_4__2_/bottom_grid_pin_11_ cbx_4__2_/bottom_grid_pin_12_
+ cbx_4__2_/bottom_grid_pin_13_ cbx_4__2_/bottom_grid_pin_14_ cbx_4__2_/bottom_grid_pin_15_
+ cbx_4__2_/bottom_grid_pin_1_ cbx_4__2_/bottom_grid_pin_2_ cbx_4__2_/bottom_grid_pin_3_
+ cbx_4__2_/bottom_grid_pin_4_ cbx_4__2_/bottom_grid_pin_5_ cbx_4__2_/bottom_grid_pin_6_
+ cbx_4__2_/bottom_grid_pin_7_ cbx_4__2_/bottom_grid_pin_8_ cbx_4__2_/bottom_grid_pin_9_
+ sb_4__2_/ccff_tail sb_3__2_/ccff_head cbx_4__2_/chanx_left_in[0] cbx_4__2_/chanx_left_in[10]
+ cbx_4__2_/chanx_left_in[11] cbx_4__2_/chanx_left_in[12] cbx_4__2_/chanx_left_in[13]
+ cbx_4__2_/chanx_left_in[14] cbx_4__2_/chanx_left_in[15] cbx_4__2_/chanx_left_in[16]
+ cbx_4__2_/chanx_left_in[17] cbx_4__2_/chanx_left_in[18] cbx_4__2_/chanx_left_in[19]
+ cbx_4__2_/chanx_left_in[1] cbx_4__2_/chanx_left_in[2] cbx_4__2_/chanx_left_in[3]
+ cbx_4__2_/chanx_left_in[4] cbx_4__2_/chanx_left_in[5] cbx_4__2_/chanx_left_in[6]
+ cbx_4__2_/chanx_left_in[7] cbx_4__2_/chanx_left_in[8] cbx_4__2_/chanx_left_in[9]
+ sb_3__2_/chanx_right_in[0] sb_3__2_/chanx_right_in[10] sb_3__2_/chanx_right_in[11]
+ sb_3__2_/chanx_right_in[12] sb_3__2_/chanx_right_in[13] sb_3__2_/chanx_right_in[14]
+ sb_3__2_/chanx_right_in[15] sb_3__2_/chanx_right_in[16] sb_3__2_/chanx_right_in[17]
+ sb_3__2_/chanx_right_in[18] sb_3__2_/chanx_right_in[19] sb_3__2_/chanx_right_in[1]
+ sb_3__2_/chanx_right_in[2] sb_3__2_/chanx_right_in[3] sb_3__2_/chanx_right_in[4]
+ sb_3__2_/chanx_right_in[5] sb_3__2_/chanx_right_in[6] sb_3__2_/chanx_right_in[7]
+ sb_3__2_/chanx_right_in[8] sb_3__2_/chanx_right_in[9] sb_4__2_/chanx_left_out[0]
+ sb_4__2_/chanx_left_out[10] sb_4__2_/chanx_left_out[11] sb_4__2_/chanx_left_out[12]
+ sb_4__2_/chanx_left_out[13] sb_4__2_/chanx_left_out[14] sb_4__2_/chanx_left_out[15]
+ sb_4__2_/chanx_left_out[16] sb_4__2_/chanx_left_out[17] sb_4__2_/chanx_left_out[18]
+ sb_4__2_/chanx_left_out[19] sb_4__2_/chanx_left_out[1] sb_4__2_/chanx_left_out[2]
+ sb_4__2_/chanx_left_out[3] sb_4__2_/chanx_left_out[4] sb_4__2_/chanx_left_out[5]
+ sb_4__2_/chanx_left_out[6] sb_4__2_/chanx_left_out[7] sb_4__2_/chanx_left_out[8]
+ sb_4__2_/chanx_left_out[9] sb_4__2_/chanx_left_in[0] sb_4__2_/chanx_left_in[10]
+ sb_4__2_/chanx_left_in[11] sb_4__2_/chanx_left_in[12] sb_4__2_/chanx_left_in[13]
+ sb_4__2_/chanx_left_in[14] sb_4__2_/chanx_left_in[15] sb_4__2_/chanx_left_in[16]
+ sb_4__2_/chanx_left_in[17] sb_4__2_/chanx_left_in[18] sb_4__2_/chanx_left_in[19]
+ sb_4__2_/chanx_left_in[1] sb_4__2_/chanx_left_in[2] sb_4__2_/chanx_left_in[3] sb_4__2_/chanx_left_in[4]
+ sb_4__2_/chanx_left_in[5] sb_4__2_/chanx_left_in[6] sb_4__2_/chanx_left_in[7] sb_4__2_/chanx_left_in[8]
+ sb_4__2_/chanx_left_in[9] cbx_4__2_/clk_1_N_out cbx_4__2_/clk_1_S_out cbx_4__2_/clk_1_W_in
+ cbx_4__2_/clk_2_E_out cbx_4__2_/clk_2_W_in cbx_4__2_/clk_2_W_out cbx_4__2_/clk_3_E_out
+ cbx_4__2_/clk_3_W_in cbx_4__2_/clk_3_W_out cbx_4__2_/prog_clk_0_N_in cbx_4__2_/prog_clk_0_W_out
+ cbx_4__2_/prog_clk_1_N_out cbx_4__2_/prog_clk_1_S_out cbx_4__2_/prog_clk_1_W_in
+ cbx_4__2_/prog_clk_2_E_out cbx_4__2_/prog_clk_2_W_in cbx_4__2_/prog_clk_2_W_out
+ cbx_4__2_/prog_clk_3_E_out cbx_4__2_/prog_clk_3_W_in cbx_4__2_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_1__4_ sb_1__4_/Test_en_N_out sb_1__4_/Test_en_S_in VGND VPWR sb_1__4_/bottom_left_grid_pin_42_
+ sb_1__4_/bottom_left_grid_pin_43_ sb_1__4_/bottom_left_grid_pin_44_ sb_1__4_/bottom_left_grid_pin_45_
+ sb_1__4_/bottom_left_grid_pin_46_ sb_1__4_/bottom_left_grid_pin_47_ sb_1__4_/bottom_left_grid_pin_48_
+ sb_1__4_/bottom_left_grid_pin_49_ sb_1__4_/ccff_head sb_1__4_/ccff_tail sb_1__4_/chanx_left_in[0]
+ sb_1__4_/chanx_left_in[10] sb_1__4_/chanx_left_in[11] sb_1__4_/chanx_left_in[12]
+ sb_1__4_/chanx_left_in[13] sb_1__4_/chanx_left_in[14] sb_1__4_/chanx_left_in[15]
+ sb_1__4_/chanx_left_in[16] sb_1__4_/chanx_left_in[17] sb_1__4_/chanx_left_in[18]
+ sb_1__4_/chanx_left_in[19] sb_1__4_/chanx_left_in[1] sb_1__4_/chanx_left_in[2] sb_1__4_/chanx_left_in[3]
+ sb_1__4_/chanx_left_in[4] sb_1__4_/chanx_left_in[5] sb_1__4_/chanx_left_in[6] sb_1__4_/chanx_left_in[7]
+ sb_1__4_/chanx_left_in[8] sb_1__4_/chanx_left_in[9] sb_1__4_/chanx_left_out[0] sb_1__4_/chanx_left_out[10]
+ sb_1__4_/chanx_left_out[11] sb_1__4_/chanx_left_out[12] sb_1__4_/chanx_left_out[13]
+ sb_1__4_/chanx_left_out[14] sb_1__4_/chanx_left_out[15] sb_1__4_/chanx_left_out[16]
+ sb_1__4_/chanx_left_out[17] sb_1__4_/chanx_left_out[18] sb_1__4_/chanx_left_out[19]
+ sb_1__4_/chanx_left_out[1] sb_1__4_/chanx_left_out[2] sb_1__4_/chanx_left_out[3]
+ sb_1__4_/chanx_left_out[4] sb_1__4_/chanx_left_out[5] sb_1__4_/chanx_left_out[6]
+ sb_1__4_/chanx_left_out[7] sb_1__4_/chanx_left_out[8] sb_1__4_/chanx_left_out[9]
+ sb_1__4_/chanx_right_in[0] sb_1__4_/chanx_right_in[10] sb_1__4_/chanx_right_in[11]
+ sb_1__4_/chanx_right_in[12] sb_1__4_/chanx_right_in[13] sb_1__4_/chanx_right_in[14]
+ sb_1__4_/chanx_right_in[15] sb_1__4_/chanx_right_in[16] sb_1__4_/chanx_right_in[17]
+ sb_1__4_/chanx_right_in[18] sb_1__4_/chanx_right_in[19] sb_1__4_/chanx_right_in[1]
+ sb_1__4_/chanx_right_in[2] sb_1__4_/chanx_right_in[3] sb_1__4_/chanx_right_in[4]
+ sb_1__4_/chanx_right_in[5] sb_1__4_/chanx_right_in[6] sb_1__4_/chanx_right_in[7]
+ sb_1__4_/chanx_right_in[8] sb_1__4_/chanx_right_in[9] cbx_2__4_/chanx_left_in[0]
+ cbx_2__4_/chanx_left_in[10] cbx_2__4_/chanx_left_in[11] cbx_2__4_/chanx_left_in[12]
+ cbx_2__4_/chanx_left_in[13] cbx_2__4_/chanx_left_in[14] cbx_2__4_/chanx_left_in[15]
+ cbx_2__4_/chanx_left_in[16] cbx_2__4_/chanx_left_in[17] cbx_2__4_/chanx_left_in[18]
+ cbx_2__4_/chanx_left_in[19] cbx_2__4_/chanx_left_in[1] cbx_2__4_/chanx_left_in[2]
+ cbx_2__4_/chanx_left_in[3] cbx_2__4_/chanx_left_in[4] cbx_2__4_/chanx_left_in[5]
+ cbx_2__4_/chanx_left_in[6] cbx_2__4_/chanx_left_in[7] cbx_2__4_/chanx_left_in[8]
+ cbx_2__4_/chanx_left_in[9] cby_1__4_/chany_top_out[0] cby_1__4_/chany_top_out[10]
+ cby_1__4_/chany_top_out[11] cby_1__4_/chany_top_out[12] cby_1__4_/chany_top_out[13]
+ cby_1__4_/chany_top_out[14] cby_1__4_/chany_top_out[15] cby_1__4_/chany_top_out[16]
+ cby_1__4_/chany_top_out[17] cby_1__4_/chany_top_out[18] cby_1__4_/chany_top_out[19]
+ cby_1__4_/chany_top_out[1] cby_1__4_/chany_top_out[2] cby_1__4_/chany_top_out[3]
+ cby_1__4_/chany_top_out[4] cby_1__4_/chany_top_out[5] cby_1__4_/chany_top_out[6]
+ cby_1__4_/chany_top_out[7] cby_1__4_/chany_top_out[8] cby_1__4_/chany_top_out[9]
+ cby_1__4_/chany_top_in[0] cby_1__4_/chany_top_in[10] cby_1__4_/chany_top_in[11]
+ cby_1__4_/chany_top_in[12] cby_1__4_/chany_top_in[13] cby_1__4_/chany_top_in[14]
+ cby_1__4_/chany_top_in[15] cby_1__4_/chany_top_in[16] cby_1__4_/chany_top_in[17]
+ cby_1__4_/chany_top_in[18] cby_1__4_/chany_top_in[19] cby_1__4_/chany_top_in[1]
+ cby_1__4_/chany_top_in[2] cby_1__4_/chany_top_in[3] cby_1__4_/chany_top_in[4] cby_1__4_/chany_top_in[5]
+ cby_1__4_/chany_top_in[6] cby_1__4_/chany_top_in[7] cby_1__4_/chany_top_in[8] cby_1__4_/chany_top_in[9]
+ sb_1__4_/chany_top_in[0] sb_1__4_/chany_top_in[10] sb_1__4_/chany_top_in[11] sb_1__4_/chany_top_in[12]
+ sb_1__4_/chany_top_in[13] sb_1__4_/chany_top_in[14] sb_1__4_/chany_top_in[15] sb_1__4_/chany_top_in[16]
+ sb_1__4_/chany_top_in[17] sb_1__4_/chany_top_in[18] sb_1__4_/chany_top_in[19] sb_1__4_/chany_top_in[1]
+ sb_1__4_/chany_top_in[2] sb_1__4_/chany_top_in[3] sb_1__4_/chany_top_in[4] sb_1__4_/chany_top_in[5]
+ sb_1__4_/chany_top_in[6] sb_1__4_/chany_top_in[7] sb_1__4_/chany_top_in[8] sb_1__4_/chany_top_in[9]
+ sb_1__4_/chany_top_out[0] sb_1__4_/chany_top_out[10] sb_1__4_/chany_top_out[11]
+ sb_1__4_/chany_top_out[12] sb_1__4_/chany_top_out[13] sb_1__4_/chany_top_out[14]
+ sb_1__4_/chany_top_out[15] sb_1__4_/chany_top_out[16] sb_1__4_/chany_top_out[17]
+ sb_1__4_/chany_top_out[18] sb_1__4_/chany_top_out[19] sb_1__4_/chany_top_out[1]
+ sb_1__4_/chany_top_out[2] sb_1__4_/chany_top_out[3] sb_1__4_/chany_top_out[4] sb_1__4_/chany_top_out[5]
+ sb_1__4_/chany_top_out[6] sb_1__4_/chany_top_out[7] sb_1__4_/chany_top_out[8] sb_1__4_/chany_top_out[9]
+ sb_1__4_/clk_1_E_out sb_1__4_/clk_1_N_in sb_1__4_/clk_1_W_out sb_1__4_/clk_2_E_out
+ sb_1__4_/clk_2_N_in sb_1__4_/clk_2_N_out sb_1__4_/clk_2_S_out sb_1__4_/clk_2_W_out
+ sb_1__4_/clk_3_E_out sb_1__4_/clk_3_N_in sb_1__4_/clk_3_N_out sb_1__4_/clk_3_S_out
+ sb_1__4_/clk_3_W_out sb_1__4_/left_bottom_grid_pin_34_ sb_1__4_/left_bottom_grid_pin_35_
+ sb_1__4_/left_bottom_grid_pin_36_ sb_1__4_/left_bottom_grid_pin_37_ sb_1__4_/left_bottom_grid_pin_38_
+ sb_1__4_/left_bottom_grid_pin_39_ sb_1__4_/left_bottom_grid_pin_40_ sb_1__4_/left_bottom_grid_pin_41_
+ sb_1__4_/prog_clk_0_N_in sb_1__4_/prog_clk_1_E_out sb_1__4_/prog_clk_1_N_in sb_1__4_/prog_clk_1_W_out
+ sb_1__4_/prog_clk_2_E_out sb_1__4_/prog_clk_2_N_in sb_1__4_/prog_clk_2_N_out sb_1__4_/prog_clk_2_S_out
+ sb_1__4_/prog_clk_2_W_out sb_1__4_/prog_clk_3_E_out sb_1__4_/prog_clk_3_N_in sb_1__4_/prog_clk_3_N_out
+ sb_1__4_/prog_clk_3_S_out sb_1__4_/prog_clk_3_W_out sb_1__4_/right_bottom_grid_pin_34_
+ sb_1__4_/right_bottom_grid_pin_35_ sb_1__4_/right_bottom_grid_pin_36_ sb_1__4_/right_bottom_grid_pin_37_
+ sb_1__4_/right_bottom_grid_pin_38_ sb_1__4_/right_bottom_grid_pin_39_ sb_1__4_/right_bottom_grid_pin_40_
+ sb_1__4_/right_bottom_grid_pin_41_ sb_1__4_/top_left_grid_pin_42_ sb_1__4_/top_left_grid_pin_43_
+ sb_1__4_/top_left_grid_pin_44_ sb_1__4_/top_left_grid_pin_45_ sb_1__4_/top_left_grid_pin_46_
+ sb_1__4_/top_left_grid_pin_47_ sb_1__4_/top_left_grid_pin_48_ sb_1__4_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_7__3_ cby_7__3_/Test_en_W_in cby_7__3_/Test_en_E_out cby_7__3_/Test_en_N_out
+ cby_7__3_/Test_en_W_in cby_7__3_/Test_en_W_in cby_7__3_/Test_en_W_out VGND VPWR
+ cby_7__3_/ccff_head cby_7__3_/ccff_tail sb_7__2_/chany_top_out[0] sb_7__2_/chany_top_out[10]
+ sb_7__2_/chany_top_out[11] sb_7__2_/chany_top_out[12] sb_7__2_/chany_top_out[13]
+ sb_7__2_/chany_top_out[14] sb_7__2_/chany_top_out[15] sb_7__2_/chany_top_out[16]
+ sb_7__2_/chany_top_out[17] sb_7__2_/chany_top_out[18] sb_7__2_/chany_top_out[19]
+ sb_7__2_/chany_top_out[1] sb_7__2_/chany_top_out[2] sb_7__2_/chany_top_out[3] sb_7__2_/chany_top_out[4]
+ sb_7__2_/chany_top_out[5] sb_7__2_/chany_top_out[6] sb_7__2_/chany_top_out[7] sb_7__2_/chany_top_out[8]
+ sb_7__2_/chany_top_out[9] sb_7__2_/chany_top_in[0] sb_7__2_/chany_top_in[10] sb_7__2_/chany_top_in[11]
+ sb_7__2_/chany_top_in[12] sb_7__2_/chany_top_in[13] sb_7__2_/chany_top_in[14] sb_7__2_/chany_top_in[15]
+ sb_7__2_/chany_top_in[16] sb_7__2_/chany_top_in[17] sb_7__2_/chany_top_in[18] sb_7__2_/chany_top_in[19]
+ sb_7__2_/chany_top_in[1] sb_7__2_/chany_top_in[2] sb_7__2_/chany_top_in[3] sb_7__2_/chany_top_in[4]
+ sb_7__2_/chany_top_in[5] sb_7__2_/chany_top_in[6] sb_7__2_/chany_top_in[7] sb_7__2_/chany_top_in[8]
+ sb_7__2_/chany_top_in[9] cby_7__3_/chany_top_in[0] cby_7__3_/chany_top_in[10] cby_7__3_/chany_top_in[11]
+ cby_7__3_/chany_top_in[12] cby_7__3_/chany_top_in[13] cby_7__3_/chany_top_in[14]
+ cby_7__3_/chany_top_in[15] cby_7__3_/chany_top_in[16] cby_7__3_/chany_top_in[17]
+ cby_7__3_/chany_top_in[18] cby_7__3_/chany_top_in[19] cby_7__3_/chany_top_in[1]
+ cby_7__3_/chany_top_in[2] cby_7__3_/chany_top_in[3] cby_7__3_/chany_top_in[4] cby_7__3_/chany_top_in[5]
+ cby_7__3_/chany_top_in[6] cby_7__3_/chany_top_in[7] cby_7__3_/chany_top_in[8] cby_7__3_/chany_top_in[9]
+ cby_7__3_/chany_top_out[0] cby_7__3_/chany_top_out[10] cby_7__3_/chany_top_out[11]
+ cby_7__3_/chany_top_out[12] cby_7__3_/chany_top_out[13] cby_7__3_/chany_top_out[14]
+ cby_7__3_/chany_top_out[15] cby_7__3_/chany_top_out[16] cby_7__3_/chany_top_out[17]
+ cby_7__3_/chany_top_out[18] cby_7__3_/chany_top_out[19] cby_7__3_/chany_top_out[1]
+ cby_7__3_/chany_top_out[2] cby_7__3_/chany_top_out[3] cby_7__3_/chany_top_out[4]
+ cby_7__3_/chany_top_out[5] cby_7__3_/chany_top_out[6] cby_7__3_/chany_top_out[7]
+ cby_7__3_/chany_top_out[8] cby_7__3_/chany_top_out[9] sb_7__3_/clk_1_N_in sb_7__2_/clk_2_N_out
+ cby_7__3_/clk_2_S_out cby_7__3_/clk_3_N_out cby_7__3_/clk_3_S_in cby_7__3_/clk_3_S_out
+ cby_7__3_/left_grid_pin_16_ cby_7__3_/left_grid_pin_17_ cby_7__3_/left_grid_pin_18_
+ cby_7__3_/left_grid_pin_19_ cby_7__3_/left_grid_pin_20_ cby_7__3_/left_grid_pin_21_
+ cby_7__3_/left_grid_pin_22_ cby_7__3_/left_grid_pin_23_ cby_7__3_/left_grid_pin_24_
+ cby_7__3_/left_grid_pin_25_ cby_7__3_/left_grid_pin_26_ cby_7__3_/left_grid_pin_27_
+ cby_7__3_/left_grid_pin_28_ cby_7__3_/left_grid_pin_29_ cby_7__3_/left_grid_pin_30_
+ cby_7__3_/left_grid_pin_31_ cby_7__3_/prog_clk_0_N_out sb_7__2_/prog_clk_0_N_in
+ cby_7__3_/prog_clk_0_W_in sb_7__3_/prog_clk_1_N_in sb_7__2_/prog_clk_2_N_out cby_7__3_/prog_clk_2_S_out
+ cby_7__3_/prog_clk_3_N_out cby_7__3_/prog_clk_3_S_in cby_7__3_/prog_clk_3_S_out
+ cby_1__1_
Xcby_0__8_ IO_ISOL_N VGND VPWR sb_0__8_/ccff_tail cby_0__8_/ccff_tail sb_0__7_/chany_top_out[0]
+ sb_0__7_/chany_top_out[10] sb_0__7_/chany_top_out[11] sb_0__7_/chany_top_out[12]
+ sb_0__7_/chany_top_out[13] sb_0__7_/chany_top_out[14] sb_0__7_/chany_top_out[15]
+ sb_0__7_/chany_top_out[16] sb_0__7_/chany_top_out[17] sb_0__7_/chany_top_out[18]
+ sb_0__7_/chany_top_out[19] sb_0__7_/chany_top_out[1] sb_0__7_/chany_top_out[2] sb_0__7_/chany_top_out[3]
+ sb_0__7_/chany_top_out[4] sb_0__7_/chany_top_out[5] sb_0__7_/chany_top_out[6] sb_0__7_/chany_top_out[7]
+ sb_0__7_/chany_top_out[8] sb_0__7_/chany_top_out[9] sb_0__7_/chany_top_in[0] sb_0__7_/chany_top_in[10]
+ sb_0__7_/chany_top_in[11] sb_0__7_/chany_top_in[12] sb_0__7_/chany_top_in[13] sb_0__7_/chany_top_in[14]
+ sb_0__7_/chany_top_in[15] sb_0__7_/chany_top_in[16] sb_0__7_/chany_top_in[17] sb_0__7_/chany_top_in[18]
+ sb_0__7_/chany_top_in[19] sb_0__7_/chany_top_in[1] sb_0__7_/chany_top_in[2] sb_0__7_/chany_top_in[3]
+ sb_0__7_/chany_top_in[4] sb_0__7_/chany_top_in[5] sb_0__7_/chany_top_in[6] sb_0__7_/chany_top_in[7]
+ sb_0__7_/chany_top_in[8] sb_0__7_/chany_top_in[9] cby_0__8_/chany_top_in[0] cby_0__8_/chany_top_in[10]
+ cby_0__8_/chany_top_in[11] cby_0__8_/chany_top_in[12] cby_0__8_/chany_top_in[13]
+ cby_0__8_/chany_top_in[14] cby_0__8_/chany_top_in[15] cby_0__8_/chany_top_in[16]
+ cby_0__8_/chany_top_in[17] cby_0__8_/chany_top_in[18] cby_0__8_/chany_top_in[19]
+ cby_0__8_/chany_top_in[1] cby_0__8_/chany_top_in[2] cby_0__8_/chany_top_in[3] cby_0__8_/chany_top_in[4]
+ cby_0__8_/chany_top_in[5] cby_0__8_/chany_top_in[6] cby_0__8_/chany_top_in[7] cby_0__8_/chany_top_in[8]
+ cby_0__8_/chany_top_in[9] cby_0__8_/chany_top_out[0] cby_0__8_/chany_top_out[10]
+ cby_0__8_/chany_top_out[11] cby_0__8_/chany_top_out[12] cby_0__8_/chany_top_out[13]
+ cby_0__8_/chany_top_out[14] cby_0__8_/chany_top_out[15] cby_0__8_/chany_top_out[16]
+ cby_0__8_/chany_top_out[17] cby_0__8_/chany_top_out[18] cby_0__8_/chany_top_out[19]
+ cby_0__8_/chany_top_out[1] cby_0__8_/chany_top_out[2] cby_0__8_/chany_top_out[3]
+ cby_0__8_/chany_top_out[4] cby_0__8_/chany_top_out[5] cby_0__8_/chany_top_out[6]
+ cby_0__8_/chany_top_out[7] cby_0__8_/chany_top_out[8] cby_0__8_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
+ cby_0__8_/left_grid_pin_0_ cby_0__8_/prog_clk_0_E_in cby_0__8_/left_grid_pin_0_
+ sb_0__7_/top_left_grid_pin_1_ sb_0__8_/bottom_left_grid_pin_1_ cby_0__1_
Xcbx_7__4_ cbx_7__4_/REGIN_FEEDTHROUGH cbx_7__4_/REGOUT_FEEDTHROUGH cbx_7__4_/SC_IN_BOT
+ cbx_7__4_/SC_IN_TOP cbx_7__4_/SC_OUT_BOT cbx_7__4_/SC_OUT_TOP VGND VPWR cbx_7__4_/bottom_grid_pin_0_
+ cbx_7__4_/bottom_grid_pin_10_ cbx_7__4_/bottom_grid_pin_11_ cbx_7__4_/bottom_grid_pin_12_
+ cbx_7__4_/bottom_grid_pin_13_ cbx_7__4_/bottom_grid_pin_14_ cbx_7__4_/bottom_grid_pin_15_
+ cbx_7__4_/bottom_grid_pin_1_ cbx_7__4_/bottom_grid_pin_2_ cbx_7__4_/bottom_grid_pin_3_
+ cbx_7__4_/bottom_grid_pin_4_ cbx_7__4_/bottom_grid_pin_5_ cbx_7__4_/bottom_grid_pin_6_
+ cbx_7__4_/bottom_grid_pin_7_ cbx_7__4_/bottom_grid_pin_8_ cbx_7__4_/bottom_grid_pin_9_
+ sb_7__4_/ccff_tail sb_6__4_/ccff_head cbx_7__4_/chanx_left_in[0] cbx_7__4_/chanx_left_in[10]
+ cbx_7__4_/chanx_left_in[11] cbx_7__4_/chanx_left_in[12] cbx_7__4_/chanx_left_in[13]
+ cbx_7__4_/chanx_left_in[14] cbx_7__4_/chanx_left_in[15] cbx_7__4_/chanx_left_in[16]
+ cbx_7__4_/chanx_left_in[17] cbx_7__4_/chanx_left_in[18] cbx_7__4_/chanx_left_in[19]
+ cbx_7__4_/chanx_left_in[1] cbx_7__4_/chanx_left_in[2] cbx_7__4_/chanx_left_in[3]
+ cbx_7__4_/chanx_left_in[4] cbx_7__4_/chanx_left_in[5] cbx_7__4_/chanx_left_in[6]
+ cbx_7__4_/chanx_left_in[7] cbx_7__4_/chanx_left_in[8] cbx_7__4_/chanx_left_in[9]
+ sb_6__4_/chanx_right_in[0] sb_6__4_/chanx_right_in[10] sb_6__4_/chanx_right_in[11]
+ sb_6__4_/chanx_right_in[12] sb_6__4_/chanx_right_in[13] sb_6__4_/chanx_right_in[14]
+ sb_6__4_/chanx_right_in[15] sb_6__4_/chanx_right_in[16] sb_6__4_/chanx_right_in[17]
+ sb_6__4_/chanx_right_in[18] sb_6__4_/chanx_right_in[19] sb_6__4_/chanx_right_in[1]
+ sb_6__4_/chanx_right_in[2] sb_6__4_/chanx_right_in[3] sb_6__4_/chanx_right_in[4]
+ sb_6__4_/chanx_right_in[5] sb_6__4_/chanx_right_in[6] sb_6__4_/chanx_right_in[7]
+ sb_6__4_/chanx_right_in[8] sb_6__4_/chanx_right_in[9] sb_7__4_/chanx_left_out[0]
+ sb_7__4_/chanx_left_out[10] sb_7__4_/chanx_left_out[11] sb_7__4_/chanx_left_out[12]
+ sb_7__4_/chanx_left_out[13] sb_7__4_/chanx_left_out[14] sb_7__4_/chanx_left_out[15]
+ sb_7__4_/chanx_left_out[16] sb_7__4_/chanx_left_out[17] sb_7__4_/chanx_left_out[18]
+ sb_7__4_/chanx_left_out[19] sb_7__4_/chanx_left_out[1] sb_7__4_/chanx_left_out[2]
+ sb_7__4_/chanx_left_out[3] sb_7__4_/chanx_left_out[4] sb_7__4_/chanx_left_out[5]
+ sb_7__4_/chanx_left_out[6] sb_7__4_/chanx_left_out[7] sb_7__4_/chanx_left_out[8]
+ sb_7__4_/chanx_left_out[9] sb_7__4_/chanx_left_in[0] sb_7__4_/chanx_left_in[10]
+ sb_7__4_/chanx_left_in[11] sb_7__4_/chanx_left_in[12] sb_7__4_/chanx_left_in[13]
+ sb_7__4_/chanx_left_in[14] sb_7__4_/chanx_left_in[15] sb_7__4_/chanx_left_in[16]
+ sb_7__4_/chanx_left_in[17] sb_7__4_/chanx_left_in[18] sb_7__4_/chanx_left_in[19]
+ sb_7__4_/chanx_left_in[1] sb_7__4_/chanx_left_in[2] sb_7__4_/chanx_left_in[3] sb_7__4_/chanx_left_in[4]
+ sb_7__4_/chanx_left_in[5] sb_7__4_/chanx_left_in[6] sb_7__4_/chanx_left_in[7] sb_7__4_/chanx_left_in[8]
+ sb_7__4_/chanx_left_in[9] cbx_7__4_/clk_1_N_out cbx_7__4_/clk_1_S_out cbx_7__4_/clk_1_W_in
+ cbx_7__4_/clk_2_E_out cbx_7__4_/clk_2_W_in cbx_7__4_/clk_2_W_out cbx_7__4_/clk_3_E_out
+ cbx_7__4_/clk_3_W_in cbx_7__4_/clk_3_W_out cbx_7__4_/prog_clk_0_N_in cbx_7__4_/prog_clk_0_W_out
+ cbx_7__4_/prog_clk_1_N_out cbx_7__4_/prog_clk_1_S_out cbx_7__4_/prog_clk_1_W_in
+ cbx_7__4_/prog_clk_2_E_out cbx_7__4_/prog_clk_2_W_in cbx_7__4_/prog_clk_2_W_out
+ cbx_7__4_/prog_clk_3_E_out cbx_7__4_/prog_clk_3_W_in cbx_7__4_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_6__4_ cbx_6__3_/SC_OUT_TOP grid_clb_6__4_/SC_OUT_BOT cbx_6__4_/SC_IN_BOT
+ cby_5__4_/Test_en_E_out cby_6__4_/Test_en_W_in cby_5__4_/Test_en_E_out grid_clb_6__4_/Test_en_W_out
+ VGND VPWR cbx_6__3_/REGIN_FEEDTHROUGH grid_clb_6__4_/bottom_width_0_height_0__pin_51_
+ cby_5__4_/ccff_tail cby_6__4_/ccff_head cbx_6__3_/clk_1_N_out cbx_6__3_/clk_1_N_out
+ cby_6__4_/prog_clk_0_W_in cbx_6__3_/prog_clk_1_N_out grid_clb_6__4_/prog_clk_0_N_out
+ cbx_6__3_/prog_clk_1_N_out cbx_6__3_/prog_clk_0_N_in grid_clb_6__4_/prog_clk_0_W_out
+ cby_6__4_/left_grid_pin_16_ cby_6__4_/left_grid_pin_17_ cby_6__4_/left_grid_pin_18_
+ cby_6__4_/left_grid_pin_19_ cby_6__4_/left_grid_pin_20_ cby_6__4_/left_grid_pin_21_
+ cby_6__4_/left_grid_pin_22_ cby_6__4_/left_grid_pin_23_ cby_6__4_/left_grid_pin_24_
+ cby_6__4_/left_grid_pin_25_ cby_6__4_/left_grid_pin_26_ cby_6__4_/left_grid_pin_27_
+ cby_6__4_/left_grid_pin_28_ cby_6__4_/left_grid_pin_29_ cby_6__4_/left_grid_pin_30_
+ cby_6__4_/left_grid_pin_31_ sb_6__3_/top_left_grid_pin_42_ sb_6__4_/bottom_left_grid_pin_42_
+ sb_6__3_/top_left_grid_pin_43_ sb_6__4_/bottom_left_grid_pin_43_ sb_6__3_/top_left_grid_pin_44_
+ sb_6__4_/bottom_left_grid_pin_44_ sb_6__3_/top_left_grid_pin_45_ sb_6__4_/bottom_left_grid_pin_45_
+ sb_6__3_/top_left_grid_pin_46_ sb_6__4_/bottom_left_grid_pin_46_ sb_6__3_/top_left_grid_pin_47_
+ sb_6__4_/bottom_left_grid_pin_47_ sb_6__3_/top_left_grid_pin_48_ sb_6__4_/bottom_left_grid_pin_48_
+ sb_6__3_/top_left_grid_pin_49_ sb_6__4_/bottom_left_grid_pin_49_ cbx_6__4_/bottom_grid_pin_0_
+ cbx_6__4_/bottom_grid_pin_10_ cbx_6__4_/bottom_grid_pin_11_ cbx_6__4_/bottom_grid_pin_12_
+ cbx_6__4_/bottom_grid_pin_13_ cbx_6__4_/bottom_grid_pin_14_ cbx_6__4_/bottom_grid_pin_15_
+ cbx_6__4_/bottom_grid_pin_1_ cbx_6__4_/bottom_grid_pin_2_ cbx_6__4_/REGOUT_FEEDTHROUGH
+ grid_clb_6__4_/top_width_0_height_0__pin_33_ sb_6__4_/left_bottom_grid_pin_34_ sb_5__4_/right_bottom_grid_pin_34_
+ sb_6__4_/left_bottom_grid_pin_35_ sb_5__4_/right_bottom_grid_pin_35_ sb_6__4_/left_bottom_grid_pin_36_
+ sb_5__4_/right_bottom_grid_pin_36_ sb_6__4_/left_bottom_grid_pin_37_ sb_5__4_/right_bottom_grid_pin_37_
+ sb_6__4_/left_bottom_grid_pin_38_ sb_5__4_/right_bottom_grid_pin_38_ sb_6__4_/left_bottom_grid_pin_39_
+ sb_5__4_/right_bottom_grid_pin_39_ cbx_6__4_/bottom_grid_pin_3_ sb_6__4_/left_bottom_grid_pin_40_
+ sb_5__4_/right_bottom_grid_pin_40_ sb_6__4_/left_bottom_grid_pin_41_ sb_5__4_/right_bottom_grid_pin_41_
+ cbx_6__4_/bottom_grid_pin_4_ cbx_6__4_/bottom_grid_pin_5_ cbx_6__4_/bottom_grid_pin_6_
+ cbx_6__4_/bottom_grid_pin_7_ cbx_6__4_/bottom_grid_pin_8_ cbx_6__4_/bottom_grid_pin_9_
+ grid_clb
Xcbx_4__1_ cbx_4__1_/REGIN_FEEDTHROUGH cbx_4__1_/REGOUT_FEEDTHROUGH cbx_4__1_/SC_IN_BOT
+ cbx_4__1_/SC_IN_TOP cbx_4__1_/SC_OUT_BOT cbx_4__1_/SC_OUT_TOP VGND VPWR cbx_4__1_/bottom_grid_pin_0_
+ cbx_4__1_/bottom_grid_pin_10_ cbx_4__1_/bottom_grid_pin_11_ cbx_4__1_/bottom_grid_pin_12_
+ cbx_4__1_/bottom_grid_pin_13_ cbx_4__1_/bottom_grid_pin_14_ cbx_4__1_/bottom_grid_pin_15_
+ cbx_4__1_/bottom_grid_pin_1_ cbx_4__1_/bottom_grid_pin_2_ cbx_4__1_/bottom_grid_pin_3_
+ cbx_4__1_/bottom_grid_pin_4_ cbx_4__1_/bottom_grid_pin_5_ cbx_4__1_/bottom_grid_pin_6_
+ cbx_4__1_/bottom_grid_pin_7_ cbx_4__1_/bottom_grid_pin_8_ cbx_4__1_/bottom_grid_pin_9_
+ sb_4__1_/ccff_tail sb_3__1_/ccff_head cbx_4__1_/chanx_left_in[0] cbx_4__1_/chanx_left_in[10]
+ cbx_4__1_/chanx_left_in[11] cbx_4__1_/chanx_left_in[12] cbx_4__1_/chanx_left_in[13]
+ cbx_4__1_/chanx_left_in[14] cbx_4__1_/chanx_left_in[15] cbx_4__1_/chanx_left_in[16]
+ cbx_4__1_/chanx_left_in[17] cbx_4__1_/chanx_left_in[18] cbx_4__1_/chanx_left_in[19]
+ cbx_4__1_/chanx_left_in[1] cbx_4__1_/chanx_left_in[2] cbx_4__1_/chanx_left_in[3]
+ cbx_4__1_/chanx_left_in[4] cbx_4__1_/chanx_left_in[5] cbx_4__1_/chanx_left_in[6]
+ cbx_4__1_/chanx_left_in[7] cbx_4__1_/chanx_left_in[8] cbx_4__1_/chanx_left_in[9]
+ sb_3__1_/chanx_right_in[0] sb_3__1_/chanx_right_in[10] sb_3__1_/chanx_right_in[11]
+ sb_3__1_/chanx_right_in[12] sb_3__1_/chanx_right_in[13] sb_3__1_/chanx_right_in[14]
+ sb_3__1_/chanx_right_in[15] sb_3__1_/chanx_right_in[16] sb_3__1_/chanx_right_in[17]
+ sb_3__1_/chanx_right_in[18] sb_3__1_/chanx_right_in[19] sb_3__1_/chanx_right_in[1]
+ sb_3__1_/chanx_right_in[2] sb_3__1_/chanx_right_in[3] sb_3__1_/chanx_right_in[4]
+ sb_3__1_/chanx_right_in[5] sb_3__1_/chanx_right_in[6] sb_3__1_/chanx_right_in[7]
+ sb_3__1_/chanx_right_in[8] sb_3__1_/chanx_right_in[9] sb_4__1_/chanx_left_out[0]
+ sb_4__1_/chanx_left_out[10] sb_4__1_/chanx_left_out[11] sb_4__1_/chanx_left_out[12]
+ sb_4__1_/chanx_left_out[13] sb_4__1_/chanx_left_out[14] sb_4__1_/chanx_left_out[15]
+ sb_4__1_/chanx_left_out[16] sb_4__1_/chanx_left_out[17] sb_4__1_/chanx_left_out[18]
+ sb_4__1_/chanx_left_out[19] sb_4__1_/chanx_left_out[1] sb_4__1_/chanx_left_out[2]
+ sb_4__1_/chanx_left_out[3] sb_4__1_/chanx_left_out[4] sb_4__1_/chanx_left_out[5]
+ sb_4__1_/chanx_left_out[6] sb_4__1_/chanx_left_out[7] sb_4__1_/chanx_left_out[8]
+ sb_4__1_/chanx_left_out[9] sb_4__1_/chanx_left_in[0] sb_4__1_/chanx_left_in[10]
+ sb_4__1_/chanx_left_in[11] sb_4__1_/chanx_left_in[12] sb_4__1_/chanx_left_in[13]
+ sb_4__1_/chanx_left_in[14] sb_4__1_/chanx_left_in[15] sb_4__1_/chanx_left_in[16]
+ sb_4__1_/chanx_left_in[17] sb_4__1_/chanx_left_in[18] sb_4__1_/chanx_left_in[19]
+ sb_4__1_/chanx_left_in[1] sb_4__1_/chanx_left_in[2] sb_4__1_/chanx_left_in[3] sb_4__1_/chanx_left_in[4]
+ sb_4__1_/chanx_left_in[5] sb_4__1_/chanx_left_in[6] sb_4__1_/chanx_left_in[7] sb_4__1_/chanx_left_in[8]
+ sb_4__1_/chanx_left_in[9] cbx_4__1_/clk_1_N_out cbx_4__1_/clk_1_S_out sb_3__1_/clk_1_E_out
+ cbx_4__1_/clk_2_E_out cbx_4__1_/clk_2_W_in cbx_4__1_/clk_2_W_out cbx_4__1_/clk_3_E_out
+ cbx_4__1_/clk_3_W_in cbx_4__1_/clk_3_W_out cbx_4__1_/prog_clk_0_N_in cbx_4__1_/prog_clk_0_W_out
+ cbx_4__1_/prog_clk_1_N_out cbx_4__1_/prog_clk_1_S_out sb_3__1_/prog_clk_1_E_out
+ cbx_4__1_/prog_clk_2_E_out cbx_4__1_/prog_clk_2_W_in cbx_4__1_/prog_clk_2_W_out
+ cbx_4__1_/prog_clk_3_E_out cbx_4__1_/prog_clk_3_W_in cbx_4__1_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_4__6_ sb_4__6_/Test_en_N_out sb_4__6_/Test_en_S_in VGND VPWR sb_4__6_/bottom_left_grid_pin_42_
+ sb_4__6_/bottom_left_grid_pin_43_ sb_4__6_/bottom_left_grid_pin_44_ sb_4__6_/bottom_left_grid_pin_45_
+ sb_4__6_/bottom_left_grid_pin_46_ sb_4__6_/bottom_left_grid_pin_47_ sb_4__6_/bottom_left_grid_pin_48_
+ sb_4__6_/bottom_left_grid_pin_49_ sb_4__6_/ccff_head sb_4__6_/ccff_tail sb_4__6_/chanx_left_in[0]
+ sb_4__6_/chanx_left_in[10] sb_4__6_/chanx_left_in[11] sb_4__6_/chanx_left_in[12]
+ sb_4__6_/chanx_left_in[13] sb_4__6_/chanx_left_in[14] sb_4__6_/chanx_left_in[15]
+ sb_4__6_/chanx_left_in[16] sb_4__6_/chanx_left_in[17] sb_4__6_/chanx_left_in[18]
+ sb_4__6_/chanx_left_in[19] sb_4__6_/chanx_left_in[1] sb_4__6_/chanx_left_in[2] sb_4__6_/chanx_left_in[3]
+ sb_4__6_/chanx_left_in[4] sb_4__6_/chanx_left_in[5] sb_4__6_/chanx_left_in[6] sb_4__6_/chanx_left_in[7]
+ sb_4__6_/chanx_left_in[8] sb_4__6_/chanx_left_in[9] sb_4__6_/chanx_left_out[0] sb_4__6_/chanx_left_out[10]
+ sb_4__6_/chanx_left_out[11] sb_4__6_/chanx_left_out[12] sb_4__6_/chanx_left_out[13]
+ sb_4__6_/chanx_left_out[14] sb_4__6_/chanx_left_out[15] sb_4__6_/chanx_left_out[16]
+ sb_4__6_/chanx_left_out[17] sb_4__6_/chanx_left_out[18] sb_4__6_/chanx_left_out[19]
+ sb_4__6_/chanx_left_out[1] sb_4__6_/chanx_left_out[2] sb_4__6_/chanx_left_out[3]
+ sb_4__6_/chanx_left_out[4] sb_4__6_/chanx_left_out[5] sb_4__6_/chanx_left_out[6]
+ sb_4__6_/chanx_left_out[7] sb_4__6_/chanx_left_out[8] sb_4__6_/chanx_left_out[9]
+ sb_4__6_/chanx_right_in[0] sb_4__6_/chanx_right_in[10] sb_4__6_/chanx_right_in[11]
+ sb_4__6_/chanx_right_in[12] sb_4__6_/chanx_right_in[13] sb_4__6_/chanx_right_in[14]
+ sb_4__6_/chanx_right_in[15] sb_4__6_/chanx_right_in[16] sb_4__6_/chanx_right_in[17]
+ sb_4__6_/chanx_right_in[18] sb_4__6_/chanx_right_in[19] sb_4__6_/chanx_right_in[1]
+ sb_4__6_/chanx_right_in[2] sb_4__6_/chanx_right_in[3] sb_4__6_/chanx_right_in[4]
+ sb_4__6_/chanx_right_in[5] sb_4__6_/chanx_right_in[6] sb_4__6_/chanx_right_in[7]
+ sb_4__6_/chanx_right_in[8] sb_4__6_/chanx_right_in[9] cbx_5__6_/chanx_left_in[0]
+ cbx_5__6_/chanx_left_in[10] cbx_5__6_/chanx_left_in[11] cbx_5__6_/chanx_left_in[12]
+ cbx_5__6_/chanx_left_in[13] cbx_5__6_/chanx_left_in[14] cbx_5__6_/chanx_left_in[15]
+ cbx_5__6_/chanx_left_in[16] cbx_5__6_/chanx_left_in[17] cbx_5__6_/chanx_left_in[18]
+ cbx_5__6_/chanx_left_in[19] cbx_5__6_/chanx_left_in[1] cbx_5__6_/chanx_left_in[2]
+ cbx_5__6_/chanx_left_in[3] cbx_5__6_/chanx_left_in[4] cbx_5__6_/chanx_left_in[5]
+ cbx_5__6_/chanx_left_in[6] cbx_5__6_/chanx_left_in[7] cbx_5__6_/chanx_left_in[8]
+ cbx_5__6_/chanx_left_in[9] cby_4__6_/chany_top_out[0] cby_4__6_/chany_top_out[10]
+ cby_4__6_/chany_top_out[11] cby_4__6_/chany_top_out[12] cby_4__6_/chany_top_out[13]
+ cby_4__6_/chany_top_out[14] cby_4__6_/chany_top_out[15] cby_4__6_/chany_top_out[16]
+ cby_4__6_/chany_top_out[17] cby_4__6_/chany_top_out[18] cby_4__6_/chany_top_out[19]
+ cby_4__6_/chany_top_out[1] cby_4__6_/chany_top_out[2] cby_4__6_/chany_top_out[3]
+ cby_4__6_/chany_top_out[4] cby_4__6_/chany_top_out[5] cby_4__6_/chany_top_out[6]
+ cby_4__6_/chany_top_out[7] cby_4__6_/chany_top_out[8] cby_4__6_/chany_top_out[9]
+ cby_4__6_/chany_top_in[0] cby_4__6_/chany_top_in[10] cby_4__6_/chany_top_in[11]
+ cby_4__6_/chany_top_in[12] cby_4__6_/chany_top_in[13] cby_4__6_/chany_top_in[14]
+ cby_4__6_/chany_top_in[15] cby_4__6_/chany_top_in[16] cby_4__6_/chany_top_in[17]
+ cby_4__6_/chany_top_in[18] cby_4__6_/chany_top_in[19] cby_4__6_/chany_top_in[1]
+ cby_4__6_/chany_top_in[2] cby_4__6_/chany_top_in[3] cby_4__6_/chany_top_in[4] cby_4__6_/chany_top_in[5]
+ cby_4__6_/chany_top_in[6] cby_4__6_/chany_top_in[7] cby_4__6_/chany_top_in[8] cby_4__6_/chany_top_in[9]
+ sb_4__6_/chany_top_in[0] sb_4__6_/chany_top_in[10] sb_4__6_/chany_top_in[11] sb_4__6_/chany_top_in[12]
+ sb_4__6_/chany_top_in[13] sb_4__6_/chany_top_in[14] sb_4__6_/chany_top_in[15] sb_4__6_/chany_top_in[16]
+ sb_4__6_/chany_top_in[17] sb_4__6_/chany_top_in[18] sb_4__6_/chany_top_in[19] sb_4__6_/chany_top_in[1]
+ sb_4__6_/chany_top_in[2] sb_4__6_/chany_top_in[3] sb_4__6_/chany_top_in[4] sb_4__6_/chany_top_in[5]
+ sb_4__6_/chany_top_in[6] sb_4__6_/chany_top_in[7] sb_4__6_/chany_top_in[8] sb_4__6_/chany_top_in[9]
+ sb_4__6_/chany_top_out[0] sb_4__6_/chany_top_out[10] sb_4__6_/chany_top_out[11]
+ sb_4__6_/chany_top_out[12] sb_4__6_/chany_top_out[13] sb_4__6_/chany_top_out[14]
+ sb_4__6_/chany_top_out[15] sb_4__6_/chany_top_out[16] sb_4__6_/chany_top_out[17]
+ sb_4__6_/chany_top_out[18] sb_4__6_/chany_top_out[19] sb_4__6_/chany_top_out[1]
+ sb_4__6_/chany_top_out[2] sb_4__6_/chany_top_out[3] sb_4__6_/chany_top_out[4] sb_4__6_/chany_top_out[5]
+ sb_4__6_/chany_top_out[6] sb_4__6_/chany_top_out[7] sb_4__6_/chany_top_out[8] sb_4__6_/chany_top_out[9]
+ sb_4__6_/clk_1_E_out sb_4__6_/clk_1_N_in sb_4__6_/clk_1_W_out sb_4__6_/clk_2_E_out
+ sb_4__6_/clk_2_N_in sb_4__6_/clk_2_N_out sb_4__6_/clk_2_S_out sb_4__6_/clk_2_W_out
+ sb_4__6_/clk_3_E_out sb_4__6_/clk_3_N_in sb_4__6_/clk_3_N_out sb_4__6_/clk_3_S_out
+ sb_4__6_/clk_3_W_out sb_4__6_/left_bottom_grid_pin_34_ sb_4__6_/left_bottom_grid_pin_35_
+ sb_4__6_/left_bottom_grid_pin_36_ sb_4__6_/left_bottom_grid_pin_37_ sb_4__6_/left_bottom_grid_pin_38_
+ sb_4__6_/left_bottom_grid_pin_39_ sb_4__6_/left_bottom_grid_pin_40_ sb_4__6_/left_bottom_grid_pin_41_
+ sb_4__6_/prog_clk_0_N_in sb_4__6_/prog_clk_1_E_out sb_4__6_/prog_clk_1_N_in sb_4__6_/prog_clk_1_W_out
+ sb_4__6_/prog_clk_2_E_out sb_4__6_/prog_clk_2_N_in sb_4__6_/prog_clk_2_N_out sb_4__6_/prog_clk_2_S_out
+ sb_4__6_/prog_clk_2_W_out sb_4__6_/prog_clk_3_E_out sb_4__6_/prog_clk_3_N_in sb_4__6_/prog_clk_3_N_out
+ sb_4__6_/prog_clk_3_S_out sb_4__6_/prog_clk_3_W_out sb_4__6_/right_bottom_grid_pin_34_
+ sb_4__6_/right_bottom_grid_pin_35_ sb_4__6_/right_bottom_grid_pin_36_ sb_4__6_/right_bottom_grid_pin_37_
+ sb_4__6_/right_bottom_grid_pin_38_ sb_4__6_/right_bottom_grid_pin_39_ sb_4__6_/right_bottom_grid_pin_40_
+ sb_4__6_/right_bottom_grid_pin_41_ sb_4__6_/top_left_grid_pin_42_ sb_4__6_/top_left_grid_pin_43_
+ sb_4__6_/top_left_grid_pin_44_ sb_4__6_/top_left_grid_pin_45_ sb_4__6_/top_left_grid_pin_46_
+ sb_4__6_/top_left_grid_pin_47_ sb_4__6_/top_left_grid_pin_48_ sb_4__6_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_1__3_ sb_1__3_/Test_en_N_out sb_1__3_/Test_en_S_in VGND VPWR sb_1__3_/bottom_left_grid_pin_42_
+ sb_1__3_/bottom_left_grid_pin_43_ sb_1__3_/bottom_left_grid_pin_44_ sb_1__3_/bottom_left_grid_pin_45_
+ sb_1__3_/bottom_left_grid_pin_46_ sb_1__3_/bottom_left_grid_pin_47_ sb_1__3_/bottom_left_grid_pin_48_
+ sb_1__3_/bottom_left_grid_pin_49_ sb_1__3_/ccff_head sb_1__3_/ccff_tail sb_1__3_/chanx_left_in[0]
+ sb_1__3_/chanx_left_in[10] sb_1__3_/chanx_left_in[11] sb_1__3_/chanx_left_in[12]
+ sb_1__3_/chanx_left_in[13] sb_1__3_/chanx_left_in[14] sb_1__3_/chanx_left_in[15]
+ sb_1__3_/chanx_left_in[16] sb_1__3_/chanx_left_in[17] sb_1__3_/chanx_left_in[18]
+ sb_1__3_/chanx_left_in[19] sb_1__3_/chanx_left_in[1] sb_1__3_/chanx_left_in[2] sb_1__3_/chanx_left_in[3]
+ sb_1__3_/chanx_left_in[4] sb_1__3_/chanx_left_in[5] sb_1__3_/chanx_left_in[6] sb_1__3_/chanx_left_in[7]
+ sb_1__3_/chanx_left_in[8] sb_1__3_/chanx_left_in[9] sb_1__3_/chanx_left_out[0] sb_1__3_/chanx_left_out[10]
+ sb_1__3_/chanx_left_out[11] sb_1__3_/chanx_left_out[12] sb_1__3_/chanx_left_out[13]
+ sb_1__3_/chanx_left_out[14] sb_1__3_/chanx_left_out[15] sb_1__3_/chanx_left_out[16]
+ sb_1__3_/chanx_left_out[17] sb_1__3_/chanx_left_out[18] sb_1__3_/chanx_left_out[19]
+ sb_1__3_/chanx_left_out[1] sb_1__3_/chanx_left_out[2] sb_1__3_/chanx_left_out[3]
+ sb_1__3_/chanx_left_out[4] sb_1__3_/chanx_left_out[5] sb_1__3_/chanx_left_out[6]
+ sb_1__3_/chanx_left_out[7] sb_1__3_/chanx_left_out[8] sb_1__3_/chanx_left_out[9]
+ sb_1__3_/chanx_right_in[0] sb_1__3_/chanx_right_in[10] sb_1__3_/chanx_right_in[11]
+ sb_1__3_/chanx_right_in[12] sb_1__3_/chanx_right_in[13] sb_1__3_/chanx_right_in[14]
+ sb_1__3_/chanx_right_in[15] sb_1__3_/chanx_right_in[16] sb_1__3_/chanx_right_in[17]
+ sb_1__3_/chanx_right_in[18] sb_1__3_/chanx_right_in[19] sb_1__3_/chanx_right_in[1]
+ sb_1__3_/chanx_right_in[2] sb_1__3_/chanx_right_in[3] sb_1__3_/chanx_right_in[4]
+ sb_1__3_/chanx_right_in[5] sb_1__3_/chanx_right_in[6] sb_1__3_/chanx_right_in[7]
+ sb_1__3_/chanx_right_in[8] sb_1__3_/chanx_right_in[9] cbx_2__3_/chanx_left_in[0]
+ cbx_2__3_/chanx_left_in[10] cbx_2__3_/chanx_left_in[11] cbx_2__3_/chanx_left_in[12]
+ cbx_2__3_/chanx_left_in[13] cbx_2__3_/chanx_left_in[14] cbx_2__3_/chanx_left_in[15]
+ cbx_2__3_/chanx_left_in[16] cbx_2__3_/chanx_left_in[17] cbx_2__3_/chanx_left_in[18]
+ cbx_2__3_/chanx_left_in[19] cbx_2__3_/chanx_left_in[1] cbx_2__3_/chanx_left_in[2]
+ cbx_2__3_/chanx_left_in[3] cbx_2__3_/chanx_left_in[4] cbx_2__3_/chanx_left_in[5]
+ cbx_2__3_/chanx_left_in[6] cbx_2__3_/chanx_left_in[7] cbx_2__3_/chanx_left_in[8]
+ cbx_2__3_/chanx_left_in[9] cby_1__3_/chany_top_out[0] cby_1__3_/chany_top_out[10]
+ cby_1__3_/chany_top_out[11] cby_1__3_/chany_top_out[12] cby_1__3_/chany_top_out[13]
+ cby_1__3_/chany_top_out[14] cby_1__3_/chany_top_out[15] cby_1__3_/chany_top_out[16]
+ cby_1__3_/chany_top_out[17] cby_1__3_/chany_top_out[18] cby_1__3_/chany_top_out[19]
+ cby_1__3_/chany_top_out[1] cby_1__3_/chany_top_out[2] cby_1__3_/chany_top_out[3]
+ cby_1__3_/chany_top_out[4] cby_1__3_/chany_top_out[5] cby_1__3_/chany_top_out[6]
+ cby_1__3_/chany_top_out[7] cby_1__3_/chany_top_out[8] cby_1__3_/chany_top_out[9]
+ cby_1__3_/chany_top_in[0] cby_1__3_/chany_top_in[10] cby_1__3_/chany_top_in[11]
+ cby_1__3_/chany_top_in[12] cby_1__3_/chany_top_in[13] cby_1__3_/chany_top_in[14]
+ cby_1__3_/chany_top_in[15] cby_1__3_/chany_top_in[16] cby_1__3_/chany_top_in[17]
+ cby_1__3_/chany_top_in[18] cby_1__3_/chany_top_in[19] cby_1__3_/chany_top_in[1]
+ cby_1__3_/chany_top_in[2] cby_1__3_/chany_top_in[3] cby_1__3_/chany_top_in[4] cby_1__3_/chany_top_in[5]
+ cby_1__3_/chany_top_in[6] cby_1__3_/chany_top_in[7] cby_1__3_/chany_top_in[8] cby_1__3_/chany_top_in[9]
+ sb_1__3_/chany_top_in[0] sb_1__3_/chany_top_in[10] sb_1__3_/chany_top_in[11] sb_1__3_/chany_top_in[12]
+ sb_1__3_/chany_top_in[13] sb_1__3_/chany_top_in[14] sb_1__3_/chany_top_in[15] sb_1__3_/chany_top_in[16]
+ sb_1__3_/chany_top_in[17] sb_1__3_/chany_top_in[18] sb_1__3_/chany_top_in[19] sb_1__3_/chany_top_in[1]
+ sb_1__3_/chany_top_in[2] sb_1__3_/chany_top_in[3] sb_1__3_/chany_top_in[4] sb_1__3_/chany_top_in[5]
+ sb_1__3_/chany_top_in[6] sb_1__3_/chany_top_in[7] sb_1__3_/chany_top_in[8] sb_1__3_/chany_top_in[9]
+ sb_1__3_/chany_top_out[0] sb_1__3_/chany_top_out[10] sb_1__3_/chany_top_out[11]
+ sb_1__3_/chany_top_out[12] sb_1__3_/chany_top_out[13] sb_1__3_/chany_top_out[14]
+ sb_1__3_/chany_top_out[15] sb_1__3_/chany_top_out[16] sb_1__3_/chany_top_out[17]
+ sb_1__3_/chany_top_out[18] sb_1__3_/chany_top_out[19] sb_1__3_/chany_top_out[1]
+ sb_1__3_/chany_top_out[2] sb_1__3_/chany_top_out[3] sb_1__3_/chany_top_out[4] sb_1__3_/chany_top_out[5]
+ sb_1__3_/chany_top_out[6] sb_1__3_/chany_top_out[7] sb_1__3_/chany_top_out[8] sb_1__3_/chany_top_out[9]
+ sb_1__3_/clk_1_E_out sb_1__3_/clk_1_N_in sb_1__3_/clk_1_W_out sb_1__3_/clk_2_E_out
+ sb_1__3_/clk_2_N_in sb_1__3_/clk_2_N_out sb_1__3_/clk_2_S_out sb_1__3_/clk_2_W_out
+ sb_1__3_/clk_3_E_out sb_1__3_/clk_3_N_in sb_1__3_/clk_3_N_out sb_1__3_/clk_3_S_out
+ sb_1__3_/clk_3_W_out sb_1__3_/left_bottom_grid_pin_34_ sb_1__3_/left_bottom_grid_pin_35_
+ sb_1__3_/left_bottom_grid_pin_36_ sb_1__3_/left_bottom_grid_pin_37_ sb_1__3_/left_bottom_grid_pin_38_
+ sb_1__3_/left_bottom_grid_pin_39_ sb_1__3_/left_bottom_grid_pin_40_ sb_1__3_/left_bottom_grid_pin_41_
+ sb_1__3_/prog_clk_0_N_in sb_1__3_/prog_clk_1_E_out sb_1__3_/prog_clk_1_N_in sb_1__3_/prog_clk_1_W_out
+ sb_1__3_/prog_clk_2_E_out sb_1__3_/prog_clk_2_N_in sb_1__3_/prog_clk_2_N_out sb_1__3_/prog_clk_2_S_out
+ sb_1__3_/prog_clk_2_W_out sb_1__3_/prog_clk_3_E_out sb_1__3_/prog_clk_3_N_in sb_1__3_/prog_clk_3_N_out
+ sb_1__3_/prog_clk_3_S_out sb_1__3_/prog_clk_3_W_out sb_1__3_/right_bottom_grid_pin_34_
+ sb_1__3_/right_bottom_grid_pin_35_ sb_1__3_/right_bottom_grid_pin_36_ sb_1__3_/right_bottom_grid_pin_37_
+ sb_1__3_/right_bottom_grid_pin_38_ sb_1__3_/right_bottom_grid_pin_39_ sb_1__3_/right_bottom_grid_pin_40_
+ sb_1__3_/right_bottom_grid_pin_41_ sb_1__3_/top_left_grid_pin_42_ sb_1__3_/top_left_grid_pin_43_
+ sb_1__3_/top_left_grid_pin_44_ sb_1__3_/top_left_grid_pin_45_ sb_1__3_/top_left_grid_pin_46_
+ sb_1__3_/top_left_grid_pin_47_ sb_1__3_/top_left_grid_pin_48_ sb_1__3_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_3__1_ cbx_3__1_/SC_OUT_BOT cbx_3__0_/SC_IN_TOP grid_clb_3__1_/SC_OUT_TOP
+ cby_3__1_/Test_en_W_out grid_clb_3__1_/Test_en_E_out cby_3__1_/Test_en_W_out cby_2__1_/Test_en_W_in
+ VGND VPWR grid_clb_3__1_/bottom_width_0_height_0__pin_50_ grid_clb_3__1_/bottom_width_0_height_0__pin_51_
+ cby_2__1_/ccff_tail cby_3__1_/ccff_head cbx_3__1_/clk_1_S_out cbx_3__1_/clk_1_S_out
+ cby_3__1_/prog_clk_0_W_in cbx_3__1_/prog_clk_1_S_out grid_clb_3__1_/prog_clk_0_N_out
+ cbx_3__1_/prog_clk_1_S_out cbx_3__0_/prog_clk_0_N_in grid_clb_3__1_/prog_clk_0_W_out
+ cby_3__1_/left_grid_pin_16_ cby_3__1_/left_grid_pin_17_ cby_3__1_/left_grid_pin_18_
+ cby_3__1_/left_grid_pin_19_ cby_3__1_/left_grid_pin_20_ cby_3__1_/left_grid_pin_21_
+ cby_3__1_/left_grid_pin_22_ cby_3__1_/left_grid_pin_23_ cby_3__1_/left_grid_pin_24_
+ cby_3__1_/left_grid_pin_25_ cby_3__1_/left_grid_pin_26_ cby_3__1_/left_grid_pin_27_
+ cby_3__1_/left_grid_pin_28_ cby_3__1_/left_grid_pin_29_ cby_3__1_/left_grid_pin_30_
+ cby_3__1_/left_grid_pin_31_ sb_3__0_/top_left_grid_pin_42_ sb_3__1_/bottom_left_grid_pin_42_
+ sb_3__0_/top_left_grid_pin_43_ sb_3__1_/bottom_left_grid_pin_43_ sb_3__0_/top_left_grid_pin_44_
+ sb_3__1_/bottom_left_grid_pin_44_ sb_3__0_/top_left_grid_pin_45_ sb_3__1_/bottom_left_grid_pin_45_
+ sb_3__0_/top_left_grid_pin_46_ sb_3__1_/bottom_left_grid_pin_46_ sb_3__0_/top_left_grid_pin_47_
+ sb_3__1_/bottom_left_grid_pin_47_ sb_3__0_/top_left_grid_pin_48_ sb_3__1_/bottom_left_grid_pin_48_
+ sb_3__0_/top_left_grid_pin_49_ sb_3__1_/bottom_left_grid_pin_49_ cbx_3__1_/bottom_grid_pin_0_
+ cbx_3__1_/bottom_grid_pin_10_ cbx_3__1_/bottom_grid_pin_11_ cbx_3__1_/bottom_grid_pin_12_
+ cbx_3__1_/bottom_grid_pin_13_ cbx_3__1_/bottom_grid_pin_14_ cbx_3__1_/bottom_grid_pin_15_
+ cbx_3__1_/bottom_grid_pin_1_ cbx_3__1_/bottom_grid_pin_2_ cbx_3__1_/REGOUT_FEEDTHROUGH
+ grid_clb_3__1_/top_width_0_height_0__pin_33_ sb_3__1_/left_bottom_grid_pin_34_ sb_2__1_/right_bottom_grid_pin_34_
+ sb_3__1_/left_bottom_grid_pin_35_ sb_2__1_/right_bottom_grid_pin_35_ sb_3__1_/left_bottom_grid_pin_36_
+ sb_2__1_/right_bottom_grid_pin_36_ sb_3__1_/left_bottom_grid_pin_37_ sb_2__1_/right_bottom_grid_pin_37_
+ sb_3__1_/left_bottom_grid_pin_38_ sb_2__1_/right_bottom_grid_pin_38_ sb_3__1_/left_bottom_grid_pin_39_
+ sb_2__1_/right_bottom_grid_pin_39_ cbx_3__1_/bottom_grid_pin_3_ sb_3__1_/left_bottom_grid_pin_40_
+ sb_2__1_/right_bottom_grid_pin_40_ sb_3__1_/left_bottom_grid_pin_41_ sb_2__1_/right_bottom_grid_pin_41_
+ cbx_3__1_/bottom_grid_pin_4_ cbx_3__1_/bottom_grid_pin_5_ cbx_3__1_/bottom_grid_pin_6_
+ cbx_3__1_/bottom_grid_pin_7_ cbx_3__1_/bottom_grid_pin_8_ cbx_3__1_/bottom_grid_pin_9_
+ grid_clb
Xcby_7__2_ cby_7__2_/Test_en_W_in cby_7__2_/Test_en_E_out cby_7__2_/Test_en_N_out
+ cby_7__2_/Test_en_W_in cby_7__2_/Test_en_W_in cby_7__2_/Test_en_W_out VGND VPWR
+ cby_7__2_/ccff_head cby_7__2_/ccff_tail sb_7__1_/chany_top_out[0] sb_7__1_/chany_top_out[10]
+ sb_7__1_/chany_top_out[11] sb_7__1_/chany_top_out[12] sb_7__1_/chany_top_out[13]
+ sb_7__1_/chany_top_out[14] sb_7__1_/chany_top_out[15] sb_7__1_/chany_top_out[16]
+ sb_7__1_/chany_top_out[17] sb_7__1_/chany_top_out[18] sb_7__1_/chany_top_out[19]
+ sb_7__1_/chany_top_out[1] sb_7__1_/chany_top_out[2] sb_7__1_/chany_top_out[3] sb_7__1_/chany_top_out[4]
+ sb_7__1_/chany_top_out[5] sb_7__1_/chany_top_out[6] sb_7__1_/chany_top_out[7] sb_7__1_/chany_top_out[8]
+ sb_7__1_/chany_top_out[9] sb_7__1_/chany_top_in[0] sb_7__1_/chany_top_in[10] sb_7__1_/chany_top_in[11]
+ sb_7__1_/chany_top_in[12] sb_7__1_/chany_top_in[13] sb_7__1_/chany_top_in[14] sb_7__1_/chany_top_in[15]
+ sb_7__1_/chany_top_in[16] sb_7__1_/chany_top_in[17] sb_7__1_/chany_top_in[18] sb_7__1_/chany_top_in[19]
+ sb_7__1_/chany_top_in[1] sb_7__1_/chany_top_in[2] sb_7__1_/chany_top_in[3] sb_7__1_/chany_top_in[4]
+ sb_7__1_/chany_top_in[5] sb_7__1_/chany_top_in[6] sb_7__1_/chany_top_in[7] sb_7__1_/chany_top_in[8]
+ sb_7__1_/chany_top_in[9] cby_7__2_/chany_top_in[0] cby_7__2_/chany_top_in[10] cby_7__2_/chany_top_in[11]
+ cby_7__2_/chany_top_in[12] cby_7__2_/chany_top_in[13] cby_7__2_/chany_top_in[14]
+ cby_7__2_/chany_top_in[15] cby_7__2_/chany_top_in[16] cby_7__2_/chany_top_in[17]
+ cby_7__2_/chany_top_in[18] cby_7__2_/chany_top_in[19] cby_7__2_/chany_top_in[1]
+ cby_7__2_/chany_top_in[2] cby_7__2_/chany_top_in[3] cby_7__2_/chany_top_in[4] cby_7__2_/chany_top_in[5]
+ cby_7__2_/chany_top_in[6] cby_7__2_/chany_top_in[7] cby_7__2_/chany_top_in[8] cby_7__2_/chany_top_in[9]
+ cby_7__2_/chany_top_out[0] cby_7__2_/chany_top_out[10] cby_7__2_/chany_top_out[11]
+ cby_7__2_/chany_top_out[12] cby_7__2_/chany_top_out[13] cby_7__2_/chany_top_out[14]
+ cby_7__2_/chany_top_out[15] cby_7__2_/chany_top_out[16] cby_7__2_/chany_top_out[17]
+ cby_7__2_/chany_top_out[18] cby_7__2_/chany_top_out[19] cby_7__2_/chany_top_out[1]
+ cby_7__2_/chany_top_out[2] cby_7__2_/chany_top_out[3] cby_7__2_/chany_top_out[4]
+ cby_7__2_/chany_top_out[5] cby_7__2_/chany_top_out[6] cby_7__2_/chany_top_out[7]
+ cby_7__2_/chany_top_out[8] cby_7__2_/chany_top_out[9] cby_7__2_/clk_2_N_out sb_7__2_/clk_2_S_out
+ sb_7__1_/clk_1_N_in cby_7__2_/clk_3_N_out cby_7__2_/clk_3_S_in cby_7__2_/clk_3_S_out
+ cby_7__2_/left_grid_pin_16_ cby_7__2_/left_grid_pin_17_ cby_7__2_/left_grid_pin_18_
+ cby_7__2_/left_grid_pin_19_ cby_7__2_/left_grid_pin_20_ cby_7__2_/left_grid_pin_21_
+ cby_7__2_/left_grid_pin_22_ cby_7__2_/left_grid_pin_23_ cby_7__2_/left_grid_pin_24_
+ cby_7__2_/left_grid_pin_25_ cby_7__2_/left_grid_pin_26_ cby_7__2_/left_grid_pin_27_
+ cby_7__2_/left_grid_pin_28_ cby_7__2_/left_grid_pin_29_ cby_7__2_/left_grid_pin_30_
+ cby_7__2_/left_grid_pin_31_ cby_7__2_/prog_clk_0_N_out sb_7__1_/prog_clk_0_N_in
+ cby_7__2_/prog_clk_0_W_in cby_7__2_/prog_clk_2_N_out sb_7__2_/prog_clk_2_S_out sb_7__1_/prog_clk_1_N_in
+ cby_7__2_/prog_clk_3_N_out cby_7__2_/prog_clk_3_S_in cby_7__2_/prog_clk_3_S_out
+ cby_1__1_
Xcby_0__7_ IO_ISOL_N VGND VPWR sb_0__7_/ccff_tail cby_0__7_/ccff_tail sb_0__6_/chany_top_out[0]
+ sb_0__6_/chany_top_out[10] sb_0__6_/chany_top_out[11] sb_0__6_/chany_top_out[12]
+ sb_0__6_/chany_top_out[13] sb_0__6_/chany_top_out[14] sb_0__6_/chany_top_out[15]
+ sb_0__6_/chany_top_out[16] sb_0__6_/chany_top_out[17] sb_0__6_/chany_top_out[18]
+ sb_0__6_/chany_top_out[19] sb_0__6_/chany_top_out[1] sb_0__6_/chany_top_out[2] sb_0__6_/chany_top_out[3]
+ sb_0__6_/chany_top_out[4] sb_0__6_/chany_top_out[5] sb_0__6_/chany_top_out[6] sb_0__6_/chany_top_out[7]
+ sb_0__6_/chany_top_out[8] sb_0__6_/chany_top_out[9] sb_0__6_/chany_top_in[0] sb_0__6_/chany_top_in[10]
+ sb_0__6_/chany_top_in[11] sb_0__6_/chany_top_in[12] sb_0__6_/chany_top_in[13] sb_0__6_/chany_top_in[14]
+ sb_0__6_/chany_top_in[15] sb_0__6_/chany_top_in[16] sb_0__6_/chany_top_in[17] sb_0__6_/chany_top_in[18]
+ sb_0__6_/chany_top_in[19] sb_0__6_/chany_top_in[1] sb_0__6_/chany_top_in[2] sb_0__6_/chany_top_in[3]
+ sb_0__6_/chany_top_in[4] sb_0__6_/chany_top_in[5] sb_0__6_/chany_top_in[6] sb_0__6_/chany_top_in[7]
+ sb_0__6_/chany_top_in[8] sb_0__6_/chany_top_in[9] cby_0__7_/chany_top_in[0] cby_0__7_/chany_top_in[10]
+ cby_0__7_/chany_top_in[11] cby_0__7_/chany_top_in[12] cby_0__7_/chany_top_in[13]
+ cby_0__7_/chany_top_in[14] cby_0__7_/chany_top_in[15] cby_0__7_/chany_top_in[16]
+ cby_0__7_/chany_top_in[17] cby_0__7_/chany_top_in[18] cby_0__7_/chany_top_in[19]
+ cby_0__7_/chany_top_in[1] cby_0__7_/chany_top_in[2] cby_0__7_/chany_top_in[3] cby_0__7_/chany_top_in[4]
+ cby_0__7_/chany_top_in[5] cby_0__7_/chany_top_in[6] cby_0__7_/chany_top_in[7] cby_0__7_/chany_top_in[8]
+ cby_0__7_/chany_top_in[9] cby_0__7_/chany_top_out[0] cby_0__7_/chany_top_out[10]
+ cby_0__7_/chany_top_out[11] cby_0__7_/chany_top_out[12] cby_0__7_/chany_top_out[13]
+ cby_0__7_/chany_top_out[14] cby_0__7_/chany_top_out[15] cby_0__7_/chany_top_out[16]
+ cby_0__7_/chany_top_out[17] cby_0__7_/chany_top_out[18] cby_0__7_/chany_top_out[19]
+ cby_0__7_/chany_top_out[1] cby_0__7_/chany_top_out[2] cby_0__7_/chany_top_out[3]
+ cby_0__7_/chany_top_out[4] cby_0__7_/chany_top_out[5] cby_0__7_/chany_top_out[6]
+ cby_0__7_/chany_top_out[7] cby_0__7_/chany_top_out[8] cby_0__7_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
+ cby_0__7_/left_grid_pin_0_ cby_0__7_/prog_clk_0_E_in cby_0__7_/left_grid_pin_0_
+ sb_0__6_/top_left_grid_pin_1_ sb_0__7_/bottom_left_grid_pin_1_ cby_0__1_
Xcbx_7__3_ cbx_7__3_/REGIN_FEEDTHROUGH cbx_7__3_/REGOUT_FEEDTHROUGH cbx_7__3_/SC_IN_BOT
+ cbx_7__3_/SC_IN_TOP cbx_7__3_/SC_OUT_BOT cbx_7__3_/SC_OUT_TOP VGND VPWR cbx_7__3_/bottom_grid_pin_0_
+ cbx_7__3_/bottom_grid_pin_10_ cbx_7__3_/bottom_grid_pin_11_ cbx_7__3_/bottom_grid_pin_12_
+ cbx_7__3_/bottom_grid_pin_13_ cbx_7__3_/bottom_grid_pin_14_ cbx_7__3_/bottom_grid_pin_15_
+ cbx_7__3_/bottom_grid_pin_1_ cbx_7__3_/bottom_grid_pin_2_ cbx_7__3_/bottom_grid_pin_3_
+ cbx_7__3_/bottom_grid_pin_4_ cbx_7__3_/bottom_grid_pin_5_ cbx_7__3_/bottom_grid_pin_6_
+ cbx_7__3_/bottom_grid_pin_7_ cbx_7__3_/bottom_grid_pin_8_ cbx_7__3_/bottom_grid_pin_9_
+ sb_7__3_/ccff_tail sb_6__3_/ccff_head cbx_7__3_/chanx_left_in[0] cbx_7__3_/chanx_left_in[10]
+ cbx_7__3_/chanx_left_in[11] cbx_7__3_/chanx_left_in[12] cbx_7__3_/chanx_left_in[13]
+ cbx_7__3_/chanx_left_in[14] cbx_7__3_/chanx_left_in[15] cbx_7__3_/chanx_left_in[16]
+ cbx_7__3_/chanx_left_in[17] cbx_7__3_/chanx_left_in[18] cbx_7__3_/chanx_left_in[19]
+ cbx_7__3_/chanx_left_in[1] cbx_7__3_/chanx_left_in[2] cbx_7__3_/chanx_left_in[3]
+ cbx_7__3_/chanx_left_in[4] cbx_7__3_/chanx_left_in[5] cbx_7__3_/chanx_left_in[6]
+ cbx_7__3_/chanx_left_in[7] cbx_7__3_/chanx_left_in[8] cbx_7__3_/chanx_left_in[9]
+ sb_6__3_/chanx_right_in[0] sb_6__3_/chanx_right_in[10] sb_6__3_/chanx_right_in[11]
+ sb_6__3_/chanx_right_in[12] sb_6__3_/chanx_right_in[13] sb_6__3_/chanx_right_in[14]
+ sb_6__3_/chanx_right_in[15] sb_6__3_/chanx_right_in[16] sb_6__3_/chanx_right_in[17]
+ sb_6__3_/chanx_right_in[18] sb_6__3_/chanx_right_in[19] sb_6__3_/chanx_right_in[1]
+ sb_6__3_/chanx_right_in[2] sb_6__3_/chanx_right_in[3] sb_6__3_/chanx_right_in[4]
+ sb_6__3_/chanx_right_in[5] sb_6__3_/chanx_right_in[6] sb_6__3_/chanx_right_in[7]
+ sb_6__3_/chanx_right_in[8] sb_6__3_/chanx_right_in[9] sb_7__3_/chanx_left_out[0]
+ sb_7__3_/chanx_left_out[10] sb_7__3_/chanx_left_out[11] sb_7__3_/chanx_left_out[12]
+ sb_7__3_/chanx_left_out[13] sb_7__3_/chanx_left_out[14] sb_7__3_/chanx_left_out[15]
+ sb_7__3_/chanx_left_out[16] sb_7__3_/chanx_left_out[17] sb_7__3_/chanx_left_out[18]
+ sb_7__3_/chanx_left_out[19] sb_7__3_/chanx_left_out[1] sb_7__3_/chanx_left_out[2]
+ sb_7__3_/chanx_left_out[3] sb_7__3_/chanx_left_out[4] sb_7__3_/chanx_left_out[5]
+ sb_7__3_/chanx_left_out[6] sb_7__3_/chanx_left_out[7] sb_7__3_/chanx_left_out[8]
+ sb_7__3_/chanx_left_out[9] sb_7__3_/chanx_left_in[0] sb_7__3_/chanx_left_in[10]
+ sb_7__3_/chanx_left_in[11] sb_7__3_/chanx_left_in[12] sb_7__3_/chanx_left_in[13]
+ sb_7__3_/chanx_left_in[14] sb_7__3_/chanx_left_in[15] sb_7__3_/chanx_left_in[16]
+ sb_7__3_/chanx_left_in[17] sb_7__3_/chanx_left_in[18] sb_7__3_/chanx_left_in[19]
+ sb_7__3_/chanx_left_in[1] sb_7__3_/chanx_left_in[2] sb_7__3_/chanx_left_in[3] sb_7__3_/chanx_left_in[4]
+ sb_7__3_/chanx_left_in[5] sb_7__3_/chanx_left_in[6] sb_7__3_/chanx_left_in[7] sb_7__3_/chanx_left_in[8]
+ sb_7__3_/chanx_left_in[9] cbx_7__3_/clk_1_N_out cbx_7__3_/clk_1_S_out sb_7__3_/clk_1_W_out
+ cbx_7__3_/clk_2_E_out cbx_7__3_/clk_2_W_in cbx_7__3_/clk_2_W_out cbx_7__3_/clk_3_E_out
+ cbx_7__3_/clk_3_W_in cbx_7__3_/clk_3_W_out cbx_7__3_/prog_clk_0_N_in cbx_7__3_/prog_clk_0_W_out
+ cbx_7__3_/prog_clk_1_N_out cbx_7__3_/prog_clk_1_S_out sb_7__3_/prog_clk_1_W_out
+ cbx_7__3_/prog_clk_2_E_out cbx_7__3_/prog_clk_2_W_in cbx_7__3_/prog_clk_2_W_out
+ cbx_7__3_/prog_clk_3_E_out cbx_7__3_/prog_clk_3_W_in cbx_7__3_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_7__8_ sb_7__8_/SC_IN_BOT sb_7__8_/SC_OUT_BOT VGND VPWR sb_7__8_/bottom_left_grid_pin_42_
+ sb_7__8_/bottom_left_grid_pin_43_ sb_7__8_/bottom_left_grid_pin_44_ sb_7__8_/bottom_left_grid_pin_45_
+ sb_7__8_/bottom_left_grid_pin_46_ sb_7__8_/bottom_left_grid_pin_47_ sb_7__8_/bottom_left_grid_pin_48_
+ sb_7__8_/bottom_left_grid_pin_49_ sb_7__8_/ccff_head sb_7__8_/ccff_tail sb_7__8_/chanx_left_in[0]
+ sb_7__8_/chanx_left_in[10] sb_7__8_/chanx_left_in[11] sb_7__8_/chanx_left_in[12]
+ sb_7__8_/chanx_left_in[13] sb_7__8_/chanx_left_in[14] sb_7__8_/chanx_left_in[15]
+ sb_7__8_/chanx_left_in[16] sb_7__8_/chanx_left_in[17] sb_7__8_/chanx_left_in[18]
+ sb_7__8_/chanx_left_in[19] sb_7__8_/chanx_left_in[1] sb_7__8_/chanx_left_in[2] sb_7__8_/chanx_left_in[3]
+ sb_7__8_/chanx_left_in[4] sb_7__8_/chanx_left_in[5] sb_7__8_/chanx_left_in[6] sb_7__8_/chanx_left_in[7]
+ sb_7__8_/chanx_left_in[8] sb_7__8_/chanx_left_in[9] sb_7__8_/chanx_left_out[0] sb_7__8_/chanx_left_out[10]
+ sb_7__8_/chanx_left_out[11] sb_7__8_/chanx_left_out[12] sb_7__8_/chanx_left_out[13]
+ sb_7__8_/chanx_left_out[14] sb_7__8_/chanx_left_out[15] sb_7__8_/chanx_left_out[16]
+ sb_7__8_/chanx_left_out[17] sb_7__8_/chanx_left_out[18] sb_7__8_/chanx_left_out[19]
+ sb_7__8_/chanx_left_out[1] sb_7__8_/chanx_left_out[2] sb_7__8_/chanx_left_out[3]
+ sb_7__8_/chanx_left_out[4] sb_7__8_/chanx_left_out[5] sb_7__8_/chanx_left_out[6]
+ sb_7__8_/chanx_left_out[7] sb_7__8_/chanx_left_out[8] sb_7__8_/chanx_left_out[9]
+ sb_7__8_/chanx_right_in[0] sb_7__8_/chanx_right_in[10] sb_7__8_/chanx_right_in[11]
+ sb_7__8_/chanx_right_in[12] sb_7__8_/chanx_right_in[13] sb_7__8_/chanx_right_in[14]
+ sb_7__8_/chanx_right_in[15] sb_7__8_/chanx_right_in[16] sb_7__8_/chanx_right_in[17]
+ sb_7__8_/chanx_right_in[18] sb_7__8_/chanx_right_in[19] sb_7__8_/chanx_right_in[1]
+ sb_7__8_/chanx_right_in[2] sb_7__8_/chanx_right_in[3] sb_7__8_/chanx_right_in[4]
+ sb_7__8_/chanx_right_in[5] sb_7__8_/chanx_right_in[6] sb_7__8_/chanx_right_in[7]
+ sb_7__8_/chanx_right_in[8] sb_7__8_/chanx_right_in[9] cbx_8__8_/chanx_left_in[0]
+ cbx_8__8_/chanx_left_in[10] cbx_8__8_/chanx_left_in[11] cbx_8__8_/chanx_left_in[12]
+ cbx_8__8_/chanx_left_in[13] cbx_8__8_/chanx_left_in[14] cbx_8__8_/chanx_left_in[15]
+ cbx_8__8_/chanx_left_in[16] cbx_8__8_/chanx_left_in[17] cbx_8__8_/chanx_left_in[18]
+ cbx_8__8_/chanx_left_in[19] cbx_8__8_/chanx_left_in[1] cbx_8__8_/chanx_left_in[2]
+ cbx_8__8_/chanx_left_in[3] cbx_8__8_/chanx_left_in[4] cbx_8__8_/chanx_left_in[5]
+ cbx_8__8_/chanx_left_in[6] cbx_8__8_/chanx_left_in[7] cbx_8__8_/chanx_left_in[8]
+ cbx_8__8_/chanx_left_in[9] cby_7__8_/chany_top_out[0] cby_7__8_/chany_top_out[10]
+ cby_7__8_/chany_top_out[11] cby_7__8_/chany_top_out[12] cby_7__8_/chany_top_out[13]
+ cby_7__8_/chany_top_out[14] cby_7__8_/chany_top_out[15] cby_7__8_/chany_top_out[16]
+ cby_7__8_/chany_top_out[17] cby_7__8_/chany_top_out[18] cby_7__8_/chany_top_out[19]
+ cby_7__8_/chany_top_out[1] cby_7__8_/chany_top_out[2] cby_7__8_/chany_top_out[3]
+ cby_7__8_/chany_top_out[4] cby_7__8_/chany_top_out[5] cby_7__8_/chany_top_out[6]
+ cby_7__8_/chany_top_out[7] cby_7__8_/chany_top_out[8] cby_7__8_/chany_top_out[9]
+ cby_7__8_/chany_top_in[0] cby_7__8_/chany_top_in[10] cby_7__8_/chany_top_in[11]
+ cby_7__8_/chany_top_in[12] cby_7__8_/chany_top_in[13] cby_7__8_/chany_top_in[14]
+ cby_7__8_/chany_top_in[15] cby_7__8_/chany_top_in[16] cby_7__8_/chany_top_in[17]
+ cby_7__8_/chany_top_in[18] cby_7__8_/chany_top_in[19] cby_7__8_/chany_top_in[1]
+ cby_7__8_/chany_top_in[2] cby_7__8_/chany_top_in[3] cby_7__8_/chany_top_in[4] cby_7__8_/chany_top_in[5]
+ cby_7__8_/chany_top_in[6] cby_7__8_/chany_top_in[7] cby_7__8_/chany_top_in[8] cby_7__8_/chany_top_in[9]
+ sb_7__8_/left_bottom_grid_pin_34_ sb_7__8_/left_bottom_grid_pin_35_ sb_7__8_/left_bottom_grid_pin_36_
+ sb_7__8_/left_bottom_grid_pin_37_ sb_7__8_/left_bottom_grid_pin_38_ sb_7__8_/left_bottom_grid_pin_39_
+ sb_7__8_/left_bottom_grid_pin_40_ sb_7__8_/left_bottom_grid_pin_41_ sb_7__8_/left_top_grid_pin_1_
+ sb_7__8_/prog_clk_0_S_in sb_7__8_/right_bottom_grid_pin_34_ sb_7__8_/right_bottom_grid_pin_35_
+ sb_7__8_/right_bottom_grid_pin_36_ sb_7__8_/right_bottom_grid_pin_37_ sb_7__8_/right_bottom_grid_pin_38_
+ sb_7__8_/right_bottom_grid_pin_39_ sb_7__8_/right_bottom_grid_pin_40_ sb_7__8_/right_bottom_grid_pin_41_
+ sb_7__8_/right_top_grid_pin_1_ sb_1__2_
Xsb_4__5_ sb_4__5_/Test_en_N_out sb_4__5_/Test_en_S_in VGND VPWR sb_4__5_/bottom_left_grid_pin_42_
+ sb_4__5_/bottom_left_grid_pin_43_ sb_4__5_/bottom_left_grid_pin_44_ sb_4__5_/bottom_left_grid_pin_45_
+ sb_4__5_/bottom_left_grid_pin_46_ sb_4__5_/bottom_left_grid_pin_47_ sb_4__5_/bottom_left_grid_pin_48_
+ sb_4__5_/bottom_left_grid_pin_49_ sb_4__5_/ccff_head sb_4__5_/ccff_tail sb_4__5_/chanx_left_in[0]
+ sb_4__5_/chanx_left_in[10] sb_4__5_/chanx_left_in[11] sb_4__5_/chanx_left_in[12]
+ sb_4__5_/chanx_left_in[13] sb_4__5_/chanx_left_in[14] sb_4__5_/chanx_left_in[15]
+ sb_4__5_/chanx_left_in[16] sb_4__5_/chanx_left_in[17] sb_4__5_/chanx_left_in[18]
+ sb_4__5_/chanx_left_in[19] sb_4__5_/chanx_left_in[1] sb_4__5_/chanx_left_in[2] sb_4__5_/chanx_left_in[3]
+ sb_4__5_/chanx_left_in[4] sb_4__5_/chanx_left_in[5] sb_4__5_/chanx_left_in[6] sb_4__5_/chanx_left_in[7]
+ sb_4__5_/chanx_left_in[8] sb_4__5_/chanx_left_in[9] sb_4__5_/chanx_left_out[0] sb_4__5_/chanx_left_out[10]
+ sb_4__5_/chanx_left_out[11] sb_4__5_/chanx_left_out[12] sb_4__5_/chanx_left_out[13]
+ sb_4__5_/chanx_left_out[14] sb_4__5_/chanx_left_out[15] sb_4__5_/chanx_left_out[16]
+ sb_4__5_/chanx_left_out[17] sb_4__5_/chanx_left_out[18] sb_4__5_/chanx_left_out[19]
+ sb_4__5_/chanx_left_out[1] sb_4__5_/chanx_left_out[2] sb_4__5_/chanx_left_out[3]
+ sb_4__5_/chanx_left_out[4] sb_4__5_/chanx_left_out[5] sb_4__5_/chanx_left_out[6]
+ sb_4__5_/chanx_left_out[7] sb_4__5_/chanx_left_out[8] sb_4__5_/chanx_left_out[9]
+ sb_4__5_/chanx_right_in[0] sb_4__5_/chanx_right_in[10] sb_4__5_/chanx_right_in[11]
+ sb_4__5_/chanx_right_in[12] sb_4__5_/chanx_right_in[13] sb_4__5_/chanx_right_in[14]
+ sb_4__5_/chanx_right_in[15] sb_4__5_/chanx_right_in[16] sb_4__5_/chanx_right_in[17]
+ sb_4__5_/chanx_right_in[18] sb_4__5_/chanx_right_in[19] sb_4__5_/chanx_right_in[1]
+ sb_4__5_/chanx_right_in[2] sb_4__5_/chanx_right_in[3] sb_4__5_/chanx_right_in[4]
+ sb_4__5_/chanx_right_in[5] sb_4__5_/chanx_right_in[6] sb_4__5_/chanx_right_in[7]
+ sb_4__5_/chanx_right_in[8] sb_4__5_/chanx_right_in[9] cbx_5__5_/chanx_left_in[0]
+ cbx_5__5_/chanx_left_in[10] cbx_5__5_/chanx_left_in[11] cbx_5__5_/chanx_left_in[12]
+ cbx_5__5_/chanx_left_in[13] cbx_5__5_/chanx_left_in[14] cbx_5__5_/chanx_left_in[15]
+ cbx_5__5_/chanx_left_in[16] cbx_5__5_/chanx_left_in[17] cbx_5__5_/chanx_left_in[18]
+ cbx_5__5_/chanx_left_in[19] cbx_5__5_/chanx_left_in[1] cbx_5__5_/chanx_left_in[2]
+ cbx_5__5_/chanx_left_in[3] cbx_5__5_/chanx_left_in[4] cbx_5__5_/chanx_left_in[5]
+ cbx_5__5_/chanx_left_in[6] cbx_5__5_/chanx_left_in[7] cbx_5__5_/chanx_left_in[8]
+ cbx_5__5_/chanx_left_in[9] cby_4__5_/chany_top_out[0] cby_4__5_/chany_top_out[10]
+ cby_4__5_/chany_top_out[11] cby_4__5_/chany_top_out[12] cby_4__5_/chany_top_out[13]
+ cby_4__5_/chany_top_out[14] cby_4__5_/chany_top_out[15] cby_4__5_/chany_top_out[16]
+ cby_4__5_/chany_top_out[17] cby_4__5_/chany_top_out[18] cby_4__5_/chany_top_out[19]
+ cby_4__5_/chany_top_out[1] cby_4__5_/chany_top_out[2] cby_4__5_/chany_top_out[3]
+ cby_4__5_/chany_top_out[4] cby_4__5_/chany_top_out[5] cby_4__5_/chany_top_out[6]
+ cby_4__5_/chany_top_out[7] cby_4__5_/chany_top_out[8] cby_4__5_/chany_top_out[9]
+ cby_4__5_/chany_top_in[0] cby_4__5_/chany_top_in[10] cby_4__5_/chany_top_in[11]
+ cby_4__5_/chany_top_in[12] cby_4__5_/chany_top_in[13] cby_4__5_/chany_top_in[14]
+ cby_4__5_/chany_top_in[15] cby_4__5_/chany_top_in[16] cby_4__5_/chany_top_in[17]
+ cby_4__5_/chany_top_in[18] cby_4__5_/chany_top_in[19] cby_4__5_/chany_top_in[1]
+ cby_4__5_/chany_top_in[2] cby_4__5_/chany_top_in[3] cby_4__5_/chany_top_in[4] cby_4__5_/chany_top_in[5]
+ cby_4__5_/chany_top_in[6] cby_4__5_/chany_top_in[7] cby_4__5_/chany_top_in[8] cby_4__5_/chany_top_in[9]
+ sb_4__5_/chany_top_in[0] sb_4__5_/chany_top_in[10] sb_4__5_/chany_top_in[11] sb_4__5_/chany_top_in[12]
+ sb_4__5_/chany_top_in[13] sb_4__5_/chany_top_in[14] sb_4__5_/chany_top_in[15] sb_4__5_/chany_top_in[16]
+ sb_4__5_/chany_top_in[17] sb_4__5_/chany_top_in[18] sb_4__5_/chany_top_in[19] sb_4__5_/chany_top_in[1]
+ sb_4__5_/chany_top_in[2] sb_4__5_/chany_top_in[3] sb_4__5_/chany_top_in[4] sb_4__5_/chany_top_in[5]
+ sb_4__5_/chany_top_in[6] sb_4__5_/chany_top_in[7] sb_4__5_/chany_top_in[8] sb_4__5_/chany_top_in[9]
+ sb_4__5_/chany_top_out[0] sb_4__5_/chany_top_out[10] sb_4__5_/chany_top_out[11]
+ sb_4__5_/chany_top_out[12] sb_4__5_/chany_top_out[13] sb_4__5_/chany_top_out[14]
+ sb_4__5_/chany_top_out[15] sb_4__5_/chany_top_out[16] sb_4__5_/chany_top_out[17]
+ sb_4__5_/chany_top_out[18] sb_4__5_/chany_top_out[19] sb_4__5_/chany_top_out[1]
+ sb_4__5_/chany_top_out[2] sb_4__5_/chany_top_out[3] sb_4__5_/chany_top_out[4] sb_4__5_/chany_top_out[5]
+ sb_4__5_/chany_top_out[6] sb_4__5_/chany_top_out[7] sb_4__5_/chany_top_out[8] sb_4__5_/chany_top_out[9]
+ sb_4__5_/clk_1_E_out sb_4__5_/clk_1_N_in sb_4__5_/clk_1_W_out sb_4__5_/clk_2_E_out
+ sb_4__5_/clk_2_N_in sb_4__5_/clk_2_N_out sb_4__5_/clk_2_S_out sb_4__5_/clk_2_W_out
+ sb_4__5_/clk_3_E_out sb_4__5_/clk_3_N_in sb_4__5_/clk_3_N_out sb_4__5_/clk_3_S_out
+ sb_4__5_/clk_3_W_out sb_4__5_/left_bottom_grid_pin_34_ sb_4__5_/left_bottom_grid_pin_35_
+ sb_4__5_/left_bottom_grid_pin_36_ sb_4__5_/left_bottom_grid_pin_37_ sb_4__5_/left_bottom_grid_pin_38_
+ sb_4__5_/left_bottom_grid_pin_39_ sb_4__5_/left_bottom_grid_pin_40_ sb_4__5_/left_bottom_grid_pin_41_
+ sb_4__5_/prog_clk_0_N_in sb_4__5_/prog_clk_1_E_out sb_4__5_/prog_clk_1_N_in sb_4__5_/prog_clk_1_W_out
+ sb_4__5_/prog_clk_2_E_out sb_4__5_/prog_clk_2_N_in sb_4__5_/prog_clk_2_N_out sb_4__5_/prog_clk_2_S_out
+ sb_4__5_/prog_clk_2_W_out sb_4__5_/prog_clk_3_E_out sb_4__5_/prog_clk_3_N_in sb_4__5_/prog_clk_3_N_out
+ sb_4__5_/prog_clk_3_S_out sb_4__5_/prog_clk_3_W_out sb_4__5_/right_bottom_grid_pin_34_
+ sb_4__5_/right_bottom_grid_pin_35_ sb_4__5_/right_bottom_grid_pin_36_ sb_4__5_/right_bottom_grid_pin_37_
+ sb_4__5_/right_bottom_grid_pin_38_ sb_4__5_/right_bottom_grid_pin_39_ sb_4__5_/right_bottom_grid_pin_40_
+ sb_4__5_/right_bottom_grid_pin_41_ sb_4__5_/top_left_grid_pin_42_ sb_4__5_/top_left_grid_pin_43_
+ sb_4__5_/top_left_grid_pin_44_ sb_4__5_/top_left_grid_pin_45_ sb_4__5_/top_left_grid_pin_46_
+ sb_4__5_/top_left_grid_pin_47_ sb_4__5_/top_left_grid_pin_48_ sb_4__5_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_6__3_ cbx_6__2_/SC_OUT_TOP grid_clb_6__3_/SC_OUT_BOT cbx_6__3_/SC_IN_BOT
+ cby_5__3_/Test_en_E_out cby_6__3_/Test_en_W_in cby_5__3_/Test_en_E_out grid_clb_6__3_/Test_en_W_out
+ VGND VPWR cbx_6__2_/REGIN_FEEDTHROUGH grid_clb_6__3_/bottom_width_0_height_0__pin_51_
+ cby_5__3_/ccff_tail cby_6__3_/ccff_head cbx_6__3_/clk_1_S_out cbx_6__3_/clk_1_S_out
+ cby_6__3_/prog_clk_0_W_in cbx_6__3_/prog_clk_1_S_out grid_clb_6__3_/prog_clk_0_N_out
+ cbx_6__3_/prog_clk_1_S_out cbx_6__2_/prog_clk_0_N_in grid_clb_6__3_/prog_clk_0_W_out
+ cby_6__3_/left_grid_pin_16_ cby_6__3_/left_grid_pin_17_ cby_6__3_/left_grid_pin_18_
+ cby_6__3_/left_grid_pin_19_ cby_6__3_/left_grid_pin_20_ cby_6__3_/left_grid_pin_21_
+ cby_6__3_/left_grid_pin_22_ cby_6__3_/left_grid_pin_23_ cby_6__3_/left_grid_pin_24_
+ cby_6__3_/left_grid_pin_25_ cby_6__3_/left_grid_pin_26_ cby_6__3_/left_grid_pin_27_
+ cby_6__3_/left_grid_pin_28_ cby_6__3_/left_grid_pin_29_ cby_6__3_/left_grid_pin_30_
+ cby_6__3_/left_grid_pin_31_ sb_6__2_/top_left_grid_pin_42_ sb_6__3_/bottom_left_grid_pin_42_
+ sb_6__2_/top_left_grid_pin_43_ sb_6__3_/bottom_left_grid_pin_43_ sb_6__2_/top_left_grid_pin_44_
+ sb_6__3_/bottom_left_grid_pin_44_ sb_6__2_/top_left_grid_pin_45_ sb_6__3_/bottom_left_grid_pin_45_
+ sb_6__2_/top_left_grid_pin_46_ sb_6__3_/bottom_left_grid_pin_46_ sb_6__2_/top_left_grid_pin_47_
+ sb_6__3_/bottom_left_grid_pin_47_ sb_6__2_/top_left_grid_pin_48_ sb_6__3_/bottom_left_grid_pin_48_
+ sb_6__2_/top_left_grid_pin_49_ sb_6__3_/bottom_left_grid_pin_49_ cbx_6__3_/bottom_grid_pin_0_
+ cbx_6__3_/bottom_grid_pin_10_ cbx_6__3_/bottom_grid_pin_11_ cbx_6__3_/bottom_grid_pin_12_
+ cbx_6__3_/bottom_grid_pin_13_ cbx_6__3_/bottom_grid_pin_14_ cbx_6__3_/bottom_grid_pin_15_
+ cbx_6__3_/bottom_grid_pin_1_ cbx_6__3_/bottom_grid_pin_2_ cbx_6__3_/REGOUT_FEEDTHROUGH
+ grid_clb_6__3_/top_width_0_height_0__pin_33_ sb_6__3_/left_bottom_grid_pin_34_ sb_5__3_/right_bottom_grid_pin_34_
+ sb_6__3_/left_bottom_grid_pin_35_ sb_5__3_/right_bottom_grid_pin_35_ sb_6__3_/left_bottom_grid_pin_36_
+ sb_5__3_/right_bottom_grid_pin_36_ sb_6__3_/left_bottom_grid_pin_37_ sb_5__3_/right_bottom_grid_pin_37_
+ sb_6__3_/left_bottom_grid_pin_38_ sb_5__3_/right_bottom_grid_pin_38_ sb_6__3_/left_bottom_grid_pin_39_
+ sb_5__3_/right_bottom_grid_pin_39_ cbx_6__3_/bottom_grid_pin_3_ sb_6__3_/left_bottom_grid_pin_40_
+ sb_5__3_/right_bottom_grid_pin_40_ sb_6__3_/left_bottom_grid_pin_41_ sb_5__3_/right_bottom_grid_pin_41_
+ cbx_6__3_/bottom_grid_pin_4_ cbx_6__3_/bottom_grid_pin_5_ cbx_6__3_/bottom_grid_pin_6_
+ cbx_6__3_/bottom_grid_pin_7_ cbx_6__3_/bottom_grid_pin_8_ cbx_6__3_/bottom_grid_pin_9_
+ grid_clb
Xcbx_4__0_ IO_ISOL_N sb_3__0_/SC_OUT_TOP cbx_4__0_/SC_IN_TOP cbx_4__0_/SC_OUT_BOT
+ cbx_4__0_/SC_OUT_TOP VGND VPWR cbx_4__0_/bottom_grid_pin_0_ cbx_4__0_/bottom_grid_pin_10_
+ cbx_4__0_/bottom_grid_pin_12_ cbx_4__0_/bottom_grid_pin_14_ cbx_4__0_/bottom_grid_pin_16_
+ cbx_4__0_/bottom_grid_pin_2_ cbx_4__0_/bottom_grid_pin_4_ cbx_4__0_/bottom_grid_pin_6_
+ cbx_4__0_/bottom_grid_pin_8_ sb_4__0_/ccff_tail sb_3__0_/ccff_head cbx_4__0_/chanx_left_in[0]
+ cbx_4__0_/chanx_left_in[10] cbx_4__0_/chanx_left_in[11] cbx_4__0_/chanx_left_in[12]
+ cbx_4__0_/chanx_left_in[13] cbx_4__0_/chanx_left_in[14] cbx_4__0_/chanx_left_in[15]
+ cbx_4__0_/chanx_left_in[16] cbx_4__0_/chanx_left_in[17] cbx_4__0_/chanx_left_in[18]
+ cbx_4__0_/chanx_left_in[19] cbx_4__0_/chanx_left_in[1] cbx_4__0_/chanx_left_in[2]
+ cbx_4__0_/chanx_left_in[3] cbx_4__0_/chanx_left_in[4] cbx_4__0_/chanx_left_in[5]
+ cbx_4__0_/chanx_left_in[6] cbx_4__0_/chanx_left_in[7] cbx_4__0_/chanx_left_in[8]
+ cbx_4__0_/chanx_left_in[9] sb_3__0_/chanx_right_in[0] sb_3__0_/chanx_right_in[10]
+ sb_3__0_/chanx_right_in[11] sb_3__0_/chanx_right_in[12] sb_3__0_/chanx_right_in[13]
+ sb_3__0_/chanx_right_in[14] sb_3__0_/chanx_right_in[15] sb_3__0_/chanx_right_in[16]
+ sb_3__0_/chanx_right_in[17] sb_3__0_/chanx_right_in[18] sb_3__0_/chanx_right_in[19]
+ sb_3__0_/chanx_right_in[1] sb_3__0_/chanx_right_in[2] sb_3__0_/chanx_right_in[3]
+ sb_3__0_/chanx_right_in[4] sb_3__0_/chanx_right_in[5] sb_3__0_/chanx_right_in[6]
+ sb_3__0_/chanx_right_in[7] sb_3__0_/chanx_right_in[8] sb_3__0_/chanx_right_in[9]
+ sb_4__0_/chanx_left_out[0] sb_4__0_/chanx_left_out[10] sb_4__0_/chanx_left_out[11]
+ sb_4__0_/chanx_left_out[12] sb_4__0_/chanx_left_out[13] sb_4__0_/chanx_left_out[14]
+ sb_4__0_/chanx_left_out[15] sb_4__0_/chanx_left_out[16] sb_4__0_/chanx_left_out[17]
+ sb_4__0_/chanx_left_out[18] sb_4__0_/chanx_left_out[19] sb_4__0_/chanx_left_out[1]
+ sb_4__0_/chanx_left_out[2] sb_4__0_/chanx_left_out[3] sb_4__0_/chanx_left_out[4]
+ sb_4__0_/chanx_left_out[5] sb_4__0_/chanx_left_out[6] sb_4__0_/chanx_left_out[7]
+ sb_4__0_/chanx_left_out[8] sb_4__0_/chanx_left_out[9] sb_4__0_/chanx_left_in[0]
+ sb_4__0_/chanx_left_in[10] sb_4__0_/chanx_left_in[11] sb_4__0_/chanx_left_in[12]
+ sb_4__0_/chanx_left_in[13] sb_4__0_/chanx_left_in[14] sb_4__0_/chanx_left_in[15]
+ sb_4__0_/chanx_left_in[16] sb_4__0_/chanx_left_in[17] sb_4__0_/chanx_left_in[18]
+ sb_4__0_/chanx_left_in[19] sb_4__0_/chanx_left_in[1] sb_4__0_/chanx_left_in[2] sb_4__0_/chanx_left_in[3]
+ sb_4__0_/chanx_left_in[4] sb_4__0_/chanx_left_in[5] sb_4__0_/chanx_left_in[6] sb_4__0_/chanx_left_in[7]
+ sb_4__0_/chanx_left_in[8] sb_4__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60] cbx_4__0_/prog_clk_0_N_in
+ cbx_4__0_/prog_clk_0_W_out cbx_4__0_/bottom_grid_pin_0_ cbx_4__0_/bottom_grid_pin_10_
+ sb_4__0_/left_bottom_grid_pin_11_ sb_3__0_/right_bottom_grid_pin_11_ cbx_4__0_/bottom_grid_pin_12_
+ sb_4__0_/left_bottom_grid_pin_13_ sb_3__0_/right_bottom_grid_pin_13_ cbx_4__0_/bottom_grid_pin_14_
+ sb_4__0_/left_bottom_grid_pin_15_ sb_3__0_/right_bottom_grid_pin_15_ cbx_4__0_/bottom_grid_pin_16_
+ sb_4__0_/left_bottom_grid_pin_17_ sb_3__0_/right_bottom_grid_pin_17_ sb_4__0_/left_bottom_grid_pin_1_
+ sb_3__0_/right_bottom_grid_pin_1_ cbx_4__0_/bottom_grid_pin_2_ sb_4__0_/left_bottom_grid_pin_3_
+ sb_3__0_/right_bottom_grid_pin_3_ cbx_4__0_/bottom_grid_pin_4_ sb_4__0_/left_bottom_grid_pin_5_
+ sb_3__0_/right_bottom_grid_pin_5_ cbx_4__0_/bottom_grid_pin_6_ sb_4__0_/left_bottom_grid_pin_7_
+ sb_3__0_/right_bottom_grid_pin_7_ cbx_4__0_/bottom_grid_pin_8_ sb_4__0_/left_bottom_grid_pin_9_
+ sb_3__0_/right_bottom_grid_pin_9_ cbx_1__0_
Xsb_1__2_ sb_1__2_/Test_en_N_out sb_1__2_/Test_en_S_in VGND VPWR sb_1__2_/bottom_left_grid_pin_42_
+ sb_1__2_/bottom_left_grid_pin_43_ sb_1__2_/bottom_left_grid_pin_44_ sb_1__2_/bottom_left_grid_pin_45_
+ sb_1__2_/bottom_left_grid_pin_46_ sb_1__2_/bottom_left_grid_pin_47_ sb_1__2_/bottom_left_grid_pin_48_
+ sb_1__2_/bottom_left_grid_pin_49_ sb_1__2_/ccff_head sb_1__2_/ccff_tail sb_1__2_/chanx_left_in[0]
+ sb_1__2_/chanx_left_in[10] sb_1__2_/chanx_left_in[11] sb_1__2_/chanx_left_in[12]
+ sb_1__2_/chanx_left_in[13] sb_1__2_/chanx_left_in[14] sb_1__2_/chanx_left_in[15]
+ sb_1__2_/chanx_left_in[16] sb_1__2_/chanx_left_in[17] sb_1__2_/chanx_left_in[18]
+ sb_1__2_/chanx_left_in[19] sb_1__2_/chanx_left_in[1] sb_1__2_/chanx_left_in[2] sb_1__2_/chanx_left_in[3]
+ sb_1__2_/chanx_left_in[4] sb_1__2_/chanx_left_in[5] sb_1__2_/chanx_left_in[6] sb_1__2_/chanx_left_in[7]
+ sb_1__2_/chanx_left_in[8] sb_1__2_/chanx_left_in[9] sb_1__2_/chanx_left_out[0] sb_1__2_/chanx_left_out[10]
+ sb_1__2_/chanx_left_out[11] sb_1__2_/chanx_left_out[12] sb_1__2_/chanx_left_out[13]
+ sb_1__2_/chanx_left_out[14] sb_1__2_/chanx_left_out[15] sb_1__2_/chanx_left_out[16]
+ sb_1__2_/chanx_left_out[17] sb_1__2_/chanx_left_out[18] sb_1__2_/chanx_left_out[19]
+ sb_1__2_/chanx_left_out[1] sb_1__2_/chanx_left_out[2] sb_1__2_/chanx_left_out[3]
+ sb_1__2_/chanx_left_out[4] sb_1__2_/chanx_left_out[5] sb_1__2_/chanx_left_out[6]
+ sb_1__2_/chanx_left_out[7] sb_1__2_/chanx_left_out[8] sb_1__2_/chanx_left_out[9]
+ sb_1__2_/chanx_right_in[0] sb_1__2_/chanx_right_in[10] sb_1__2_/chanx_right_in[11]
+ sb_1__2_/chanx_right_in[12] sb_1__2_/chanx_right_in[13] sb_1__2_/chanx_right_in[14]
+ sb_1__2_/chanx_right_in[15] sb_1__2_/chanx_right_in[16] sb_1__2_/chanx_right_in[17]
+ sb_1__2_/chanx_right_in[18] sb_1__2_/chanx_right_in[19] sb_1__2_/chanx_right_in[1]
+ sb_1__2_/chanx_right_in[2] sb_1__2_/chanx_right_in[3] sb_1__2_/chanx_right_in[4]
+ sb_1__2_/chanx_right_in[5] sb_1__2_/chanx_right_in[6] sb_1__2_/chanx_right_in[7]
+ sb_1__2_/chanx_right_in[8] sb_1__2_/chanx_right_in[9] cbx_2__2_/chanx_left_in[0]
+ cbx_2__2_/chanx_left_in[10] cbx_2__2_/chanx_left_in[11] cbx_2__2_/chanx_left_in[12]
+ cbx_2__2_/chanx_left_in[13] cbx_2__2_/chanx_left_in[14] cbx_2__2_/chanx_left_in[15]
+ cbx_2__2_/chanx_left_in[16] cbx_2__2_/chanx_left_in[17] cbx_2__2_/chanx_left_in[18]
+ cbx_2__2_/chanx_left_in[19] cbx_2__2_/chanx_left_in[1] cbx_2__2_/chanx_left_in[2]
+ cbx_2__2_/chanx_left_in[3] cbx_2__2_/chanx_left_in[4] cbx_2__2_/chanx_left_in[5]
+ cbx_2__2_/chanx_left_in[6] cbx_2__2_/chanx_left_in[7] cbx_2__2_/chanx_left_in[8]
+ cbx_2__2_/chanx_left_in[9] cby_1__2_/chany_top_out[0] cby_1__2_/chany_top_out[10]
+ cby_1__2_/chany_top_out[11] cby_1__2_/chany_top_out[12] cby_1__2_/chany_top_out[13]
+ cby_1__2_/chany_top_out[14] cby_1__2_/chany_top_out[15] cby_1__2_/chany_top_out[16]
+ cby_1__2_/chany_top_out[17] cby_1__2_/chany_top_out[18] cby_1__2_/chany_top_out[19]
+ cby_1__2_/chany_top_out[1] cby_1__2_/chany_top_out[2] cby_1__2_/chany_top_out[3]
+ cby_1__2_/chany_top_out[4] cby_1__2_/chany_top_out[5] cby_1__2_/chany_top_out[6]
+ cby_1__2_/chany_top_out[7] cby_1__2_/chany_top_out[8] cby_1__2_/chany_top_out[9]
+ cby_1__2_/chany_top_in[0] cby_1__2_/chany_top_in[10] cby_1__2_/chany_top_in[11]
+ cby_1__2_/chany_top_in[12] cby_1__2_/chany_top_in[13] cby_1__2_/chany_top_in[14]
+ cby_1__2_/chany_top_in[15] cby_1__2_/chany_top_in[16] cby_1__2_/chany_top_in[17]
+ cby_1__2_/chany_top_in[18] cby_1__2_/chany_top_in[19] cby_1__2_/chany_top_in[1]
+ cby_1__2_/chany_top_in[2] cby_1__2_/chany_top_in[3] cby_1__2_/chany_top_in[4] cby_1__2_/chany_top_in[5]
+ cby_1__2_/chany_top_in[6] cby_1__2_/chany_top_in[7] cby_1__2_/chany_top_in[8] cby_1__2_/chany_top_in[9]
+ sb_1__2_/chany_top_in[0] sb_1__2_/chany_top_in[10] sb_1__2_/chany_top_in[11] sb_1__2_/chany_top_in[12]
+ sb_1__2_/chany_top_in[13] sb_1__2_/chany_top_in[14] sb_1__2_/chany_top_in[15] sb_1__2_/chany_top_in[16]
+ sb_1__2_/chany_top_in[17] sb_1__2_/chany_top_in[18] sb_1__2_/chany_top_in[19] sb_1__2_/chany_top_in[1]
+ sb_1__2_/chany_top_in[2] sb_1__2_/chany_top_in[3] sb_1__2_/chany_top_in[4] sb_1__2_/chany_top_in[5]
+ sb_1__2_/chany_top_in[6] sb_1__2_/chany_top_in[7] sb_1__2_/chany_top_in[8] sb_1__2_/chany_top_in[9]
+ sb_1__2_/chany_top_out[0] sb_1__2_/chany_top_out[10] sb_1__2_/chany_top_out[11]
+ sb_1__2_/chany_top_out[12] sb_1__2_/chany_top_out[13] sb_1__2_/chany_top_out[14]
+ sb_1__2_/chany_top_out[15] sb_1__2_/chany_top_out[16] sb_1__2_/chany_top_out[17]
+ sb_1__2_/chany_top_out[18] sb_1__2_/chany_top_out[19] sb_1__2_/chany_top_out[1]
+ sb_1__2_/chany_top_out[2] sb_1__2_/chany_top_out[3] sb_1__2_/chany_top_out[4] sb_1__2_/chany_top_out[5]
+ sb_1__2_/chany_top_out[6] sb_1__2_/chany_top_out[7] sb_1__2_/chany_top_out[8] sb_1__2_/chany_top_out[9]
+ sb_1__2_/clk_1_E_out sb_1__2_/clk_1_N_in sb_1__2_/clk_1_W_out sb_1__2_/clk_2_E_out
+ sb_1__2_/clk_2_N_in sb_1__2_/clk_2_N_out sb_1__2_/clk_2_S_out sb_1__2_/clk_2_W_out
+ sb_1__2_/clk_3_E_out sb_1__2_/clk_3_N_in sb_1__2_/clk_3_N_out sb_1__2_/clk_3_S_out
+ sb_1__2_/clk_3_W_out sb_1__2_/left_bottom_grid_pin_34_ sb_1__2_/left_bottom_grid_pin_35_
+ sb_1__2_/left_bottom_grid_pin_36_ sb_1__2_/left_bottom_grid_pin_37_ sb_1__2_/left_bottom_grid_pin_38_
+ sb_1__2_/left_bottom_grid_pin_39_ sb_1__2_/left_bottom_grid_pin_40_ sb_1__2_/left_bottom_grid_pin_41_
+ sb_1__2_/prog_clk_0_N_in sb_1__2_/prog_clk_1_E_out sb_1__2_/prog_clk_1_N_in sb_1__2_/prog_clk_1_W_out
+ sb_1__2_/prog_clk_2_E_out sb_1__2_/prog_clk_2_N_in sb_1__2_/prog_clk_2_N_out sb_1__2_/prog_clk_2_S_out
+ sb_1__2_/prog_clk_2_W_out sb_1__2_/prog_clk_3_E_out sb_1__2_/prog_clk_3_N_in sb_1__2_/prog_clk_3_N_out
+ sb_1__2_/prog_clk_3_S_out sb_1__2_/prog_clk_3_W_out sb_1__2_/right_bottom_grid_pin_34_
+ sb_1__2_/right_bottom_grid_pin_35_ sb_1__2_/right_bottom_grid_pin_36_ sb_1__2_/right_bottom_grid_pin_37_
+ sb_1__2_/right_bottom_grid_pin_38_ sb_1__2_/right_bottom_grid_pin_39_ sb_1__2_/right_bottom_grid_pin_40_
+ sb_1__2_/right_bottom_grid_pin_41_ sb_1__2_/top_left_grid_pin_42_ sb_1__2_/top_left_grid_pin_43_
+ sb_1__2_/top_left_grid_pin_44_ sb_1__2_/top_left_grid_pin_45_ sb_1__2_/top_left_grid_pin_46_
+ sb_1__2_/top_left_grid_pin_47_ sb_1__2_/top_left_grid_pin_48_ sb_1__2_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_7__1_ cby_7__1_/Test_en_W_in cby_7__1_/Test_en_E_out cby_7__1_/Test_en_N_out
+ cby_7__1_/Test_en_W_in cby_7__1_/Test_en_W_in cby_7__1_/Test_en_W_out VGND VPWR
+ cby_7__1_/ccff_head cby_7__1_/ccff_tail sb_7__0_/chany_top_out[0] sb_7__0_/chany_top_out[10]
+ sb_7__0_/chany_top_out[11] sb_7__0_/chany_top_out[12] sb_7__0_/chany_top_out[13]
+ sb_7__0_/chany_top_out[14] sb_7__0_/chany_top_out[15] sb_7__0_/chany_top_out[16]
+ sb_7__0_/chany_top_out[17] sb_7__0_/chany_top_out[18] sb_7__0_/chany_top_out[19]
+ sb_7__0_/chany_top_out[1] sb_7__0_/chany_top_out[2] sb_7__0_/chany_top_out[3] sb_7__0_/chany_top_out[4]
+ sb_7__0_/chany_top_out[5] sb_7__0_/chany_top_out[6] sb_7__0_/chany_top_out[7] sb_7__0_/chany_top_out[8]
+ sb_7__0_/chany_top_out[9] sb_7__0_/chany_top_in[0] sb_7__0_/chany_top_in[10] sb_7__0_/chany_top_in[11]
+ sb_7__0_/chany_top_in[12] sb_7__0_/chany_top_in[13] sb_7__0_/chany_top_in[14] sb_7__0_/chany_top_in[15]
+ sb_7__0_/chany_top_in[16] sb_7__0_/chany_top_in[17] sb_7__0_/chany_top_in[18] sb_7__0_/chany_top_in[19]
+ sb_7__0_/chany_top_in[1] sb_7__0_/chany_top_in[2] sb_7__0_/chany_top_in[3] sb_7__0_/chany_top_in[4]
+ sb_7__0_/chany_top_in[5] sb_7__0_/chany_top_in[6] sb_7__0_/chany_top_in[7] sb_7__0_/chany_top_in[8]
+ sb_7__0_/chany_top_in[9] cby_7__1_/chany_top_in[0] cby_7__1_/chany_top_in[10] cby_7__1_/chany_top_in[11]
+ cby_7__1_/chany_top_in[12] cby_7__1_/chany_top_in[13] cby_7__1_/chany_top_in[14]
+ cby_7__1_/chany_top_in[15] cby_7__1_/chany_top_in[16] cby_7__1_/chany_top_in[17]
+ cby_7__1_/chany_top_in[18] cby_7__1_/chany_top_in[19] cby_7__1_/chany_top_in[1]
+ cby_7__1_/chany_top_in[2] cby_7__1_/chany_top_in[3] cby_7__1_/chany_top_in[4] cby_7__1_/chany_top_in[5]
+ cby_7__1_/chany_top_in[6] cby_7__1_/chany_top_in[7] cby_7__1_/chany_top_in[8] cby_7__1_/chany_top_in[9]
+ cby_7__1_/chany_top_out[0] cby_7__1_/chany_top_out[10] cby_7__1_/chany_top_out[11]
+ cby_7__1_/chany_top_out[12] cby_7__1_/chany_top_out[13] cby_7__1_/chany_top_out[14]
+ cby_7__1_/chany_top_out[15] cby_7__1_/chany_top_out[16] cby_7__1_/chany_top_out[17]
+ cby_7__1_/chany_top_out[18] cby_7__1_/chany_top_out[19] cby_7__1_/chany_top_out[1]
+ cby_7__1_/chany_top_out[2] cby_7__1_/chany_top_out[3] cby_7__1_/chany_top_out[4]
+ cby_7__1_/chany_top_out[5] cby_7__1_/chany_top_out[6] cby_7__1_/chany_top_out[7]
+ cby_7__1_/chany_top_out[8] cby_7__1_/chany_top_out[9] cby_7__1_/clk_2_N_out cby_7__1_/clk_2_S_in
+ cby_7__1_/clk_2_S_out cby_7__1_/clk_3_N_out cby_7__1_/clk_3_S_in cby_7__1_/clk_3_S_out
+ cby_7__1_/left_grid_pin_16_ cby_7__1_/left_grid_pin_17_ cby_7__1_/left_grid_pin_18_
+ cby_7__1_/left_grid_pin_19_ cby_7__1_/left_grid_pin_20_ cby_7__1_/left_grid_pin_21_
+ cby_7__1_/left_grid_pin_22_ cby_7__1_/left_grid_pin_23_ cby_7__1_/left_grid_pin_24_
+ cby_7__1_/left_grid_pin_25_ cby_7__1_/left_grid_pin_26_ cby_7__1_/left_grid_pin_27_
+ cby_7__1_/left_grid_pin_28_ cby_7__1_/left_grid_pin_29_ cby_7__1_/left_grid_pin_30_
+ cby_7__1_/left_grid_pin_31_ cby_7__1_/prog_clk_0_N_out sb_7__0_/prog_clk_0_N_in
+ cby_7__1_/prog_clk_0_W_in cby_7__1_/prog_clk_2_N_out cby_7__1_/prog_clk_2_S_in cby_7__1_/prog_clk_2_S_out
+ cby_7__1_/prog_clk_3_N_out cby_7__1_/prog_clk_3_S_in cby_7__1_/prog_clk_3_S_out
+ cby_1__1_
Xcby_0__6_ IO_ISOL_N VGND VPWR sb_0__6_/ccff_tail cby_0__6_/ccff_tail sb_0__5_/chany_top_out[0]
+ sb_0__5_/chany_top_out[10] sb_0__5_/chany_top_out[11] sb_0__5_/chany_top_out[12]
+ sb_0__5_/chany_top_out[13] sb_0__5_/chany_top_out[14] sb_0__5_/chany_top_out[15]
+ sb_0__5_/chany_top_out[16] sb_0__5_/chany_top_out[17] sb_0__5_/chany_top_out[18]
+ sb_0__5_/chany_top_out[19] sb_0__5_/chany_top_out[1] sb_0__5_/chany_top_out[2] sb_0__5_/chany_top_out[3]
+ sb_0__5_/chany_top_out[4] sb_0__5_/chany_top_out[5] sb_0__5_/chany_top_out[6] sb_0__5_/chany_top_out[7]
+ sb_0__5_/chany_top_out[8] sb_0__5_/chany_top_out[9] sb_0__5_/chany_top_in[0] sb_0__5_/chany_top_in[10]
+ sb_0__5_/chany_top_in[11] sb_0__5_/chany_top_in[12] sb_0__5_/chany_top_in[13] sb_0__5_/chany_top_in[14]
+ sb_0__5_/chany_top_in[15] sb_0__5_/chany_top_in[16] sb_0__5_/chany_top_in[17] sb_0__5_/chany_top_in[18]
+ sb_0__5_/chany_top_in[19] sb_0__5_/chany_top_in[1] sb_0__5_/chany_top_in[2] sb_0__5_/chany_top_in[3]
+ sb_0__5_/chany_top_in[4] sb_0__5_/chany_top_in[5] sb_0__5_/chany_top_in[6] sb_0__5_/chany_top_in[7]
+ sb_0__5_/chany_top_in[8] sb_0__5_/chany_top_in[9] cby_0__6_/chany_top_in[0] cby_0__6_/chany_top_in[10]
+ cby_0__6_/chany_top_in[11] cby_0__6_/chany_top_in[12] cby_0__6_/chany_top_in[13]
+ cby_0__6_/chany_top_in[14] cby_0__6_/chany_top_in[15] cby_0__6_/chany_top_in[16]
+ cby_0__6_/chany_top_in[17] cby_0__6_/chany_top_in[18] cby_0__6_/chany_top_in[19]
+ cby_0__6_/chany_top_in[1] cby_0__6_/chany_top_in[2] cby_0__6_/chany_top_in[3] cby_0__6_/chany_top_in[4]
+ cby_0__6_/chany_top_in[5] cby_0__6_/chany_top_in[6] cby_0__6_/chany_top_in[7] cby_0__6_/chany_top_in[8]
+ cby_0__6_/chany_top_in[9] cby_0__6_/chany_top_out[0] cby_0__6_/chany_top_out[10]
+ cby_0__6_/chany_top_out[11] cby_0__6_/chany_top_out[12] cby_0__6_/chany_top_out[13]
+ cby_0__6_/chany_top_out[14] cby_0__6_/chany_top_out[15] cby_0__6_/chany_top_out[16]
+ cby_0__6_/chany_top_out[17] cby_0__6_/chany_top_out[18] cby_0__6_/chany_top_out[19]
+ cby_0__6_/chany_top_out[1] cby_0__6_/chany_top_out[2] cby_0__6_/chany_top_out[3]
+ cby_0__6_/chany_top_out[4] cby_0__6_/chany_top_out[5] cby_0__6_/chany_top_out[6]
+ cby_0__6_/chany_top_out[7] cby_0__6_/chany_top_out[8] cby_0__6_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
+ cby_0__6_/left_grid_pin_0_ cby_0__6_/prog_clk_0_E_in cby_0__6_/left_grid_pin_0_
+ sb_0__5_/top_left_grid_pin_1_ sb_0__6_/bottom_left_grid_pin_1_ cby_0__1_
Xgrid_clb_6__2_ cbx_6__1_/SC_OUT_TOP grid_clb_6__2_/SC_OUT_BOT cbx_6__2_/SC_IN_BOT
+ cby_5__2_/Test_en_E_out cby_6__2_/Test_en_W_in cby_5__2_/Test_en_E_out grid_clb_6__2_/Test_en_W_out
+ VGND VPWR cbx_6__1_/REGIN_FEEDTHROUGH grid_clb_6__2_/bottom_width_0_height_0__pin_51_
+ cby_5__2_/ccff_tail cby_6__2_/ccff_head cbx_6__1_/clk_1_N_out cbx_6__1_/clk_1_N_out
+ cby_6__2_/prog_clk_0_W_in cbx_6__1_/prog_clk_1_N_out grid_clb_6__2_/prog_clk_0_N_out
+ cbx_6__1_/prog_clk_1_N_out cbx_6__1_/prog_clk_0_N_in grid_clb_6__2_/prog_clk_0_W_out
+ cby_6__2_/left_grid_pin_16_ cby_6__2_/left_grid_pin_17_ cby_6__2_/left_grid_pin_18_
+ cby_6__2_/left_grid_pin_19_ cby_6__2_/left_grid_pin_20_ cby_6__2_/left_grid_pin_21_
+ cby_6__2_/left_grid_pin_22_ cby_6__2_/left_grid_pin_23_ cby_6__2_/left_grid_pin_24_
+ cby_6__2_/left_grid_pin_25_ cby_6__2_/left_grid_pin_26_ cby_6__2_/left_grid_pin_27_
+ cby_6__2_/left_grid_pin_28_ cby_6__2_/left_grid_pin_29_ cby_6__2_/left_grid_pin_30_
+ cby_6__2_/left_grid_pin_31_ sb_6__1_/top_left_grid_pin_42_ sb_6__2_/bottom_left_grid_pin_42_
+ sb_6__1_/top_left_grid_pin_43_ sb_6__2_/bottom_left_grid_pin_43_ sb_6__1_/top_left_grid_pin_44_
+ sb_6__2_/bottom_left_grid_pin_44_ sb_6__1_/top_left_grid_pin_45_ sb_6__2_/bottom_left_grid_pin_45_
+ sb_6__1_/top_left_grid_pin_46_ sb_6__2_/bottom_left_grid_pin_46_ sb_6__1_/top_left_grid_pin_47_
+ sb_6__2_/bottom_left_grid_pin_47_ sb_6__1_/top_left_grid_pin_48_ sb_6__2_/bottom_left_grid_pin_48_
+ sb_6__1_/top_left_grid_pin_49_ sb_6__2_/bottom_left_grid_pin_49_ cbx_6__2_/bottom_grid_pin_0_
+ cbx_6__2_/bottom_grid_pin_10_ cbx_6__2_/bottom_grid_pin_11_ cbx_6__2_/bottom_grid_pin_12_
+ cbx_6__2_/bottom_grid_pin_13_ cbx_6__2_/bottom_grid_pin_14_ cbx_6__2_/bottom_grid_pin_15_
+ cbx_6__2_/bottom_grid_pin_1_ cbx_6__2_/bottom_grid_pin_2_ cbx_6__2_/REGOUT_FEEDTHROUGH
+ grid_clb_6__2_/top_width_0_height_0__pin_33_ sb_6__2_/left_bottom_grid_pin_34_ sb_5__2_/right_bottom_grid_pin_34_
+ sb_6__2_/left_bottom_grid_pin_35_ sb_5__2_/right_bottom_grid_pin_35_ sb_6__2_/left_bottom_grid_pin_36_
+ sb_5__2_/right_bottom_grid_pin_36_ sb_6__2_/left_bottom_grid_pin_37_ sb_5__2_/right_bottom_grid_pin_37_
+ sb_6__2_/left_bottom_grid_pin_38_ sb_5__2_/right_bottom_grid_pin_38_ sb_6__2_/left_bottom_grid_pin_39_
+ sb_5__2_/right_bottom_grid_pin_39_ cbx_6__2_/bottom_grid_pin_3_ sb_6__2_/left_bottom_grid_pin_40_
+ sb_5__2_/right_bottom_grid_pin_40_ sb_6__2_/left_bottom_grid_pin_41_ sb_5__2_/right_bottom_grid_pin_41_
+ cbx_6__2_/bottom_grid_pin_4_ cbx_6__2_/bottom_grid_pin_5_ cbx_6__2_/bottom_grid_pin_6_
+ cbx_6__2_/bottom_grid_pin_7_ cbx_6__2_/bottom_grid_pin_8_ cbx_6__2_/bottom_grid_pin_9_
+ grid_clb
Xcbx_7__2_ cbx_7__2_/REGIN_FEEDTHROUGH cbx_7__2_/REGOUT_FEEDTHROUGH cbx_7__2_/SC_IN_BOT
+ cbx_7__2_/SC_IN_TOP cbx_7__2_/SC_OUT_BOT cbx_7__2_/SC_OUT_TOP VGND VPWR cbx_7__2_/bottom_grid_pin_0_
+ cbx_7__2_/bottom_grid_pin_10_ cbx_7__2_/bottom_grid_pin_11_ cbx_7__2_/bottom_grid_pin_12_
+ cbx_7__2_/bottom_grid_pin_13_ cbx_7__2_/bottom_grid_pin_14_ cbx_7__2_/bottom_grid_pin_15_
+ cbx_7__2_/bottom_grid_pin_1_ cbx_7__2_/bottom_grid_pin_2_ cbx_7__2_/bottom_grid_pin_3_
+ cbx_7__2_/bottom_grid_pin_4_ cbx_7__2_/bottom_grid_pin_5_ cbx_7__2_/bottom_grid_pin_6_
+ cbx_7__2_/bottom_grid_pin_7_ cbx_7__2_/bottom_grid_pin_8_ cbx_7__2_/bottom_grid_pin_9_
+ sb_7__2_/ccff_tail sb_6__2_/ccff_head cbx_7__2_/chanx_left_in[0] cbx_7__2_/chanx_left_in[10]
+ cbx_7__2_/chanx_left_in[11] cbx_7__2_/chanx_left_in[12] cbx_7__2_/chanx_left_in[13]
+ cbx_7__2_/chanx_left_in[14] cbx_7__2_/chanx_left_in[15] cbx_7__2_/chanx_left_in[16]
+ cbx_7__2_/chanx_left_in[17] cbx_7__2_/chanx_left_in[18] cbx_7__2_/chanx_left_in[19]
+ cbx_7__2_/chanx_left_in[1] cbx_7__2_/chanx_left_in[2] cbx_7__2_/chanx_left_in[3]
+ cbx_7__2_/chanx_left_in[4] cbx_7__2_/chanx_left_in[5] cbx_7__2_/chanx_left_in[6]
+ cbx_7__2_/chanx_left_in[7] cbx_7__2_/chanx_left_in[8] cbx_7__2_/chanx_left_in[9]
+ sb_6__2_/chanx_right_in[0] sb_6__2_/chanx_right_in[10] sb_6__2_/chanx_right_in[11]
+ sb_6__2_/chanx_right_in[12] sb_6__2_/chanx_right_in[13] sb_6__2_/chanx_right_in[14]
+ sb_6__2_/chanx_right_in[15] sb_6__2_/chanx_right_in[16] sb_6__2_/chanx_right_in[17]
+ sb_6__2_/chanx_right_in[18] sb_6__2_/chanx_right_in[19] sb_6__2_/chanx_right_in[1]
+ sb_6__2_/chanx_right_in[2] sb_6__2_/chanx_right_in[3] sb_6__2_/chanx_right_in[4]
+ sb_6__2_/chanx_right_in[5] sb_6__2_/chanx_right_in[6] sb_6__2_/chanx_right_in[7]
+ sb_6__2_/chanx_right_in[8] sb_6__2_/chanx_right_in[9] sb_7__2_/chanx_left_out[0]
+ sb_7__2_/chanx_left_out[10] sb_7__2_/chanx_left_out[11] sb_7__2_/chanx_left_out[12]
+ sb_7__2_/chanx_left_out[13] sb_7__2_/chanx_left_out[14] sb_7__2_/chanx_left_out[15]
+ sb_7__2_/chanx_left_out[16] sb_7__2_/chanx_left_out[17] sb_7__2_/chanx_left_out[18]
+ sb_7__2_/chanx_left_out[19] sb_7__2_/chanx_left_out[1] sb_7__2_/chanx_left_out[2]
+ sb_7__2_/chanx_left_out[3] sb_7__2_/chanx_left_out[4] sb_7__2_/chanx_left_out[5]
+ sb_7__2_/chanx_left_out[6] sb_7__2_/chanx_left_out[7] sb_7__2_/chanx_left_out[8]
+ sb_7__2_/chanx_left_out[9] sb_7__2_/chanx_left_in[0] sb_7__2_/chanx_left_in[10]
+ sb_7__2_/chanx_left_in[11] sb_7__2_/chanx_left_in[12] sb_7__2_/chanx_left_in[13]
+ sb_7__2_/chanx_left_in[14] sb_7__2_/chanx_left_in[15] sb_7__2_/chanx_left_in[16]
+ sb_7__2_/chanx_left_in[17] sb_7__2_/chanx_left_in[18] sb_7__2_/chanx_left_in[19]
+ sb_7__2_/chanx_left_in[1] sb_7__2_/chanx_left_in[2] sb_7__2_/chanx_left_in[3] sb_7__2_/chanx_left_in[4]
+ sb_7__2_/chanx_left_in[5] sb_7__2_/chanx_left_in[6] sb_7__2_/chanx_left_in[7] sb_7__2_/chanx_left_in[8]
+ sb_7__2_/chanx_left_in[9] cbx_7__2_/clk_1_N_out cbx_7__2_/clk_1_S_out cbx_7__2_/clk_1_W_in
+ sb_7__2_/clk_2_N_in sb_6__2_/clk_2_E_out cbx_7__2_/clk_2_W_out cbx_7__2_/clk_3_E_out
+ cbx_7__2_/clk_3_W_in cbx_7__2_/clk_3_W_out cbx_7__2_/prog_clk_0_N_in cbx_7__2_/prog_clk_0_W_out
+ cbx_7__2_/prog_clk_1_N_out cbx_7__2_/prog_clk_1_S_out cbx_7__2_/prog_clk_1_W_in
+ sb_7__2_/prog_clk_2_N_in sb_6__2_/prog_clk_2_E_out cbx_7__2_/prog_clk_2_W_out cbx_7__2_/prog_clk_3_E_out
+ cbx_7__2_/prog_clk_3_W_in cbx_7__2_/prog_clk_3_W_out cbx_1__1_
Xsb_7__7_ sb_7__7_/Test_en_N_out sb_7__7_/Test_en_S_in VGND VPWR sb_7__7_/bottom_left_grid_pin_42_
+ sb_7__7_/bottom_left_grid_pin_43_ sb_7__7_/bottom_left_grid_pin_44_ sb_7__7_/bottom_left_grid_pin_45_
+ sb_7__7_/bottom_left_grid_pin_46_ sb_7__7_/bottom_left_grid_pin_47_ sb_7__7_/bottom_left_grid_pin_48_
+ sb_7__7_/bottom_left_grid_pin_49_ sb_7__7_/ccff_head sb_7__7_/ccff_tail sb_7__7_/chanx_left_in[0]
+ sb_7__7_/chanx_left_in[10] sb_7__7_/chanx_left_in[11] sb_7__7_/chanx_left_in[12]
+ sb_7__7_/chanx_left_in[13] sb_7__7_/chanx_left_in[14] sb_7__7_/chanx_left_in[15]
+ sb_7__7_/chanx_left_in[16] sb_7__7_/chanx_left_in[17] sb_7__7_/chanx_left_in[18]
+ sb_7__7_/chanx_left_in[19] sb_7__7_/chanx_left_in[1] sb_7__7_/chanx_left_in[2] sb_7__7_/chanx_left_in[3]
+ sb_7__7_/chanx_left_in[4] sb_7__7_/chanx_left_in[5] sb_7__7_/chanx_left_in[6] sb_7__7_/chanx_left_in[7]
+ sb_7__7_/chanx_left_in[8] sb_7__7_/chanx_left_in[9] sb_7__7_/chanx_left_out[0] sb_7__7_/chanx_left_out[10]
+ sb_7__7_/chanx_left_out[11] sb_7__7_/chanx_left_out[12] sb_7__7_/chanx_left_out[13]
+ sb_7__7_/chanx_left_out[14] sb_7__7_/chanx_left_out[15] sb_7__7_/chanx_left_out[16]
+ sb_7__7_/chanx_left_out[17] sb_7__7_/chanx_left_out[18] sb_7__7_/chanx_left_out[19]
+ sb_7__7_/chanx_left_out[1] sb_7__7_/chanx_left_out[2] sb_7__7_/chanx_left_out[3]
+ sb_7__7_/chanx_left_out[4] sb_7__7_/chanx_left_out[5] sb_7__7_/chanx_left_out[6]
+ sb_7__7_/chanx_left_out[7] sb_7__7_/chanx_left_out[8] sb_7__7_/chanx_left_out[9]
+ sb_7__7_/chanx_right_in[0] sb_7__7_/chanx_right_in[10] sb_7__7_/chanx_right_in[11]
+ sb_7__7_/chanx_right_in[12] sb_7__7_/chanx_right_in[13] sb_7__7_/chanx_right_in[14]
+ sb_7__7_/chanx_right_in[15] sb_7__7_/chanx_right_in[16] sb_7__7_/chanx_right_in[17]
+ sb_7__7_/chanx_right_in[18] sb_7__7_/chanx_right_in[19] sb_7__7_/chanx_right_in[1]
+ sb_7__7_/chanx_right_in[2] sb_7__7_/chanx_right_in[3] sb_7__7_/chanx_right_in[4]
+ sb_7__7_/chanx_right_in[5] sb_7__7_/chanx_right_in[6] sb_7__7_/chanx_right_in[7]
+ sb_7__7_/chanx_right_in[8] sb_7__7_/chanx_right_in[9] cbx_8__7_/chanx_left_in[0]
+ cbx_8__7_/chanx_left_in[10] cbx_8__7_/chanx_left_in[11] cbx_8__7_/chanx_left_in[12]
+ cbx_8__7_/chanx_left_in[13] cbx_8__7_/chanx_left_in[14] cbx_8__7_/chanx_left_in[15]
+ cbx_8__7_/chanx_left_in[16] cbx_8__7_/chanx_left_in[17] cbx_8__7_/chanx_left_in[18]
+ cbx_8__7_/chanx_left_in[19] cbx_8__7_/chanx_left_in[1] cbx_8__7_/chanx_left_in[2]
+ cbx_8__7_/chanx_left_in[3] cbx_8__7_/chanx_left_in[4] cbx_8__7_/chanx_left_in[5]
+ cbx_8__7_/chanx_left_in[6] cbx_8__7_/chanx_left_in[7] cbx_8__7_/chanx_left_in[8]
+ cbx_8__7_/chanx_left_in[9] cby_7__7_/chany_top_out[0] cby_7__7_/chany_top_out[10]
+ cby_7__7_/chany_top_out[11] cby_7__7_/chany_top_out[12] cby_7__7_/chany_top_out[13]
+ cby_7__7_/chany_top_out[14] cby_7__7_/chany_top_out[15] cby_7__7_/chany_top_out[16]
+ cby_7__7_/chany_top_out[17] cby_7__7_/chany_top_out[18] cby_7__7_/chany_top_out[19]
+ cby_7__7_/chany_top_out[1] cby_7__7_/chany_top_out[2] cby_7__7_/chany_top_out[3]
+ cby_7__7_/chany_top_out[4] cby_7__7_/chany_top_out[5] cby_7__7_/chany_top_out[6]
+ cby_7__7_/chany_top_out[7] cby_7__7_/chany_top_out[8] cby_7__7_/chany_top_out[9]
+ cby_7__7_/chany_top_in[0] cby_7__7_/chany_top_in[10] cby_7__7_/chany_top_in[11]
+ cby_7__7_/chany_top_in[12] cby_7__7_/chany_top_in[13] cby_7__7_/chany_top_in[14]
+ cby_7__7_/chany_top_in[15] cby_7__7_/chany_top_in[16] cby_7__7_/chany_top_in[17]
+ cby_7__7_/chany_top_in[18] cby_7__7_/chany_top_in[19] cby_7__7_/chany_top_in[1]
+ cby_7__7_/chany_top_in[2] cby_7__7_/chany_top_in[3] cby_7__7_/chany_top_in[4] cby_7__7_/chany_top_in[5]
+ cby_7__7_/chany_top_in[6] cby_7__7_/chany_top_in[7] cby_7__7_/chany_top_in[8] cby_7__7_/chany_top_in[9]
+ sb_7__7_/chany_top_in[0] sb_7__7_/chany_top_in[10] sb_7__7_/chany_top_in[11] sb_7__7_/chany_top_in[12]
+ sb_7__7_/chany_top_in[13] sb_7__7_/chany_top_in[14] sb_7__7_/chany_top_in[15] sb_7__7_/chany_top_in[16]
+ sb_7__7_/chany_top_in[17] sb_7__7_/chany_top_in[18] sb_7__7_/chany_top_in[19] sb_7__7_/chany_top_in[1]
+ sb_7__7_/chany_top_in[2] sb_7__7_/chany_top_in[3] sb_7__7_/chany_top_in[4] sb_7__7_/chany_top_in[5]
+ sb_7__7_/chany_top_in[6] sb_7__7_/chany_top_in[7] sb_7__7_/chany_top_in[8] sb_7__7_/chany_top_in[9]
+ sb_7__7_/chany_top_out[0] sb_7__7_/chany_top_out[10] sb_7__7_/chany_top_out[11]
+ sb_7__7_/chany_top_out[12] sb_7__7_/chany_top_out[13] sb_7__7_/chany_top_out[14]
+ sb_7__7_/chany_top_out[15] sb_7__7_/chany_top_out[16] sb_7__7_/chany_top_out[17]
+ sb_7__7_/chany_top_out[18] sb_7__7_/chany_top_out[19] sb_7__7_/chany_top_out[1]
+ sb_7__7_/chany_top_out[2] sb_7__7_/chany_top_out[3] sb_7__7_/chany_top_out[4] sb_7__7_/chany_top_out[5]
+ sb_7__7_/chany_top_out[6] sb_7__7_/chany_top_out[7] sb_7__7_/chany_top_out[8] sb_7__7_/chany_top_out[9]
+ sb_7__7_/clk_1_E_out sb_7__7_/clk_1_N_in sb_7__7_/clk_1_W_out sb_7__7_/clk_2_E_out
+ sb_7__7_/clk_2_N_in sb_7__7_/clk_2_N_out sb_7__7_/clk_2_S_out sb_7__7_/clk_2_W_out
+ sb_7__7_/clk_3_E_out sb_7__7_/clk_3_N_in sb_7__7_/clk_3_N_out sb_7__7_/clk_3_S_out
+ sb_7__7_/clk_3_W_out sb_7__7_/left_bottom_grid_pin_34_ sb_7__7_/left_bottom_grid_pin_35_
+ sb_7__7_/left_bottom_grid_pin_36_ sb_7__7_/left_bottom_grid_pin_37_ sb_7__7_/left_bottom_grid_pin_38_
+ sb_7__7_/left_bottom_grid_pin_39_ sb_7__7_/left_bottom_grid_pin_40_ sb_7__7_/left_bottom_grid_pin_41_
+ sb_7__7_/prog_clk_0_N_in sb_7__7_/prog_clk_1_E_out sb_7__7_/prog_clk_1_N_in sb_7__7_/prog_clk_1_W_out
+ sb_7__7_/prog_clk_2_E_out sb_7__7_/prog_clk_2_N_in sb_7__7_/prog_clk_2_N_out sb_7__7_/prog_clk_2_S_out
+ sb_7__7_/prog_clk_2_W_out sb_7__7_/prog_clk_3_E_out sb_7__7_/prog_clk_3_N_in sb_7__7_/prog_clk_3_N_out
+ sb_7__7_/prog_clk_3_S_out sb_7__7_/prog_clk_3_W_out sb_7__7_/right_bottom_grid_pin_34_
+ sb_7__7_/right_bottom_grid_pin_35_ sb_7__7_/right_bottom_grid_pin_36_ sb_7__7_/right_bottom_grid_pin_37_
+ sb_7__7_/right_bottom_grid_pin_38_ sb_7__7_/right_bottom_grid_pin_39_ sb_7__7_/right_bottom_grid_pin_40_
+ sb_7__7_/right_bottom_grid_pin_41_ sb_7__7_/top_left_grid_pin_42_ sb_7__7_/top_left_grid_pin_43_
+ sb_7__7_/top_left_grid_pin_44_ sb_7__7_/top_left_grid_pin_45_ sb_7__7_/top_left_grid_pin_46_
+ sb_7__7_/top_left_grid_pin_47_ sb_7__7_/top_left_grid_pin_48_ sb_7__7_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_4__4_ sb_4__4_/Test_en_N_out sb_4__4_/Test_en_S_in VGND VPWR sb_4__4_/bottom_left_grid_pin_42_
+ sb_4__4_/bottom_left_grid_pin_43_ sb_4__4_/bottom_left_grid_pin_44_ sb_4__4_/bottom_left_grid_pin_45_
+ sb_4__4_/bottom_left_grid_pin_46_ sb_4__4_/bottom_left_grid_pin_47_ sb_4__4_/bottom_left_grid_pin_48_
+ sb_4__4_/bottom_left_grid_pin_49_ sb_4__4_/ccff_head sb_4__4_/ccff_tail sb_4__4_/chanx_left_in[0]
+ sb_4__4_/chanx_left_in[10] sb_4__4_/chanx_left_in[11] sb_4__4_/chanx_left_in[12]
+ sb_4__4_/chanx_left_in[13] sb_4__4_/chanx_left_in[14] sb_4__4_/chanx_left_in[15]
+ sb_4__4_/chanx_left_in[16] sb_4__4_/chanx_left_in[17] sb_4__4_/chanx_left_in[18]
+ sb_4__4_/chanx_left_in[19] sb_4__4_/chanx_left_in[1] sb_4__4_/chanx_left_in[2] sb_4__4_/chanx_left_in[3]
+ sb_4__4_/chanx_left_in[4] sb_4__4_/chanx_left_in[5] sb_4__4_/chanx_left_in[6] sb_4__4_/chanx_left_in[7]
+ sb_4__4_/chanx_left_in[8] sb_4__4_/chanx_left_in[9] sb_4__4_/chanx_left_out[0] sb_4__4_/chanx_left_out[10]
+ sb_4__4_/chanx_left_out[11] sb_4__4_/chanx_left_out[12] sb_4__4_/chanx_left_out[13]
+ sb_4__4_/chanx_left_out[14] sb_4__4_/chanx_left_out[15] sb_4__4_/chanx_left_out[16]
+ sb_4__4_/chanx_left_out[17] sb_4__4_/chanx_left_out[18] sb_4__4_/chanx_left_out[19]
+ sb_4__4_/chanx_left_out[1] sb_4__4_/chanx_left_out[2] sb_4__4_/chanx_left_out[3]
+ sb_4__4_/chanx_left_out[4] sb_4__4_/chanx_left_out[5] sb_4__4_/chanx_left_out[6]
+ sb_4__4_/chanx_left_out[7] sb_4__4_/chanx_left_out[8] sb_4__4_/chanx_left_out[9]
+ sb_4__4_/chanx_right_in[0] sb_4__4_/chanx_right_in[10] sb_4__4_/chanx_right_in[11]
+ sb_4__4_/chanx_right_in[12] sb_4__4_/chanx_right_in[13] sb_4__4_/chanx_right_in[14]
+ sb_4__4_/chanx_right_in[15] sb_4__4_/chanx_right_in[16] sb_4__4_/chanx_right_in[17]
+ sb_4__4_/chanx_right_in[18] sb_4__4_/chanx_right_in[19] sb_4__4_/chanx_right_in[1]
+ sb_4__4_/chanx_right_in[2] sb_4__4_/chanx_right_in[3] sb_4__4_/chanx_right_in[4]
+ sb_4__4_/chanx_right_in[5] sb_4__4_/chanx_right_in[6] sb_4__4_/chanx_right_in[7]
+ sb_4__4_/chanx_right_in[8] sb_4__4_/chanx_right_in[9] cbx_5__4_/chanx_left_in[0]
+ cbx_5__4_/chanx_left_in[10] cbx_5__4_/chanx_left_in[11] cbx_5__4_/chanx_left_in[12]
+ cbx_5__4_/chanx_left_in[13] cbx_5__4_/chanx_left_in[14] cbx_5__4_/chanx_left_in[15]
+ cbx_5__4_/chanx_left_in[16] cbx_5__4_/chanx_left_in[17] cbx_5__4_/chanx_left_in[18]
+ cbx_5__4_/chanx_left_in[19] cbx_5__4_/chanx_left_in[1] cbx_5__4_/chanx_left_in[2]
+ cbx_5__4_/chanx_left_in[3] cbx_5__4_/chanx_left_in[4] cbx_5__4_/chanx_left_in[5]
+ cbx_5__4_/chanx_left_in[6] cbx_5__4_/chanx_left_in[7] cbx_5__4_/chanx_left_in[8]
+ cbx_5__4_/chanx_left_in[9] cby_4__4_/chany_top_out[0] cby_4__4_/chany_top_out[10]
+ cby_4__4_/chany_top_out[11] cby_4__4_/chany_top_out[12] cby_4__4_/chany_top_out[13]
+ cby_4__4_/chany_top_out[14] cby_4__4_/chany_top_out[15] cby_4__4_/chany_top_out[16]
+ cby_4__4_/chany_top_out[17] cby_4__4_/chany_top_out[18] cby_4__4_/chany_top_out[19]
+ cby_4__4_/chany_top_out[1] cby_4__4_/chany_top_out[2] cby_4__4_/chany_top_out[3]
+ cby_4__4_/chany_top_out[4] cby_4__4_/chany_top_out[5] cby_4__4_/chany_top_out[6]
+ cby_4__4_/chany_top_out[7] cby_4__4_/chany_top_out[8] cby_4__4_/chany_top_out[9]
+ cby_4__4_/chany_top_in[0] cby_4__4_/chany_top_in[10] cby_4__4_/chany_top_in[11]
+ cby_4__4_/chany_top_in[12] cby_4__4_/chany_top_in[13] cby_4__4_/chany_top_in[14]
+ cby_4__4_/chany_top_in[15] cby_4__4_/chany_top_in[16] cby_4__4_/chany_top_in[17]
+ cby_4__4_/chany_top_in[18] cby_4__4_/chany_top_in[19] cby_4__4_/chany_top_in[1]
+ cby_4__4_/chany_top_in[2] cby_4__4_/chany_top_in[3] cby_4__4_/chany_top_in[4] cby_4__4_/chany_top_in[5]
+ cby_4__4_/chany_top_in[6] cby_4__4_/chany_top_in[7] cby_4__4_/chany_top_in[8] cby_4__4_/chany_top_in[9]
+ sb_4__4_/chany_top_in[0] sb_4__4_/chany_top_in[10] sb_4__4_/chany_top_in[11] sb_4__4_/chany_top_in[12]
+ sb_4__4_/chany_top_in[13] sb_4__4_/chany_top_in[14] sb_4__4_/chany_top_in[15] sb_4__4_/chany_top_in[16]
+ sb_4__4_/chany_top_in[17] sb_4__4_/chany_top_in[18] sb_4__4_/chany_top_in[19] sb_4__4_/chany_top_in[1]
+ sb_4__4_/chany_top_in[2] sb_4__4_/chany_top_in[3] sb_4__4_/chany_top_in[4] sb_4__4_/chany_top_in[5]
+ sb_4__4_/chany_top_in[6] sb_4__4_/chany_top_in[7] sb_4__4_/chany_top_in[8] sb_4__4_/chany_top_in[9]
+ sb_4__4_/chany_top_out[0] sb_4__4_/chany_top_out[10] sb_4__4_/chany_top_out[11]
+ sb_4__4_/chany_top_out[12] sb_4__4_/chany_top_out[13] sb_4__4_/chany_top_out[14]
+ sb_4__4_/chany_top_out[15] sb_4__4_/chany_top_out[16] sb_4__4_/chany_top_out[17]
+ sb_4__4_/chany_top_out[18] sb_4__4_/chany_top_out[19] sb_4__4_/chany_top_out[1]
+ sb_4__4_/chany_top_out[2] sb_4__4_/chany_top_out[3] sb_4__4_/chany_top_out[4] sb_4__4_/chany_top_out[5]
+ sb_4__4_/chany_top_out[6] sb_4__4_/chany_top_out[7] sb_4__4_/chany_top_out[8] sb_4__4_/chany_top_out[9]
+ sb_4__4_/clk_1_E_out sb_4__4_/clk_1_N_in sb_4__4_/clk_1_W_out sb_4__4_/clk_2_E_out
+ sb_4__4_/clk_2_N_in sb_4__4_/clk_2_N_out sb_4__4_/clk_2_S_out sb_4__4_/clk_2_W_out
+ sb_4__4_/clk_3_E_out sb_4__4_/clk_3_N_in sb_4__4_/clk_3_N_out sb_4__4_/clk_3_S_out
+ sb_4__4_/clk_3_W_out sb_4__4_/left_bottom_grid_pin_34_ sb_4__4_/left_bottom_grid_pin_35_
+ sb_4__4_/left_bottom_grid_pin_36_ sb_4__4_/left_bottom_grid_pin_37_ sb_4__4_/left_bottom_grid_pin_38_
+ sb_4__4_/left_bottom_grid_pin_39_ sb_4__4_/left_bottom_grid_pin_40_ sb_4__4_/left_bottom_grid_pin_41_
+ sb_4__4_/prog_clk_0_N_in sb_4__4_/prog_clk_1_E_out sb_4__4_/prog_clk_1_N_in sb_4__4_/prog_clk_1_W_out
+ sb_4__4_/prog_clk_2_E_out sb_4__4_/prog_clk_2_N_in sb_4__4_/prog_clk_2_N_out sb_4__4_/prog_clk_2_S_out
+ sb_4__4_/prog_clk_2_W_out sb_4__4_/prog_clk_3_E_out sb_4__4_/prog_clk_3_N_in sb_4__4_/prog_clk_3_N_out
+ sb_4__4_/prog_clk_3_S_out sb_4__4_/prog_clk_3_W_out sb_4__4_/right_bottom_grid_pin_34_
+ sb_4__4_/right_bottom_grid_pin_35_ sb_4__4_/right_bottom_grid_pin_36_ sb_4__4_/right_bottom_grid_pin_37_
+ sb_4__4_/right_bottom_grid_pin_38_ sb_4__4_/right_bottom_grid_pin_39_ sb_4__4_/right_bottom_grid_pin_40_
+ sb_4__4_/right_bottom_grid_pin_41_ sb_4__4_/top_left_grid_pin_42_ sb_4__4_/top_left_grid_pin_43_
+ sb_4__4_/top_left_grid_pin_44_ sb_4__4_/top_left_grid_pin_45_ sb_4__4_/top_left_grid_pin_46_
+ sb_4__4_/top_left_grid_pin_47_ sb_4__4_/top_left_grid_pin_48_ sb_4__4_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_1__1_ sb_1__1_/Test_en_N_out sb_1__1_/Test_en_S_in VGND VPWR sb_1__1_/bottom_left_grid_pin_42_
+ sb_1__1_/bottom_left_grid_pin_43_ sb_1__1_/bottom_left_grid_pin_44_ sb_1__1_/bottom_left_grid_pin_45_
+ sb_1__1_/bottom_left_grid_pin_46_ sb_1__1_/bottom_left_grid_pin_47_ sb_1__1_/bottom_left_grid_pin_48_
+ sb_1__1_/bottom_left_grid_pin_49_ sb_1__1_/ccff_head sb_1__1_/ccff_tail sb_1__1_/chanx_left_in[0]
+ sb_1__1_/chanx_left_in[10] sb_1__1_/chanx_left_in[11] sb_1__1_/chanx_left_in[12]
+ sb_1__1_/chanx_left_in[13] sb_1__1_/chanx_left_in[14] sb_1__1_/chanx_left_in[15]
+ sb_1__1_/chanx_left_in[16] sb_1__1_/chanx_left_in[17] sb_1__1_/chanx_left_in[18]
+ sb_1__1_/chanx_left_in[19] sb_1__1_/chanx_left_in[1] sb_1__1_/chanx_left_in[2] sb_1__1_/chanx_left_in[3]
+ sb_1__1_/chanx_left_in[4] sb_1__1_/chanx_left_in[5] sb_1__1_/chanx_left_in[6] sb_1__1_/chanx_left_in[7]
+ sb_1__1_/chanx_left_in[8] sb_1__1_/chanx_left_in[9] sb_1__1_/chanx_left_out[0] sb_1__1_/chanx_left_out[10]
+ sb_1__1_/chanx_left_out[11] sb_1__1_/chanx_left_out[12] sb_1__1_/chanx_left_out[13]
+ sb_1__1_/chanx_left_out[14] sb_1__1_/chanx_left_out[15] sb_1__1_/chanx_left_out[16]
+ sb_1__1_/chanx_left_out[17] sb_1__1_/chanx_left_out[18] sb_1__1_/chanx_left_out[19]
+ sb_1__1_/chanx_left_out[1] sb_1__1_/chanx_left_out[2] sb_1__1_/chanx_left_out[3]
+ sb_1__1_/chanx_left_out[4] sb_1__1_/chanx_left_out[5] sb_1__1_/chanx_left_out[6]
+ sb_1__1_/chanx_left_out[7] sb_1__1_/chanx_left_out[8] sb_1__1_/chanx_left_out[9]
+ sb_1__1_/chanx_right_in[0] sb_1__1_/chanx_right_in[10] sb_1__1_/chanx_right_in[11]
+ sb_1__1_/chanx_right_in[12] sb_1__1_/chanx_right_in[13] sb_1__1_/chanx_right_in[14]
+ sb_1__1_/chanx_right_in[15] sb_1__1_/chanx_right_in[16] sb_1__1_/chanx_right_in[17]
+ sb_1__1_/chanx_right_in[18] sb_1__1_/chanx_right_in[19] sb_1__1_/chanx_right_in[1]
+ sb_1__1_/chanx_right_in[2] sb_1__1_/chanx_right_in[3] sb_1__1_/chanx_right_in[4]
+ sb_1__1_/chanx_right_in[5] sb_1__1_/chanx_right_in[6] sb_1__1_/chanx_right_in[7]
+ sb_1__1_/chanx_right_in[8] sb_1__1_/chanx_right_in[9] cbx_2__1_/chanx_left_in[0]
+ cbx_2__1_/chanx_left_in[10] cbx_2__1_/chanx_left_in[11] cbx_2__1_/chanx_left_in[12]
+ cbx_2__1_/chanx_left_in[13] cbx_2__1_/chanx_left_in[14] cbx_2__1_/chanx_left_in[15]
+ cbx_2__1_/chanx_left_in[16] cbx_2__1_/chanx_left_in[17] cbx_2__1_/chanx_left_in[18]
+ cbx_2__1_/chanx_left_in[19] cbx_2__1_/chanx_left_in[1] cbx_2__1_/chanx_left_in[2]
+ cbx_2__1_/chanx_left_in[3] cbx_2__1_/chanx_left_in[4] cbx_2__1_/chanx_left_in[5]
+ cbx_2__1_/chanx_left_in[6] cbx_2__1_/chanx_left_in[7] cbx_2__1_/chanx_left_in[8]
+ cbx_2__1_/chanx_left_in[9] cby_1__1_/chany_top_out[0] cby_1__1_/chany_top_out[10]
+ cby_1__1_/chany_top_out[11] cby_1__1_/chany_top_out[12] cby_1__1_/chany_top_out[13]
+ cby_1__1_/chany_top_out[14] cby_1__1_/chany_top_out[15] cby_1__1_/chany_top_out[16]
+ cby_1__1_/chany_top_out[17] cby_1__1_/chany_top_out[18] cby_1__1_/chany_top_out[19]
+ cby_1__1_/chany_top_out[1] cby_1__1_/chany_top_out[2] cby_1__1_/chany_top_out[3]
+ cby_1__1_/chany_top_out[4] cby_1__1_/chany_top_out[5] cby_1__1_/chany_top_out[6]
+ cby_1__1_/chany_top_out[7] cby_1__1_/chany_top_out[8] cby_1__1_/chany_top_out[9]
+ cby_1__1_/chany_top_in[0] cby_1__1_/chany_top_in[10] cby_1__1_/chany_top_in[11]
+ cby_1__1_/chany_top_in[12] cby_1__1_/chany_top_in[13] cby_1__1_/chany_top_in[14]
+ cby_1__1_/chany_top_in[15] cby_1__1_/chany_top_in[16] cby_1__1_/chany_top_in[17]
+ cby_1__1_/chany_top_in[18] cby_1__1_/chany_top_in[19] cby_1__1_/chany_top_in[1]
+ cby_1__1_/chany_top_in[2] cby_1__1_/chany_top_in[3] cby_1__1_/chany_top_in[4] cby_1__1_/chany_top_in[5]
+ cby_1__1_/chany_top_in[6] cby_1__1_/chany_top_in[7] cby_1__1_/chany_top_in[8] cby_1__1_/chany_top_in[9]
+ sb_1__1_/chany_top_in[0] sb_1__1_/chany_top_in[10] sb_1__1_/chany_top_in[11] sb_1__1_/chany_top_in[12]
+ sb_1__1_/chany_top_in[13] sb_1__1_/chany_top_in[14] sb_1__1_/chany_top_in[15] sb_1__1_/chany_top_in[16]
+ sb_1__1_/chany_top_in[17] sb_1__1_/chany_top_in[18] sb_1__1_/chany_top_in[19] sb_1__1_/chany_top_in[1]
+ sb_1__1_/chany_top_in[2] sb_1__1_/chany_top_in[3] sb_1__1_/chany_top_in[4] sb_1__1_/chany_top_in[5]
+ sb_1__1_/chany_top_in[6] sb_1__1_/chany_top_in[7] sb_1__1_/chany_top_in[8] sb_1__1_/chany_top_in[9]
+ sb_1__1_/chany_top_out[0] sb_1__1_/chany_top_out[10] sb_1__1_/chany_top_out[11]
+ sb_1__1_/chany_top_out[12] sb_1__1_/chany_top_out[13] sb_1__1_/chany_top_out[14]
+ sb_1__1_/chany_top_out[15] sb_1__1_/chany_top_out[16] sb_1__1_/chany_top_out[17]
+ sb_1__1_/chany_top_out[18] sb_1__1_/chany_top_out[19] sb_1__1_/chany_top_out[1]
+ sb_1__1_/chany_top_out[2] sb_1__1_/chany_top_out[3] sb_1__1_/chany_top_out[4] sb_1__1_/chany_top_out[5]
+ sb_1__1_/chany_top_out[6] sb_1__1_/chany_top_out[7] sb_1__1_/chany_top_out[8] sb_1__1_/chany_top_out[9]
+ sb_1__1_/clk_1_E_out sb_1__1_/clk_1_N_in sb_1__1_/clk_1_W_out sb_1__1_/clk_2_E_out
+ sb_1__1_/clk_2_N_in sb_1__1_/clk_2_N_out sb_1__1_/clk_2_S_out sb_1__1_/clk_2_W_out
+ sb_1__1_/clk_3_E_out sb_1__1_/clk_3_N_in sb_1__1_/clk_3_N_out sb_1__1_/clk_3_S_out
+ sb_1__1_/clk_3_W_out sb_1__1_/left_bottom_grid_pin_34_ sb_1__1_/left_bottom_grid_pin_35_
+ sb_1__1_/left_bottom_grid_pin_36_ sb_1__1_/left_bottom_grid_pin_37_ sb_1__1_/left_bottom_grid_pin_38_
+ sb_1__1_/left_bottom_grid_pin_39_ sb_1__1_/left_bottom_grid_pin_40_ sb_1__1_/left_bottom_grid_pin_41_
+ sb_1__1_/prog_clk_0_N_in sb_1__1_/prog_clk_1_E_out sb_1__1_/prog_clk_1_N_in sb_1__1_/prog_clk_1_W_out
+ sb_1__1_/prog_clk_2_E_out sb_1__1_/prog_clk_2_N_in sb_1__1_/prog_clk_2_N_out sb_1__1_/prog_clk_2_S_out
+ sb_1__1_/prog_clk_2_W_out sb_1__1_/prog_clk_3_E_out sb_1__1_/prog_clk_3_N_in sb_1__1_/prog_clk_3_N_out
+ sb_1__1_/prog_clk_3_S_out sb_1__1_/prog_clk_3_W_out sb_1__1_/right_bottom_grid_pin_34_
+ sb_1__1_/right_bottom_grid_pin_35_ sb_1__1_/right_bottom_grid_pin_36_ sb_1__1_/right_bottom_grid_pin_37_
+ sb_1__1_/right_bottom_grid_pin_38_ sb_1__1_/right_bottom_grid_pin_39_ sb_1__1_/right_bottom_grid_pin_40_
+ sb_1__1_/right_bottom_grid_pin_41_ sb_1__1_/top_left_grid_pin_42_ sb_1__1_/top_left_grid_pin_43_
+ sb_1__1_/top_left_grid_pin_44_ sb_1__1_/top_left_grid_pin_45_ sb_1__1_/top_left_grid_pin_46_
+ sb_1__1_/top_left_grid_pin_47_ sb_1__1_/top_left_grid_pin_48_ sb_1__1_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_3__8_ cby_3__8_/Test_en_W_in cby_3__8_/Test_en_E_out cby_3__8_/Test_en_N_out
+ cby_3__8_/Test_en_W_in cby_3__8_/Test_en_W_in cby_3__8_/Test_en_W_out VGND VPWR
+ cby_3__8_/ccff_head cby_3__8_/ccff_tail sb_3__7_/chany_top_out[0] sb_3__7_/chany_top_out[10]
+ sb_3__7_/chany_top_out[11] sb_3__7_/chany_top_out[12] sb_3__7_/chany_top_out[13]
+ sb_3__7_/chany_top_out[14] sb_3__7_/chany_top_out[15] sb_3__7_/chany_top_out[16]
+ sb_3__7_/chany_top_out[17] sb_3__7_/chany_top_out[18] sb_3__7_/chany_top_out[19]
+ sb_3__7_/chany_top_out[1] sb_3__7_/chany_top_out[2] sb_3__7_/chany_top_out[3] sb_3__7_/chany_top_out[4]
+ sb_3__7_/chany_top_out[5] sb_3__7_/chany_top_out[6] sb_3__7_/chany_top_out[7] sb_3__7_/chany_top_out[8]
+ sb_3__7_/chany_top_out[9] sb_3__7_/chany_top_in[0] sb_3__7_/chany_top_in[10] sb_3__7_/chany_top_in[11]
+ sb_3__7_/chany_top_in[12] sb_3__7_/chany_top_in[13] sb_3__7_/chany_top_in[14] sb_3__7_/chany_top_in[15]
+ sb_3__7_/chany_top_in[16] sb_3__7_/chany_top_in[17] sb_3__7_/chany_top_in[18] sb_3__7_/chany_top_in[19]
+ sb_3__7_/chany_top_in[1] sb_3__7_/chany_top_in[2] sb_3__7_/chany_top_in[3] sb_3__7_/chany_top_in[4]
+ sb_3__7_/chany_top_in[5] sb_3__7_/chany_top_in[6] sb_3__7_/chany_top_in[7] sb_3__7_/chany_top_in[8]
+ sb_3__7_/chany_top_in[9] cby_3__8_/chany_top_in[0] cby_3__8_/chany_top_in[10] cby_3__8_/chany_top_in[11]
+ cby_3__8_/chany_top_in[12] cby_3__8_/chany_top_in[13] cby_3__8_/chany_top_in[14]
+ cby_3__8_/chany_top_in[15] cby_3__8_/chany_top_in[16] cby_3__8_/chany_top_in[17]
+ cby_3__8_/chany_top_in[18] cby_3__8_/chany_top_in[19] cby_3__8_/chany_top_in[1]
+ cby_3__8_/chany_top_in[2] cby_3__8_/chany_top_in[3] cby_3__8_/chany_top_in[4] cby_3__8_/chany_top_in[5]
+ cby_3__8_/chany_top_in[6] cby_3__8_/chany_top_in[7] cby_3__8_/chany_top_in[8] cby_3__8_/chany_top_in[9]
+ cby_3__8_/chany_top_out[0] cby_3__8_/chany_top_out[10] cby_3__8_/chany_top_out[11]
+ cby_3__8_/chany_top_out[12] cby_3__8_/chany_top_out[13] cby_3__8_/chany_top_out[14]
+ cby_3__8_/chany_top_out[15] cby_3__8_/chany_top_out[16] cby_3__8_/chany_top_out[17]
+ cby_3__8_/chany_top_out[18] cby_3__8_/chany_top_out[19] cby_3__8_/chany_top_out[1]
+ cby_3__8_/chany_top_out[2] cby_3__8_/chany_top_out[3] cby_3__8_/chany_top_out[4]
+ cby_3__8_/chany_top_out[5] cby_3__8_/chany_top_out[6] cby_3__8_/chany_top_out[7]
+ cby_3__8_/chany_top_out[8] cby_3__8_/chany_top_out[9] cby_3__8_/clk_2_N_out cby_3__8_/clk_2_S_in
+ cby_3__8_/clk_2_S_out cby_3__8_/clk_3_N_out cby_3__8_/clk_3_S_in cby_3__8_/clk_3_S_out
+ cby_3__8_/left_grid_pin_16_ cby_3__8_/left_grid_pin_17_ cby_3__8_/left_grid_pin_18_
+ cby_3__8_/left_grid_pin_19_ cby_3__8_/left_grid_pin_20_ cby_3__8_/left_grid_pin_21_
+ cby_3__8_/left_grid_pin_22_ cby_3__8_/left_grid_pin_23_ cby_3__8_/left_grid_pin_24_
+ cby_3__8_/left_grid_pin_25_ cby_3__8_/left_grid_pin_26_ cby_3__8_/left_grid_pin_27_
+ cby_3__8_/left_grid_pin_28_ cby_3__8_/left_grid_pin_29_ cby_3__8_/left_grid_pin_30_
+ cby_3__8_/left_grid_pin_31_ sb_3__8_/prog_clk_0_S_in sb_3__7_/prog_clk_0_N_in cby_3__8_/prog_clk_0_W_in
+ cby_3__8_/prog_clk_2_N_out cby_3__8_/prog_clk_2_S_in cby_3__8_/prog_clk_2_S_out
+ cby_3__8_/prog_clk_3_N_out cby_3__8_/prog_clk_3_S_in cby_3__8_/prog_clk_3_S_out
+ cby_1__1_
Xcby_0__5_ IO_ISOL_N VGND VPWR sb_0__5_/ccff_tail cby_0__5_/ccff_tail sb_0__4_/chany_top_out[0]
+ sb_0__4_/chany_top_out[10] sb_0__4_/chany_top_out[11] sb_0__4_/chany_top_out[12]
+ sb_0__4_/chany_top_out[13] sb_0__4_/chany_top_out[14] sb_0__4_/chany_top_out[15]
+ sb_0__4_/chany_top_out[16] sb_0__4_/chany_top_out[17] sb_0__4_/chany_top_out[18]
+ sb_0__4_/chany_top_out[19] sb_0__4_/chany_top_out[1] sb_0__4_/chany_top_out[2] sb_0__4_/chany_top_out[3]
+ sb_0__4_/chany_top_out[4] sb_0__4_/chany_top_out[5] sb_0__4_/chany_top_out[6] sb_0__4_/chany_top_out[7]
+ sb_0__4_/chany_top_out[8] sb_0__4_/chany_top_out[9] sb_0__4_/chany_top_in[0] sb_0__4_/chany_top_in[10]
+ sb_0__4_/chany_top_in[11] sb_0__4_/chany_top_in[12] sb_0__4_/chany_top_in[13] sb_0__4_/chany_top_in[14]
+ sb_0__4_/chany_top_in[15] sb_0__4_/chany_top_in[16] sb_0__4_/chany_top_in[17] sb_0__4_/chany_top_in[18]
+ sb_0__4_/chany_top_in[19] sb_0__4_/chany_top_in[1] sb_0__4_/chany_top_in[2] sb_0__4_/chany_top_in[3]
+ sb_0__4_/chany_top_in[4] sb_0__4_/chany_top_in[5] sb_0__4_/chany_top_in[6] sb_0__4_/chany_top_in[7]
+ sb_0__4_/chany_top_in[8] sb_0__4_/chany_top_in[9] cby_0__5_/chany_top_in[0] cby_0__5_/chany_top_in[10]
+ cby_0__5_/chany_top_in[11] cby_0__5_/chany_top_in[12] cby_0__5_/chany_top_in[13]
+ cby_0__5_/chany_top_in[14] cby_0__5_/chany_top_in[15] cby_0__5_/chany_top_in[16]
+ cby_0__5_/chany_top_in[17] cby_0__5_/chany_top_in[18] cby_0__5_/chany_top_in[19]
+ cby_0__5_/chany_top_in[1] cby_0__5_/chany_top_in[2] cby_0__5_/chany_top_in[3] cby_0__5_/chany_top_in[4]
+ cby_0__5_/chany_top_in[5] cby_0__5_/chany_top_in[6] cby_0__5_/chany_top_in[7] cby_0__5_/chany_top_in[8]
+ cby_0__5_/chany_top_in[9] cby_0__5_/chany_top_out[0] cby_0__5_/chany_top_out[10]
+ cby_0__5_/chany_top_out[11] cby_0__5_/chany_top_out[12] cby_0__5_/chany_top_out[13]
+ cby_0__5_/chany_top_out[14] cby_0__5_/chany_top_out[15] cby_0__5_/chany_top_out[16]
+ cby_0__5_/chany_top_out[17] cby_0__5_/chany_top_out[18] cby_0__5_/chany_top_out[19]
+ cby_0__5_/chany_top_out[1] cby_0__5_/chany_top_out[2] cby_0__5_/chany_top_out[3]
+ cby_0__5_/chany_top_out[4] cby_0__5_/chany_top_out[5] cby_0__5_/chany_top_out[6]
+ cby_0__5_/chany_top_out[7] cby_0__5_/chany_top_out[8] cby_0__5_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
+ cby_0__5_/left_grid_pin_0_ cby_0__5_/prog_clk_0_E_in cby_0__5_/left_grid_pin_0_
+ sb_0__4_/top_left_grid_pin_1_ sb_0__5_/bottom_left_grid_pin_1_ cby_0__1_
Xcbx_7__1_ cbx_7__1_/REGIN_FEEDTHROUGH cbx_7__1_/REGOUT_FEEDTHROUGH cbx_7__1_/SC_IN_BOT
+ cbx_7__1_/SC_IN_TOP cbx_7__1_/SC_OUT_BOT cbx_7__1_/SC_OUT_TOP VGND VPWR cbx_7__1_/bottom_grid_pin_0_
+ cbx_7__1_/bottom_grid_pin_10_ cbx_7__1_/bottom_grid_pin_11_ cbx_7__1_/bottom_grid_pin_12_
+ cbx_7__1_/bottom_grid_pin_13_ cbx_7__1_/bottom_grid_pin_14_ cbx_7__1_/bottom_grid_pin_15_
+ cbx_7__1_/bottom_grid_pin_1_ cbx_7__1_/bottom_grid_pin_2_ cbx_7__1_/bottom_grid_pin_3_
+ cbx_7__1_/bottom_grid_pin_4_ cbx_7__1_/bottom_grid_pin_5_ cbx_7__1_/bottom_grid_pin_6_
+ cbx_7__1_/bottom_grid_pin_7_ cbx_7__1_/bottom_grid_pin_8_ cbx_7__1_/bottom_grid_pin_9_
+ sb_7__1_/ccff_tail sb_6__1_/ccff_head cbx_7__1_/chanx_left_in[0] cbx_7__1_/chanx_left_in[10]
+ cbx_7__1_/chanx_left_in[11] cbx_7__1_/chanx_left_in[12] cbx_7__1_/chanx_left_in[13]
+ cbx_7__1_/chanx_left_in[14] cbx_7__1_/chanx_left_in[15] cbx_7__1_/chanx_left_in[16]
+ cbx_7__1_/chanx_left_in[17] cbx_7__1_/chanx_left_in[18] cbx_7__1_/chanx_left_in[19]
+ cbx_7__1_/chanx_left_in[1] cbx_7__1_/chanx_left_in[2] cbx_7__1_/chanx_left_in[3]
+ cbx_7__1_/chanx_left_in[4] cbx_7__1_/chanx_left_in[5] cbx_7__1_/chanx_left_in[6]
+ cbx_7__1_/chanx_left_in[7] cbx_7__1_/chanx_left_in[8] cbx_7__1_/chanx_left_in[9]
+ sb_6__1_/chanx_right_in[0] sb_6__1_/chanx_right_in[10] sb_6__1_/chanx_right_in[11]
+ sb_6__1_/chanx_right_in[12] sb_6__1_/chanx_right_in[13] sb_6__1_/chanx_right_in[14]
+ sb_6__1_/chanx_right_in[15] sb_6__1_/chanx_right_in[16] sb_6__1_/chanx_right_in[17]
+ sb_6__1_/chanx_right_in[18] sb_6__1_/chanx_right_in[19] sb_6__1_/chanx_right_in[1]
+ sb_6__1_/chanx_right_in[2] sb_6__1_/chanx_right_in[3] sb_6__1_/chanx_right_in[4]
+ sb_6__1_/chanx_right_in[5] sb_6__1_/chanx_right_in[6] sb_6__1_/chanx_right_in[7]
+ sb_6__1_/chanx_right_in[8] sb_6__1_/chanx_right_in[9] sb_7__1_/chanx_left_out[0]
+ sb_7__1_/chanx_left_out[10] sb_7__1_/chanx_left_out[11] sb_7__1_/chanx_left_out[12]
+ sb_7__1_/chanx_left_out[13] sb_7__1_/chanx_left_out[14] sb_7__1_/chanx_left_out[15]
+ sb_7__1_/chanx_left_out[16] sb_7__1_/chanx_left_out[17] sb_7__1_/chanx_left_out[18]
+ sb_7__1_/chanx_left_out[19] sb_7__1_/chanx_left_out[1] sb_7__1_/chanx_left_out[2]
+ sb_7__1_/chanx_left_out[3] sb_7__1_/chanx_left_out[4] sb_7__1_/chanx_left_out[5]
+ sb_7__1_/chanx_left_out[6] sb_7__1_/chanx_left_out[7] sb_7__1_/chanx_left_out[8]
+ sb_7__1_/chanx_left_out[9] sb_7__1_/chanx_left_in[0] sb_7__1_/chanx_left_in[10]
+ sb_7__1_/chanx_left_in[11] sb_7__1_/chanx_left_in[12] sb_7__1_/chanx_left_in[13]
+ sb_7__1_/chanx_left_in[14] sb_7__1_/chanx_left_in[15] sb_7__1_/chanx_left_in[16]
+ sb_7__1_/chanx_left_in[17] sb_7__1_/chanx_left_in[18] sb_7__1_/chanx_left_in[19]
+ sb_7__1_/chanx_left_in[1] sb_7__1_/chanx_left_in[2] sb_7__1_/chanx_left_in[3] sb_7__1_/chanx_left_in[4]
+ sb_7__1_/chanx_left_in[5] sb_7__1_/chanx_left_in[6] sb_7__1_/chanx_left_in[7] sb_7__1_/chanx_left_in[8]
+ sb_7__1_/chanx_left_in[9] cbx_7__1_/clk_1_N_out cbx_7__1_/clk_1_S_out sb_7__1_/clk_1_W_out
+ cbx_7__1_/clk_2_E_out cbx_7__1_/clk_2_W_in cbx_7__1_/clk_2_W_out cbx_7__1_/clk_3_E_out
+ cbx_7__1_/clk_3_W_in cbx_7__1_/clk_3_W_out cbx_7__1_/prog_clk_0_N_in cbx_7__1_/prog_clk_0_W_out
+ cbx_7__1_/prog_clk_1_N_out cbx_7__1_/prog_clk_1_S_out sb_7__1_/prog_clk_1_W_out
+ cbx_7__1_/prog_clk_2_E_out cbx_7__1_/prog_clk_2_W_in cbx_7__1_/prog_clk_2_W_out
+ cbx_7__1_/prog_clk_3_E_out cbx_7__1_/prog_clk_3_W_in cbx_7__1_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_7__6_ sb_7__6_/Test_en_N_out sb_7__6_/Test_en_S_in VGND VPWR sb_7__6_/bottom_left_grid_pin_42_
+ sb_7__6_/bottom_left_grid_pin_43_ sb_7__6_/bottom_left_grid_pin_44_ sb_7__6_/bottom_left_grid_pin_45_
+ sb_7__6_/bottom_left_grid_pin_46_ sb_7__6_/bottom_left_grid_pin_47_ sb_7__6_/bottom_left_grid_pin_48_
+ sb_7__6_/bottom_left_grid_pin_49_ sb_7__6_/ccff_head sb_7__6_/ccff_tail sb_7__6_/chanx_left_in[0]
+ sb_7__6_/chanx_left_in[10] sb_7__6_/chanx_left_in[11] sb_7__6_/chanx_left_in[12]
+ sb_7__6_/chanx_left_in[13] sb_7__6_/chanx_left_in[14] sb_7__6_/chanx_left_in[15]
+ sb_7__6_/chanx_left_in[16] sb_7__6_/chanx_left_in[17] sb_7__6_/chanx_left_in[18]
+ sb_7__6_/chanx_left_in[19] sb_7__6_/chanx_left_in[1] sb_7__6_/chanx_left_in[2] sb_7__6_/chanx_left_in[3]
+ sb_7__6_/chanx_left_in[4] sb_7__6_/chanx_left_in[5] sb_7__6_/chanx_left_in[6] sb_7__6_/chanx_left_in[7]
+ sb_7__6_/chanx_left_in[8] sb_7__6_/chanx_left_in[9] sb_7__6_/chanx_left_out[0] sb_7__6_/chanx_left_out[10]
+ sb_7__6_/chanx_left_out[11] sb_7__6_/chanx_left_out[12] sb_7__6_/chanx_left_out[13]
+ sb_7__6_/chanx_left_out[14] sb_7__6_/chanx_left_out[15] sb_7__6_/chanx_left_out[16]
+ sb_7__6_/chanx_left_out[17] sb_7__6_/chanx_left_out[18] sb_7__6_/chanx_left_out[19]
+ sb_7__6_/chanx_left_out[1] sb_7__6_/chanx_left_out[2] sb_7__6_/chanx_left_out[3]
+ sb_7__6_/chanx_left_out[4] sb_7__6_/chanx_left_out[5] sb_7__6_/chanx_left_out[6]
+ sb_7__6_/chanx_left_out[7] sb_7__6_/chanx_left_out[8] sb_7__6_/chanx_left_out[9]
+ sb_7__6_/chanx_right_in[0] sb_7__6_/chanx_right_in[10] sb_7__6_/chanx_right_in[11]
+ sb_7__6_/chanx_right_in[12] sb_7__6_/chanx_right_in[13] sb_7__6_/chanx_right_in[14]
+ sb_7__6_/chanx_right_in[15] sb_7__6_/chanx_right_in[16] sb_7__6_/chanx_right_in[17]
+ sb_7__6_/chanx_right_in[18] sb_7__6_/chanx_right_in[19] sb_7__6_/chanx_right_in[1]
+ sb_7__6_/chanx_right_in[2] sb_7__6_/chanx_right_in[3] sb_7__6_/chanx_right_in[4]
+ sb_7__6_/chanx_right_in[5] sb_7__6_/chanx_right_in[6] sb_7__6_/chanx_right_in[7]
+ sb_7__6_/chanx_right_in[8] sb_7__6_/chanx_right_in[9] cbx_8__6_/chanx_left_in[0]
+ cbx_8__6_/chanx_left_in[10] cbx_8__6_/chanx_left_in[11] cbx_8__6_/chanx_left_in[12]
+ cbx_8__6_/chanx_left_in[13] cbx_8__6_/chanx_left_in[14] cbx_8__6_/chanx_left_in[15]
+ cbx_8__6_/chanx_left_in[16] cbx_8__6_/chanx_left_in[17] cbx_8__6_/chanx_left_in[18]
+ cbx_8__6_/chanx_left_in[19] cbx_8__6_/chanx_left_in[1] cbx_8__6_/chanx_left_in[2]
+ cbx_8__6_/chanx_left_in[3] cbx_8__6_/chanx_left_in[4] cbx_8__6_/chanx_left_in[5]
+ cbx_8__6_/chanx_left_in[6] cbx_8__6_/chanx_left_in[7] cbx_8__6_/chanx_left_in[8]
+ cbx_8__6_/chanx_left_in[9] cby_7__6_/chany_top_out[0] cby_7__6_/chany_top_out[10]
+ cby_7__6_/chany_top_out[11] cby_7__6_/chany_top_out[12] cby_7__6_/chany_top_out[13]
+ cby_7__6_/chany_top_out[14] cby_7__6_/chany_top_out[15] cby_7__6_/chany_top_out[16]
+ cby_7__6_/chany_top_out[17] cby_7__6_/chany_top_out[18] cby_7__6_/chany_top_out[19]
+ cby_7__6_/chany_top_out[1] cby_7__6_/chany_top_out[2] cby_7__6_/chany_top_out[3]
+ cby_7__6_/chany_top_out[4] cby_7__6_/chany_top_out[5] cby_7__6_/chany_top_out[6]
+ cby_7__6_/chany_top_out[7] cby_7__6_/chany_top_out[8] cby_7__6_/chany_top_out[9]
+ cby_7__6_/chany_top_in[0] cby_7__6_/chany_top_in[10] cby_7__6_/chany_top_in[11]
+ cby_7__6_/chany_top_in[12] cby_7__6_/chany_top_in[13] cby_7__6_/chany_top_in[14]
+ cby_7__6_/chany_top_in[15] cby_7__6_/chany_top_in[16] cby_7__6_/chany_top_in[17]
+ cby_7__6_/chany_top_in[18] cby_7__6_/chany_top_in[19] cby_7__6_/chany_top_in[1]
+ cby_7__6_/chany_top_in[2] cby_7__6_/chany_top_in[3] cby_7__6_/chany_top_in[4] cby_7__6_/chany_top_in[5]
+ cby_7__6_/chany_top_in[6] cby_7__6_/chany_top_in[7] cby_7__6_/chany_top_in[8] cby_7__6_/chany_top_in[9]
+ sb_7__6_/chany_top_in[0] sb_7__6_/chany_top_in[10] sb_7__6_/chany_top_in[11] sb_7__6_/chany_top_in[12]
+ sb_7__6_/chany_top_in[13] sb_7__6_/chany_top_in[14] sb_7__6_/chany_top_in[15] sb_7__6_/chany_top_in[16]
+ sb_7__6_/chany_top_in[17] sb_7__6_/chany_top_in[18] sb_7__6_/chany_top_in[19] sb_7__6_/chany_top_in[1]
+ sb_7__6_/chany_top_in[2] sb_7__6_/chany_top_in[3] sb_7__6_/chany_top_in[4] sb_7__6_/chany_top_in[5]
+ sb_7__6_/chany_top_in[6] sb_7__6_/chany_top_in[7] sb_7__6_/chany_top_in[8] sb_7__6_/chany_top_in[9]
+ sb_7__6_/chany_top_out[0] sb_7__6_/chany_top_out[10] sb_7__6_/chany_top_out[11]
+ sb_7__6_/chany_top_out[12] sb_7__6_/chany_top_out[13] sb_7__6_/chany_top_out[14]
+ sb_7__6_/chany_top_out[15] sb_7__6_/chany_top_out[16] sb_7__6_/chany_top_out[17]
+ sb_7__6_/chany_top_out[18] sb_7__6_/chany_top_out[19] sb_7__6_/chany_top_out[1]
+ sb_7__6_/chany_top_out[2] sb_7__6_/chany_top_out[3] sb_7__6_/chany_top_out[4] sb_7__6_/chany_top_out[5]
+ sb_7__6_/chany_top_out[6] sb_7__6_/chany_top_out[7] sb_7__6_/chany_top_out[8] sb_7__6_/chany_top_out[9]
+ sb_7__6_/clk_1_E_out sb_7__6_/clk_1_N_in sb_7__6_/clk_1_W_out sb_7__6_/clk_2_E_out
+ sb_7__6_/clk_2_N_in sb_7__6_/clk_2_N_out sb_7__6_/clk_2_S_out sb_7__6_/clk_2_W_out
+ sb_7__6_/clk_3_E_out sb_7__6_/clk_3_N_in sb_7__6_/clk_3_N_out sb_7__6_/clk_3_S_out
+ sb_7__6_/clk_3_W_out sb_7__6_/left_bottom_grid_pin_34_ sb_7__6_/left_bottom_grid_pin_35_
+ sb_7__6_/left_bottom_grid_pin_36_ sb_7__6_/left_bottom_grid_pin_37_ sb_7__6_/left_bottom_grid_pin_38_
+ sb_7__6_/left_bottom_grid_pin_39_ sb_7__6_/left_bottom_grid_pin_40_ sb_7__6_/left_bottom_grid_pin_41_
+ sb_7__6_/prog_clk_0_N_in sb_7__6_/prog_clk_1_E_out sb_7__6_/prog_clk_1_N_in sb_7__6_/prog_clk_1_W_out
+ sb_7__6_/prog_clk_2_E_out sb_7__6_/prog_clk_2_N_in sb_7__6_/prog_clk_2_N_out sb_7__6_/prog_clk_2_S_out
+ sb_7__6_/prog_clk_2_W_out sb_7__6_/prog_clk_3_E_out sb_7__6_/prog_clk_3_N_in sb_7__6_/prog_clk_3_N_out
+ sb_7__6_/prog_clk_3_S_out sb_7__6_/prog_clk_3_W_out sb_7__6_/right_bottom_grid_pin_34_
+ sb_7__6_/right_bottom_grid_pin_35_ sb_7__6_/right_bottom_grid_pin_36_ sb_7__6_/right_bottom_grid_pin_37_
+ sb_7__6_/right_bottom_grid_pin_38_ sb_7__6_/right_bottom_grid_pin_39_ sb_7__6_/right_bottom_grid_pin_40_
+ sb_7__6_/right_bottom_grid_pin_41_ sb_7__6_/top_left_grid_pin_42_ sb_7__6_/top_left_grid_pin_43_
+ sb_7__6_/top_left_grid_pin_44_ sb_7__6_/top_left_grid_pin_45_ sb_7__6_/top_left_grid_pin_46_
+ sb_7__6_/top_left_grid_pin_47_ sb_7__6_/top_left_grid_pin_48_ sb_7__6_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_6__1_ cbx_6__0_/SC_OUT_TOP grid_clb_6__1_/SC_OUT_BOT cbx_6__1_/SC_IN_BOT
+ cby_5__1_/Test_en_E_out cby_6__1_/Test_en_W_in cby_5__1_/Test_en_E_out grid_clb_6__1_/Test_en_W_out
+ VGND VPWR grid_clb_6__1_/bottom_width_0_height_0__pin_50_ grid_clb_6__1_/bottom_width_0_height_0__pin_51_
+ cby_5__1_/ccff_tail cby_6__1_/ccff_head cbx_6__1_/clk_1_S_out cbx_6__1_/clk_1_S_out
+ cby_6__1_/prog_clk_0_W_in cbx_6__1_/prog_clk_1_S_out grid_clb_6__1_/prog_clk_0_N_out
+ cbx_6__1_/prog_clk_1_S_out cbx_6__0_/prog_clk_0_N_in grid_clb_6__1_/prog_clk_0_W_out
+ cby_6__1_/left_grid_pin_16_ cby_6__1_/left_grid_pin_17_ cby_6__1_/left_grid_pin_18_
+ cby_6__1_/left_grid_pin_19_ cby_6__1_/left_grid_pin_20_ cby_6__1_/left_grid_pin_21_
+ cby_6__1_/left_grid_pin_22_ cby_6__1_/left_grid_pin_23_ cby_6__1_/left_grid_pin_24_
+ cby_6__1_/left_grid_pin_25_ cby_6__1_/left_grid_pin_26_ cby_6__1_/left_grid_pin_27_
+ cby_6__1_/left_grid_pin_28_ cby_6__1_/left_grid_pin_29_ cby_6__1_/left_grid_pin_30_
+ cby_6__1_/left_grid_pin_31_ sb_6__0_/top_left_grid_pin_42_ sb_6__1_/bottom_left_grid_pin_42_
+ sb_6__0_/top_left_grid_pin_43_ sb_6__1_/bottom_left_grid_pin_43_ sb_6__0_/top_left_grid_pin_44_
+ sb_6__1_/bottom_left_grid_pin_44_ sb_6__0_/top_left_grid_pin_45_ sb_6__1_/bottom_left_grid_pin_45_
+ sb_6__0_/top_left_grid_pin_46_ sb_6__1_/bottom_left_grid_pin_46_ sb_6__0_/top_left_grid_pin_47_
+ sb_6__1_/bottom_left_grid_pin_47_ sb_6__0_/top_left_grid_pin_48_ sb_6__1_/bottom_left_grid_pin_48_
+ sb_6__0_/top_left_grid_pin_49_ sb_6__1_/bottom_left_grid_pin_49_ cbx_6__1_/bottom_grid_pin_0_
+ cbx_6__1_/bottom_grid_pin_10_ cbx_6__1_/bottom_grid_pin_11_ cbx_6__1_/bottom_grid_pin_12_
+ cbx_6__1_/bottom_grid_pin_13_ cbx_6__1_/bottom_grid_pin_14_ cbx_6__1_/bottom_grid_pin_15_
+ cbx_6__1_/bottom_grid_pin_1_ cbx_6__1_/bottom_grid_pin_2_ cbx_6__1_/REGOUT_FEEDTHROUGH
+ grid_clb_6__1_/top_width_0_height_0__pin_33_ sb_6__1_/left_bottom_grid_pin_34_ sb_5__1_/right_bottom_grid_pin_34_
+ sb_6__1_/left_bottom_grid_pin_35_ sb_5__1_/right_bottom_grid_pin_35_ sb_6__1_/left_bottom_grid_pin_36_
+ sb_5__1_/right_bottom_grid_pin_36_ sb_6__1_/left_bottom_grid_pin_37_ sb_5__1_/right_bottom_grid_pin_37_
+ sb_6__1_/left_bottom_grid_pin_38_ sb_5__1_/right_bottom_grid_pin_38_ sb_6__1_/left_bottom_grid_pin_39_
+ sb_5__1_/right_bottom_grid_pin_39_ cbx_6__1_/bottom_grid_pin_3_ sb_6__1_/left_bottom_grid_pin_40_
+ sb_5__1_/right_bottom_grid_pin_40_ sb_6__1_/left_bottom_grid_pin_41_ sb_5__1_/right_bottom_grid_pin_41_
+ cbx_6__1_/bottom_grid_pin_4_ cbx_6__1_/bottom_grid_pin_5_ cbx_6__1_/bottom_grid_pin_6_
+ cbx_6__1_/bottom_grid_pin_7_ cbx_6__1_/bottom_grid_pin_8_ cbx_6__1_/bottom_grid_pin_9_
+ grid_clb
Xsb_4__3_ sb_4__3_/Test_en_N_out sb_4__3_/Test_en_S_in VGND VPWR sb_4__3_/bottom_left_grid_pin_42_
+ sb_4__3_/bottom_left_grid_pin_43_ sb_4__3_/bottom_left_grid_pin_44_ sb_4__3_/bottom_left_grid_pin_45_
+ sb_4__3_/bottom_left_grid_pin_46_ sb_4__3_/bottom_left_grid_pin_47_ sb_4__3_/bottom_left_grid_pin_48_
+ sb_4__3_/bottom_left_grid_pin_49_ sb_4__3_/ccff_head sb_4__3_/ccff_tail sb_4__3_/chanx_left_in[0]
+ sb_4__3_/chanx_left_in[10] sb_4__3_/chanx_left_in[11] sb_4__3_/chanx_left_in[12]
+ sb_4__3_/chanx_left_in[13] sb_4__3_/chanx_left_in[14] sb_4__3_/chanx_left_in[15]
+ sb_4__3_/chanx_left_in[16] sb_4__3_/chanx_left_in[17] sb_4__3_/chanx_left_in[18]
+ sb_4__3_/chanx_left_in[19] sb_4__3_/chanx_left_in[1] sb_4__3_/chanx_left_in[2] sb_4__3_/chanx_left_in[3]
+ sb_4__3_/chanx_left_in[4] sb_4__3_/chanx_left_in[5] sb_4__3_/chanx_left_in[6] sb_4__3_/chanx_left_in[7]
+ sb_4__3_/chanx_left_in[8] sb_4__3_/chanx_left_in[9] sb_4__3_/chanx_left_out[0] sb_4__3_/chanx_left_out[10]
+ sb_4__3_/chanx_left_out[11] sb_4__3_/chanx_left_out[12] sb_4__3_/chanx_left_out[13]
+ sb_4__3_/chanx_left_out[14] sb_4__3_/chanx_left_out[15] sb_4__3_/chanx_left_out[16]
+ sb_4__3_/chanx_left_out[17] sb_4__3_/chanx_left_out[18] sb_4__3_/chanx_left_out[19]
+ sb_4__3_/chanx_left_out[1] sb_4__3_/chanx_left_out[2] sb_4__3_/chanx_left_out[3]
+ sb_4__3_/chanx_left_out[4] sb_4__3_/chanx_left_out[5] sb_4__3_/chanx_left_out[6]
+ sb_4__3_/chanx_left_out[7] sb_4__3_/chanx_left_out[8] sb_4__3_/chanx_left_out[9]
+ sb_4__3_/chanx_right_in[0] sb_4__3_/chanx_right_in[10] sb_4__3_/chanx_right_in[11]
+ sb_4__3_/chanx_right_in[12] sb_4__3_/chanx_right_in[13] sb_4__3_/chanx_right_in[14]
+ sb_4__3_/chanx_right_in[15] sb_4__3_/chanx_right_in[16] sb_4__3_/chanx_right_in[17]
+ sb_4__3_/chanx_right_in[18] sb_4__3_/chanx_right_in[19] sb_4__3_/chanx_right_in[1]
+ sb_4__3_/chanx_right_in[2] sb_4__3_/chanx_right_in[3] sb_4__3_/chanx_right_in[4]
+ sb_4__3_/chanx_right_in[5] sb_4__3_/chanx_right_in[6] sb_4__3_/chanx_right_in[7]
+ sb_4__3_/chanx_right_in[8] sb_4__3_/chanx_right_in[9] cbx_5__3_/chanx_left_in[0]
+ cbx_5__3_/chanx_left_in[10] cbx_5__3_/chanx_left_in[11] cbx_5__3_/chanx_left_in[12]
+ cbx_5__3_/chanx_left_in[13] cbx_5__3_/chanx_left_in[14] cbx_5__3_/chanx_left_in[15]
+ cbx_5__3_/chanx_left_in[16] cbx_5__3_/chanx_left_in[17] cbx_5__3_/chanx_left_in[18]
+ cbx_5__3_/chanx_left_in[19] cbx_5__3_/chanx_left_in[1] cbx_5__3_/chanx_left_in[2]
+ cbx_5__3_/chanx_left_in[3] cbx_5__3_/chanx_left_in[4] cbx_5__3_/chanx_left_in[5]
+ cbx_5__3_/chanx_left_in[6] cbx_5__3_/chanx_left_in[7] cbx_5__3_/chanx_left_in[8]
+ cbx_5__3_/chanx_left_in[9] cby_4__3_/chany_top_out[0] cby_4__3_/chany_top_out[10]
+ cby_4__3_/chany_top_out[11] cby_4__3_/chany_top_out[12] cby_4__3_/chany_top_out[13]
+ cby_4__3_/chany_top_out[14] cby_4__3_/chany_top_out[15] cby_4__3_/chany_top_out[16]
+ cby_4__3_/chany_top_out[17] cby_4__3_/chany_top_out[18] cby_4__3_/chany_top_out[19]
+ cby_4__3_/chany_top_out[1] cby_4__3_/chany_top_out[2] cby_4__3_/chany_top_out[3]
+ cby_4__3_/chany_top_out[4] cby_4__3_/chany_top_out[5] cby_4__3_/chany_top_out[6]
+ cby_4__3_/chany_top_out[7] cby_4__3_/chany_top_out[8] cby_4__3_/chany_top_out[9]
+ cby_4__3_/chany_top_in[0] cby_4__3_/chany_top_in[10] cby_4__3_/chany_top_in[11]
+ cby_4__3_/chany_top_in[12] cby_4__3_/chany_top_in[13] cby_4__3_/chany_top_in[14]
+ cby_4__3_/chany_top_in[15] cby_4__3_/chany_top_in[16] cby_4__3_/chany_top_in[17]
+ cby_4__3_/chany_top_in[18] cby_4__3_/chany_top_in[19] cby_4__3_/chany_top_in[1]
+ cby_4__3_/chany_top_in[2] cby_4__3_/chany_top_in[3] cby_4__3_/chany_top_in[4] cby_4__3_/chany_top_in[5]
+ cby_4__3_/chany_top_in[6] cby_4__3_/chany_top_in[7] cby_4__3_/chany_top_in[8] cby_4__3_/chany_top_in[9]
+ sb_4__3_/chany_top_in[0] sb_4__3_/chany_top_in[10] sb_4__3_/chany_top_in[11] sb_4__3_/chany_top_in[12]
+ sb_4__3_/chany_top_in[13] sb_4__3_/chany_top_in[14] sb_4__3_/chany_top_in[15] sb_4__3_/chany_top_in[16]
+ sb_4__3_/chany_top_in[17] sb_4__3_/chany_top_in[18] sb_4__3_/chany_top_in[19] sb_4__3_/chany_top_in[1]
+ sb_4__3_/chany_top_in[2] sb_4__3_/chany_top_in[3] sb_4__3_/chany_top_in[4] sb_4__3_/chany_top_in[5]
+ sb_4__3_/chany_top_in[6] sb_4__3_/chany_top_in[7] sb_4__3_/chany_top_in[8] sb_4__3_/chany_top_in[9]
+ sb_4__3_/chany_top_out[0] sb_4__3_/chany_top_out[10] sb_4__3_/chany_top_out[11]
+ sb_4__3_/chany_top_out[12] sb_4__3_/chany_top_out[13] sb_4__3_/chany_top_out[14]
+ sb_4__3_/chany_top_out[15] sb_4__3_/chany_top_out[16] sb_4__3_/chany_top_out[17]
+ sb_4__3_/chany_top_out[18] sb_4__3_/chany_top_out[19] sb_4__3_/chany_top_out[1]
+ sb_4__3_/chany_top_out[2] sb_4__3_/chany_top_out[3] sb_4__3_/chany_top_out[4] sb_4__3_/chany_top_out[5]
+ sb_4__3_/chany_top_out[6] sb_4__3_/chany_top_out[7] sb_4__3_/chany_top_out[8] sb_4__3_/chany_top_out[9]
+ sb_4__3_/clk_1_E_out sb_4__3_/clk_1_N_in sb_4__3_/clk_1_W_out sb_4__3_/clk_2_E_out
+ sb_4__3_/clk_2_N_in sb_4__3_/clk_2_N_out sb_4__3_/clk_2_S_out sb_4__3_/clk_2_W_out
+ sb_4__3_/clk_3_E_out sb_4__3_/clk_3_N_in sb_4__3_/clk_3_N_out sb_4__3_/clk_3_S_out
+ sb_4__3_/clk_3_W_out sb_4__3_/left_bottom_grid_pin_34_ sb_4__3_/left_bottom_grid_pin_35_
+ sb_4__3_/left_bottom_grid_pin_36_ sb_4__3_/left_bottom_grid_pin_37_ sb_4__3_/left_bottom_grid_pin_38_
+ sb_4__3_/left_bottom_grid_pin_39_ sb_4__3_/left_bottom_grid_pin_40_ sb_4__3_/left_bottom_grid_pin_41_
+ sb_4__3_/prog_clk_0_N_in sb_4__3_/prog_clk_1_E_out sb_4__3_/prog_clk_1_N_in sb_4__3_/prog_clk_1_W_out
+ sb_4__3_/prog_clk_2_E_out sb_4__3_/prog_clk_2_N_in sb_4__3_/prog_clk_2_N_out sb_4__3_/prog_clk_2_S_out
+ sb_4__3_/prog_clk_2_W_out sb_4__3_/prog_clk_3_E_out sb_4__3_/prog_clk_3_N_in sb_4__3_/prog_clk_3_N_out
+ sb_4__3_/prog_clk_3_S_out sb_4__3_/prog_clk_3_W_out sb_4__3_/right_bottom_grid_pin_34_
+ sb_4__3_/right_bottom_grid_pin_35_ sb_4__3_/right_bottom_grid_pin_36_ sb_4__3_/right_bottom_grid_pin_37_
+ sb_4__3_/right_bottom_grid_pin_38_ sb_4__3_/right_bottom_grid_pin_39_ sb_4__3_/right_bottom_grid_pin_40_
+ sb_4__3_/right_bottom_grid_pin_41_ sb_4__3_/top_left_grid_pin_42_ sb_4__3_/top_left_grid_pin_43_
+ sb_4__3_/top_left_grid_pin_44_ sb_4__3_/top_left_grid_pin_45_ sb_4__3_/top_left_grid_pin_46_
+ sb_4__3_/top_left_grid_pin_47_ sb_4__3_/top_left_grid_pin_48_ sb_4__3_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_1__0_ sb_1__0_/SC_IN_TOP sb_1__0_/SC_OUT_TOP sb_1__0_/Test_en_N_out sb_1__0_/Test_en_S_in
+ VGND VPWR sb_1__0_/ccff_head sb_1__0_/ccff_tail sb_1__0_/chanx_left_in[0] sb_1__0_/chanx_left_in[10]
+ sb_1__0_/chanx_left_in[11] sb_1__0_/chanx_left_in[12] sb_1__0_/chanx_left_in[13]
+ sb_1__0_/chanx_left_in[14] sb_1__0_/chanx_left_in[15] sb_1__0_/chanx_left_in[16]
+ sb_1__0_/chanx_left_in[17] sb_1__0_/chanx_left_in[18] sb_1__0_/chanx_left_in[19]
+ sb_1__0_/chanx_left_in[1] sb_1__0_/chanx_left_in[2] sb_1__0_/chanx_left_in[3] sb_1__0_/chanx_left_in[4]
+ sb_1__0_/chanx_left_in[5] sb_1__0_/chanx_left_in[6] sb_1__0_/chanx_left_in[7] sb_1__0_/chanx_left_in[8]
+ sb_1__0_/chanx_left_in[9] sb_1__0_/chanx_left_out[0] sb_1__0_/chanx_left_out[10]
+ sb_1__0_/chanx_left_out[11] sb_1__0_/chanx_left_out[12] sb_1__0_/chanx_left_out[13]
+ sb_1__0_/chanx_left_out[14] sb_1__0_/chanx_left_out[15] sb_1__0_/chanx_left_out[16]
+ sb_1__0_/chanx_left_out[17] sb_1__0_/chanx_left_out[18] sb_1__0_/chanx_left_out[19]
+ sb_1__0_/chanx_left_out[1] sb_1__0_/chanx_left_out[2] sb_1__0_/chanx_left_out[3]
+ sb_1__0_/chanx_left_out[4] sb_1__0_/chanx_left_out[5] sb_1__0_/chanx_left_out[6]
+ sb_1__0_/chanx_left_out[7] sb_1__0_/chanx_left_out[8] sb_1__0_/chanx_left_out[9]
+ sb_1__0_/chanx_right_in[0] sb_1__0_/chanx_right_in[10] sb_1__0_/chanx_right_in[11]
+ sb_1__0_/chanx_right_in[12] sb_1__0_/chanx_right_in[13] sb_1__0_/chanx_right_in[14]
+ sb_1__0_/chanx_right_in[15] sb_1__0_/chanx_right_in[16] sb_1__0_/chanx_right_in[17]
+ sb_1__0_/chanx_right_in[18] sb_1__0_/chanx_right_in[19] sb_1__0_/chanx_right_in[1]
+ sb_1__0_/chanx_right_in[2] sb_1__0_/chanx_right_in[3] sb_1__0_/chanx_right_in[4]
+ sb_1__0_/chanx_right_in[5] sb_1__0_/chanx_right_in[6] sb_1__0_/chanx_right_in[7]
+ sb_1__0_/chanx_right_in[8] sb_1__0_/chanx_right_in[9] cbx_2__0_/chanx_left_in[0]
+ cbx_2__0_/chanx_left_in[10] cbx_2__0_/chanx_left_in[11] cbx_2__0_/chanx_left_in[12]
+ cbx_2__0_/chanx_left_in[13] cbx_2__0_/chanx_left_in[14] cbx_2__0_/chanx_left_in[15]
+ cbx_2__0_/chanx_left_in[16] cbx_2__0_/chanx_left_in[17] cbx_2__0_/chanx_left_in[18]
+ cbx_2__0_/chanx_left_in[19] cbx_2__0_/chanx_left_in[1] cbx_2__0_/chanx_left_in[2]
+ cbx_2__0_/chanx_left_in[3] cbx_2__0_/chanx_left_in[4] cbx_2__0_/chanx_left_in[5]
+ cbx_2__0_/chanx_left_in[6] cbx_2__0_/chanx_left_in[7] cbx_2__0_/chanx_left_in[8]
+ cbx_2__0_/chanx_left_in[9] sb_1__0_/chany_top_in[0] sb_1__0_/chany_top_in[10] sb_1__0_/chany_top_in[11]
+ sb_1__0_/chany_top_in[12] sb_1__0_/chany_top_in[13] sb_1__0_/chany_top_in[14] sb_1__0_/chany_top_in[15]
+ sb_1__0_/chany_top_in[16] sb_1__0_/chany_top_in[17] sb_1__0_/chany_top_in[18] sb_1__0_/chany_top_in[19]
+ sb_1__0_/chany_top_in[1] sb_1__0_/chany_top_in[2] sb_1__0_/chany_top_in[3] sb_1__0_/chany_top_in[4]
+ sb_1__0_/chany_top_in[5] sb_1__0_/chany_top_in[6] sb_1__0_/chany_top_in[7] sb_1__0_/chany_top_in[8]
+ sb_1__0_/chany_top_in[9] sb_1__0_/chany_top_out[0] sb_1__0_/chany_top_out[10] sb_1__0_/chany_top_out[11]
+ sb_1__0_/chany_top_out[12] sb_1__0_/chany_top_out[13] sb_1__0_/chany_top_out[14]
+ sb_1__0_/chany_top_out[15] sb_1__0_/chany_top_out[16] sb_1__0_/chany_top_out[17]
+ sb_1__0_/chany_top_out[18] sb_1__0_/chany_top_out[19] sb_1__0_/chany_top_out[1]
+ sb_1__0_/chany_top_out[2] sb_1__0_/chany_top_out[3] sb_1__0_/chany_top_out[4] sb_1__0_/chany_top_out[5]
+ sb_1__0_/chany_top_out[6] sb_1__0_/chany_top_out[7] sb_1__0_/chany_top_out[8] sb_1__0_/chany_top_out[9]
+ sb_1__0_/clk_3_N_out sb_1__0_/clk_3_S_in sb_1__0_/left_bottom_grid_pin_11_ sb_1__0_/left_bottom_grid_pin_13_
+ sb_1__0_/left_bottom_grid_pin_15_ sb_1__0_/left_bottom_grid_pin_17_ sb_1__0_/left_bottom_grid_pin_1_
+ sb_1__0_/left_bottom_grid_pin_3_ sb_1__0_/left_bottom_grid_pin_5_ sb_1__0_/left_bottom_grid_pin_7_
+ sb_1__0_/left_bottom_grid_pin_9_ sb_1__0_/prog_clk_0_N_in sb_1__0_/prog_clk_3_N_out
+ sb_1__0_/prog_clk_3_S_in sb_1__0_/right_bottom_grid_pin_11_ sb_1__0_/right_bottom_grid_pin_13_
+ sb_1__0_/right_bottom_grid_pin_15_ sb_1__0_/right_bottom_grid_pin_17_ sb_1__0_/right_bottom_grid_pin_1_
+ sb_1__0_/right_bottom_grid_pin_3_ sb_1__0_/right_bottom_grid_pin_5_ sb_1__0_/right_bottom_grid_pin_7_
+ sb_1__0_/right_bottom_grid_pin_9_ sb_1__0_/top_left_grid_pin_42_ sb_1__0_/top_left_grid_pin_43_
+ sb_1__0_/top_left_grid_pin_44_ sb_1__0_/top_left_grid_pin_45_ sb_1__0_/top_left_grid_pin_46_
+ sb_1__0_/top_left_grid_pin_47_ sb_1__0_/top_left_grid_pin_48_ sb_1__0_/top_left_grid_pin_49_
+ sb_1__0_
Xcby_3__7_ cby_3__7_/Test_en_W_in cby_3__7_/Test_en_E_out cby_3__7_/Test_en_N_out
+ cby_3__7_/Test_en_W_in cby_3__7_/Test_en_W_in cby_3__7_/Test_en_W_out VGND VPWR
+ cby_3__7_/ccff_head cby_3__7_/ccff_tail sb_3__6_/chany_top_out[0] sb_3__6_/chany_top_out[10]
+ sb_3__6_/chany_top_out[11] sb_3__6_/chany_top_out[12] sb_3__6_/chany_top_out[13]
+ sb_3__6_/chany_top_out[14] sb_3__6_/chany_top_out[15] sb_3__6_/chany_top_out[16]
+ sb_3__6_/chany_top_out[17] sb_3__6_/chany_top_out[18] sb_3__6_/chany_top_out[19]
+ sb_3__6_/chany_top_out[1] sb_3__6_/chany_top_out[2] sb_3__6_/chany_top_out[3] sb_3__6_/chany_top_out[4]
+ sb_3__6_/chany_top_out[5] sb_3__6_/chany_top_out[6] sb_3__6_/chany_top_out[7] sb_3__6_/chany_top_out[8]
+ sb_3__6_/chany_top_out[9] sb_3__6_/chany_top_in[0] sb_3__6_/chany_top_in[10] sb_3__6_/chany_top_in[11]
+ sb_3__6_/chany_top_in[12] sb_3__6_/chany_top_in[13] sb_3__6_/chany_top_in[14] sb_3__6_/chany_top_in[15]
+ sb_3__6_/chany_top_in[16] sb_3__6_/chany_top_in[17] sb_3__6_/chany_top_in[18] sb_3__6_/chany_top_in[19]
+ sb_3__6_/chany_top_in[1] sb_3__6_/chany_top_in[2] sb_3__6_/chany_top_in[3] sb_3__6_/chany_top_in[4]
+ sb_3__6_/chany_top_in[5] sb_3__6_/chany_top_in[6] sb_3__6_/chany_top_in[7] sb_3__6_/chany_top_in[8]
+ sb_3__6_/chany_top_in[9] cby_3__7_/chany_top_in[0] cby_3__7_/chany_top_in[10] cby_3__7_/chany_top_in[11]
+ cby_3__7_/chany_top_in[12] cby_3__7_/chany_top_in[13] cby_3__7_/chany_top_in[14]
+ cby_3__7_/chany_top_in[15] cby_3__7_/chany_top_in[16] cby_3__7_/chany_top_in[17]
+ cby_3__7_/chany_top_in[18] cby_3__7_/chany_top_in[19] cby_3__7_/chany_top_in[1]
+ cby_3__7_/chany_top_in[2] cby_3__7_/chany_top_in[3] cby_3__7_/chany_top_in[4] cby_3__7_/chany_top_in[5]
+ cby_3__7_/chany_top_in[6] cby_3__7_/chany_top_in[7] cby_3__7_/chany_top_in[8] cby_3__7_/chany_top_in[9]
+ cby_3__7_/chany_top_out[0] cby_3__7_/chany_top_out[10] cby_3__7_/chany_top_out[11]
+ cby_3__7_/chany_top_out[12] cby_3__7_/chany_top_out[13] cby_3__7_/chany_top_out[14]
+ cby_3__7_/chany_top_out[15] cby_3__7_/chany_top_out[16] cby_3__7_/chany_top_out[17]
+ cby_3__7_/chany_top_out[18] cby_3__7_/chany_top_out[19] cby_3__7_/chany_top_out[1]
+ cby_3__7_/chany_top_out[2] cby_3__7_/chany_top_out[3] cby_3__7_/chany_top_out[4]
+ cby_3__7_/chany_top_out[5] cby_3__7_/chany_top_out[6] cby_3__7_/chany_top_out[7]
+ cby_3__7_/chany_top_out[8] cby_3__7_/chany_top_out[9] sb_3__7_/clk_1_N_in sb_3__6_/clk_2_N_out
+ cby_3__7_/clk_2_S_out cby_3__7_/clk_3_N_out cby_3__7_/clk_3_S_in cby_3__7_/clk_3_S_out
+ cby_3__7_/left_grid_pin_16_ cby_3__7_/left_grid_pin_17_ cby_3__7_/left_grid_pin_18_
+ cby_3__7_/left_grid_pin_19_ cby_3__7_/left_grid_pin_20_ cby_3__7_/left_grid_pin_21_
+ cby_3__7_/left_grid_pin_22_ cby_3__7_/left_grid_pin_23_ cby_3__7_/left_grid_pin_24_
+ cby_3__7_/left_grid_pin_25_ cby_3__7_/left_grid_pin_26_ cby_3__7_/left_grid_pin_27_
+ cby_3__7_/left_grid_pin_28_ cby_3__7_/left_grid_pin_29_ cby_3__7_/left_grid_pin_30_
+ cby_3__7_/left_grid_pin_31_ cby_3__7_/prog_clk_0_N_out sb_3__6_/prog_clk_0_N_in
+ cby_3__7_/prog_clk_0_W_in sb_3__7_/prog_clk_1_N_in sb_3__6_/prog_clk_2_N_out cby_3__7_/prog_clk_2_S_out
+ cby_3__7_/prog_clk_3_N_out cby_3__7_/prog_clk_3_S_in cby_3__7_/prog_clk_3_S_out
+ cby_1__1_
Xcby_0__4_ IO_ISOL_N VGND VPWR sb_0__4_/ccff_tail cby_0__4_/ccff_tail sb_0__3_/chany_top_out[0]
+ sb_0__3_/chany_top_out[10] sb_0__3_/chany_top_out[11] sb_0__3_/chany_top_out[12]
+ sb_0__3_/chany_top_out[13] sb_0__3_/chany_top_out[14] sb_0__3_/chany_top_out[15]
+ sb_0__3_/chany_top_out[16] sb_0__3_/chany_top_out[17] sb_0__3_/chany_top_out[18]
+ sb_0__3_/chany_top_out[19] sb_0__3_/chany_top_out[1] sb_0__3_/chany_top_out[2] sb_0__3_/chany_top_out[3]
+ sb_0__3_/chany_top_out[4] sb_0__3_/chany_top_out[5] sb_0__3_/chany_top_out[6] sb_0__3_/chany_top_out[7]
+ sb_0__3_/chany_top_out[8] sb_0__3_/chany_top_out[9] sb_0__3_/chany_top_in[0] sb_0__3_/chany_top_in[10]
+ sb_0__3_/chany_top_in[11] sb_0__3_/chany_top_in[12] sb_0__3_/chany_top_in[13] sb_0__3_/chany_top_in[14]
+ sb_0__3_/chany_top_in[15] sb_0__3_/chany_top_in[16] sb_0__3_/chany_top_in[17] sb_0__3_/chany_top_in[18]
+ sb_0__3_/chany_top_in[19] sb_0__3_/chany_top_in[1] sb_0__3_/chany_top_in[2] sb_0__3_/chany_top_in[3]
+ sb_0__3_/chany_top_in[4] sb_0__3_/chany_top_in[5] sb_0__3_/chany_top_in[6] sb_0__3_/chany_top_in[7]
+ sb_0__3_/chany_top_in[8] sb_0__3_/chany_top_in[9] cby_0__4_/chany_top_in[0] cby_0__4_/chany_top_in[10]
+ cby_0__4_/chany_top_in[11] cby_0__4_/chany_top_in[12] cby_0__4_/chany_top_in[13]
+ cby_0__4_/chany_top_in[14] cby_0__4_/chany_top_in[15] cby_0__4_/chany_top_in[16]
+ cby_0__4_/chany_top_in[17] cby_0__4_/chany_top_in[18] cby_0__4_/chany_top_in[19]
+ cby_0__4_/chany_top_in[1] cby_0__4_/chany_top_in[2] cby_0__4_/chany_top_in[3] cby_0__4_/chany_top_in[4]
+ cby_0__4_/chany_top_in[5] cby_0__4_/chany_top_in[6] cby_0__4_/chany_top_in[7] cby_0__4_/chany_top_in[8]
+ cby_0__4_/chany_top_in[9] cby_0__4_/chany_top_out[0] cby_0__4_/chany_top_out[10]
+ cby_0__4_/chany_top_out[11] cby_0__4_/chany_top_out[12] cby_0__4_/chany_top_out[13]
+ cby_0__4_/chany_top_out[14] cby_0__4_/chany_top_out[15] cby_0__4_/chany_top_out[16]
+ cby_0__4_/chany_top_out[17] cby_0__4_/chany_top_out[18] cby_0__4_/chany_top_out[19]
+ cby_0__4_/chany_top_out[1] cby_0__4_/chany_top_out[2] cby_0__4_/chany_top_out[3]
+ cby_0__4_/chany_top_out[4] cby_0__4_/chany_top_out[5] cby_0__4_/chany_top_out[6]
+ cby_0__4_/chany_top_out[7] cby_0__4_/chany_top_out[8] cby_0__4_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
+ cby_0__4_/left_grid_pin_0_ cby_0__4_/prog_clk_0_E_in cby_0__4_/left_grid_pin_0_
+ sb_0__3_/top_left_grid_pin_1_ sb_0__4_/bottom_left_grid_pin_1_ cby_0__1_
Xcbx_7__0_ IO_ISOL_N cbx_7__0_/SC_IN_BOT cbx_7__0_/SC_IN_TOP sb_7__0_/SC_IN_TOP cbx_7__0_/SC_OUT_TOP
+ VGND VPWR cbx_7__0_/bottom_grid_pin_0_ cbx_7__0_/bottom_grid_pin_10_ cbx_7__0_/bottom_grid_pin_12_
+ cbx_7__0_/bottom_grid_pin_14_ cbx_7__0_/bottom_grid_pin_16_ cbx_7__0_/bottom_grid_pin_2_
+ cbx_7__0_/bottom_grid_pin_4_ cbx_7__0_/bottom_grid_pin_6_ cbx_7__0_/bottom_grid_pin_8_
+ sb_7__0_/ccff_tail sb_6__0_/ccff_head cbx_7__0_/chanx_left_in[0] cbx_7__0_/chanx_left_in[10]
+ cbx_7__0_/chanx_left_in[11] cbx_7__0_/chanx_left_in[12] cbx_7__0_/chanx_left_in[13]
+ cbx_7__0_/chanx_left_in[14] cbx_7__0_/chanx_left_in[15] cbx_7__0_/chanx_left_in[16]
+ cbx_7__0_/chanx_left_in[17] cbx_7__0_/chanx_left_in[18] cbx_7__0_/chanx_left_in[19]
+ cbx_7__0_/chanx_left_in[1] cbx_7__0_/chanx_left_in[2] cbx_7__0_/chanx_left_in[3]
+ cbx_7__0_/chanx_left_in[4] cbx_7__0_/chanx_left_in[5] cbx_7__0_/chanx_left_in[6]
+ cbx_7__0_/chanx_left_in[7] cbx_7__0_/chanx_left_in[8] cbx_7__0_/chanx_left_in[9]
+ sb_6__0_/chanx_right_in[0] sb_6__0_/chanx_right_in[10] sb_6__0_/chanx_right_in[11]
+ sb_6__0_/chanx_right_in[12] sb_6__0_/chanx_right_in[13] sb_6__0_/chanx_right_in[14]
+ sb_6__0_/chanx_right_in[15] sb_6__0_/chanx_right_in[16] sb_6__0_/chanx_right_in[17]
+ sb_6__0_/chanx_right_in[18] sb_6__0_/chanx_right_in[19] sb_6__0_/chanx_right_in[1]
+ sb_6__0_/chanx_right_in[2] sb_6__0_/chanx_right_in[3] sb_6__0_/chanx_right_in[4]
+ sb_6__0_/chanx_right_in[5] sb_6__0_/chanx_right_in[6] sb_6__0_/chanx_right_in[7]
+ sb_6__0_/chanx_right_in[8] sb_6__0_/chanx_right_in[9] sb_7__0_/chanx_left_out[0]
+ sb_7__0_/chanx_left_out[10] sb_7__0_/chanx_left_out[11] sb_7__0_/chanx_left_out[12]
+ sb_7__0_/chanx_left_out[13] sb_7__0_/chanx_left_out[14] sb_7__0_/chanx_left_out[15]
+ sb_7__0_/chanx_left_out[16] sb_7__0_/chanx_left_out[17] sb_7__0_/chanx_left_out[18]
+ sb_7__0_/chanx_left_out[19] sb_7__0_/chanx_left_out[1] sb_7__0_/chanx_left_out[2]
+ sb_7__0_/chanx_left_out[3] sb_7__0_/chanx_left_out[4] sb_7__0_/chanx_left_out[5]
+ sb_7__0_/chanx_left_out[6] sb_7__0_/chanx_left_out[7] sb_7__0_/chanx_left_out[8]
+ sb_7__0_/chanx_left_out[9] sb_7__0_/chanx_left_in[0] sb_7__0_/chanx_left_in[10]
+ sb_7__0_/chanx_left_in[11] sb_7__0_/chanx_left_in[12] sb_7__0_/chanx_left_in[13]
+ sb_7__0_/chanx_left_in[14] sb_7__0_/chanx_left_in[15] sb_7__0_/chanx_left_in[16]
+ sb_7__0_/chanx_left_in[17] sb_7__0_/chanx_left_in[18] sb_7__0_/chanx_left_in[19]
+ sb_7__0_/chanx_left_in[1] sb_7__0_/chanx_left_in[2] sb_7__0_/chanx_left_in[3] sb_7__0_/chanx_left_in[4]
+ sb_7__0_/chanx_left_in[5] sb_7__0_/chanx_left_in[6] sb_7__0_/chanx_left_in[7] sb_7__0_/chanx_left_in[8]
+ sb_7__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33] cbx_7__0_/prog_clk_0_N_in cbx_7__0_/prog_clk_0_W_out
+ cbx_7__0_/bottom_grid_pin_0_ cbx_7__0_/bottom_grid_pin_10_ sb_7__0_/left_bottom_grid_pin_11_
+ sb_6__0_/right_bottom_grid_pin_11_ cbx_7__0_/bottom_grid_pin_12_ sb_7__0_/left_bottom_grid_pin_13_
+ sb_6__0_/right_bottom_grid_pin_13_ cbx_7__0_/bottom_grid_pin_14_ sb_7__0_/left_bottom_grid_pin_15_
+ sb_6__0_/right_bottom_grid_pin_15_ cbx_7__0_/bottom_grid_pin_16_ sb_7__0_/left_bottom_grid_pin_17_
+ sb_6__0_/right_bottom_grid_pin_17_ sb_7__0_/left_bottom_grid_pin_1_ sb_6__0_/right_bottom_grid_pin_1_
+ cbx_7__0_/bottom_grid_pin_2_ sb_7__0_/left_bottom_grid_pin_3_ sb_6__0_/right_bottom_grid_pin_3_
+ cbx_7__0_/bottom_grid_pin_4_ sb_7__0_/left_bottom_grid_pin_5_ sb_6__0_/right_bottom_grid_pin_5_
+ cbx_7__0_/bottom_grid_pin_6_ sb_7__0_/left_bottom_grid_pin_7_ sb_6__0_/right_bottom_grid_pin_7_
+ cbx_7__0_/bottom_grid_pin_8_ sb_7__0_/left_bottom_grid_pin_9_ sb_6__0_/right_bottom_grid_pin_9_
+ cbx_1__0_
Xcbx_3__8_ IO_ISOL_N cbx_3__8_/SC_IN_BOT sb_2__8_/SC_OUT_BOT cbx_3__8_/SC_OUT_BOT
+ cbx_3__8_/SC_OUT_TOP VGND VPWR cbx_3__8_/bottom_grid_pin_0_ cbx_3__8_/bottom_grid_pin_10_
+ cbx_3__8_/bottom_grid_pin_11_ cbx_3__8_/bottom_grid_pin_12_ cbx_3__8_/bottom_grid_pin_13_
+ cbx_3__8_/bottom_grid_pin_14_ cbx_3__8_/bottom_grid_pin_15_ cbx_3__8_/bottom_grid_pin_1_
+ cbx_3__8_/bottom_grid_pin_2_ cbx_3__8_/bottom_grid_pin_3_ cbx_3__8_/bottom_grid_pin_4_
+ cbx_3__8_/bottom_grid_pin_5_ cbx_3__8_/bottom_grid_pin_6_ cbx_3__8_/bottom_grid_pin_7_
+ cbx_3__8_/bottom_grid_pin_8_ cbx_3__8_/bottom_grid_pin_9_ cbx_3__8_/top_grid_pin_0_
+ sb_3__8_/left_top_grid_pin_1_ sb_2__8_/right_top_grid_pin_1_ sb_3__8_/ccff_tail
+ sb_2__8_/ccff_head cbx_3__8_/chanx_left_in[0] cbx_3__8_/chanx_left_in[10] cbx_3__8_/chanx_left_in[11]
+ cbx_3__8_/chanx_left_in[12] cbx_3__8_/chanx_left_in[13] cbx_3__8_/chanx_left_in[14]
+ cbx_3__8_/chanx_left_in[15] cbx_3__8_/chanx_left_in[16] cbx_3__8_/chanx_left_in[17]
+ cbx_3__8_/chanx_left_in[18] cbx_3__8_/chanx_left_in[19] cbx_3__8_/chanx_left_in[1]
+ cbx_3__8_/chanx_left_in[2] cbx_3__8_/chanx_left_in[3] cbx_3__8_/chanx_left_in[4]
+ cbx_3__8_/chanx_left_in[5] cbx_3__8_/chanx_left_in[6] cbx_3__8_/chanx_left_in[7]
+ cbx_3__8_/chanx_left_in[8] cbx_3__8_/chanx_left_in[9] sb_2__8_/chanx_right_in[0]
+ sb_2__8_/chanx_right_in[10] sb_2__8_/chanx_right_in[11] sb_2__8_/chanx_right_in[12]
+ sb_2__8_/chanx_right_in[13] sb_2__8_/chanx_right_in[14] sb_2__8_/chanx_right_in[15]
+ sb_2__8_/chanx_right_in[16] sb_2__8_/chanx_right_in[17] sb_2__8_/chanx_right_in[18]
+ sb_2__8_/chanx_right_in[19] sb_2__8_/chanx_right_in[1] sb_2__8_/chanx_right_in[2]
+ sb_2__8_/chanx_right_in[3] sb_2__8_/chanx_right_in[4] sb_2__8_/chanx_right_in[5]
+ sb_2__8_/chanx_right_in[6] sb_2__8_/chanx_right_in[7] sb_2__8_/chanx_right_in[8]
+ sb_2__8_/chanx_right_in[9] sb_3__8_/chanx_left_out[0] sb_3__8_/chanx_left_out[10]
+ sb_3__8_/chanx_left_out[11] sb_3__8_/chanx_left_out[12] sb_3__8_/chanx_left_out[13]
+ sb_3__8_/chanx_left_out[14] sb_3__8_/chanx_left_out[15] sb_3__8_/chanx_left_out[16]
+ sb_3__8_/chanx_left_out[17] sb_3__8_/chanx_left_out[18] sb_3__8_/chanx_left_out[19]
+ sb_3__8_/chanx_left_out[1] sb_3__8_/chanx_left_out[2] sb_3__8_/chanx_left_out[3]
+ sb_3__8_/chanx_left_out[4] sb_3__8_/chanx_left_out[5] sb_3__8_/chanx_left_out[6]
+ sb_3__8_/chanx_left_out[7] sb_3__8_/chanx_left_out[8] sb_3__8_/chanx_left_out[9]
+ sb_3__8_/chanx_left_in[0] sb_3__8_/chanx_left_in[10] sb_3__8_/chanx_left_in[11]
+ sb_3__8_/chanx_left_in[12] sb_3__8_/chanx_left_in[13] sb_3__8_/chanx_left_in[14]
+ sb_3__8_/chanx_left_in[15] sb_3__8_/chanx_left_in[16] sb_3__8_/chanx_left_in[17]
+ sb_3__8_/chanx_left_in[18] sb_3__8_/chanx_left_in[19] sb_3__8_/chanx_left_in[1]
+ sb_3__8_/chanx_left_in[2] sb_3__8_/chanx_left_in[3] sb_3__8_/chanx_left_in[4] sb_3__8_/chanx_left_in[5]
+ sb_3__8_/chanx_left_in[6] sb_3__8_/chanx_left_in[7] sb_3__8_/chanx_left_in[8] sb_3__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
+ cbx_3__8_/prog_clk_0_S_in cbx_3__8_/prog_clk_0_W_out cbx_3__8_/top_grid_pin_0_ cbx_1__2_
Xgrid_clb_2__8_ cbx_2__7_/SC_OUT_TOP grid_clb_2__8_/SC_OUT_BOT cbx_2__8_/SC_IN_BOT
+ cby_2__8_/Test_en_W_out grid_clb_2__8_/Test_en_E_out cby_2__8_/Test_en_W_out cby_1__8_/Test_en_W_in
+ VGND VPWR cbx_2__7_/REGIN_FEEDTHROUGH grid_clb_2__8_/bottom_width_0_height_0__pin_51_
+ cby_1__8_/ccff_tail cby_2__8_/ccff_head cbx_2__7_/clk_1_N_out cbx_2__7_/clk_1_N_out
+ cby_2__8_/prog_clk_0_W_in cbx_2__7_/prog_clk_1_N_out cbx_2__8_/prog_clk_0_S_in cbx_2__7_/prog_clk_1_N_out
+ cbx_2__7_/prog_clk_0_N_in grid_clb_2__8_/prog_clk_0_W_out cby_2__8_/left_grid_pin_16_
+ cby_2__8_/left_grid_pin_17_ cby_2__8_/left_grid_pin_18_ cby_2__8_/left_grid_pin_19_
+ cby_2__8_/left_grid_pin_20_ cby_2__8_/left_grid_pin_21_ cby_2__8_/left_grid_pin_22_
+ cby_2__8_/left_grid_pin_23_ cby_2__8_/left_grid_pin_24_ cby_2__8_/left_grid_pin_25_
+ cby_2__8_/left_grid_pin_26_ cby_2__8_/left_grid_pin_27_ cby_2__8_/left_grid_pin_28_
+ cby_2__8_/left_grid_pin_29_ cby_2__8_/left_grid_pin_30_ cby_2__8_/left_grid_pin_31_
+ sb_2__7_/top_left_grid_pin_42_ sb_2__8_/bottom_left_grid_pin_42_ sb_2__7_/top_left_grid_pin_43_
+ sb_2__8_/bottom_left_grid_pin_43_ sb_2__7_/top_left_grid_pin_44_ sb_2__8_/bottom_left_grid_pin_44_
+ sb_2__7_/top_left_grid_pin_45_ sb_2__8_/bottom_left_grid_pin_45_ sb_2__7_/top_left_grid_pin_46_
+ sb_2__8_/bottom_left_grid_pin_46_ sb_2__7_/top_left_grid_pin_47_ sb_2__8_/bottom_left_grid_pin_47_
+ sb_2__7_/top_left_grid_pin_48_ sb_2__8_/bottom_left_grid_pin_48_ sb_2__7_/top_left_grid_pin_49_
+ sb_2__8_/bottom_left_grid_pin_49_ cbx_2__8_/bottom_grid_pin_0_ cbx_2__8_/bottom_grid_pin_10_
+ cbx_2__8_/bottom_grid_pin_11_ cbx_2__8_/bottom_grid_pin_12_ cbx_2__8_/bottom_grid_pin_13_
+ cbx_2__8_/bottom_grid_pin_14_ cbx_2__8_/bottom_grid_pin_15_ cbx_2__8_/bottom_grid_pin_1_
+ cbx_2__8_/bottom_grid_pin_2_ tie_array/x[1] grid_clb_2__8_/top_width_0_height_0__pin_33_
+ sb_2__8_/left_bottom_grid_pin_34_ sb_1__8_/right_bottom_grid_pin_34_ sb_2__8_/left_bottom_grid_pin_35_
+ sb_1__8_/right_bottom_grid_pin_35_ sb_2__8_/left_bottom_grid_pin_36_ sb_1__8_/right_bottom_grid_pin_36_
+ sb_2__8_/left_bottom_grid_pin_37_ sb_1__8_/right_bottom_grid_pin_37_ sb_2__8_/left_bottom_grid_pin_38_
+ sb_1__8_/right_bottom_grid_pin_38_ sb_2__8_/left_bottom_grid_pin_39_ sb_1__8_/right_bottom_grid_pin_39_
+ cbx_2__8_/bottom_grid_pin_3_ sb_2__8_/left_bottom_grid_pin_40_ sb_1__8_/right_bottom_grid_pin_40_
+ sb_2__8_/left_bottom_grid_pin_41_ sb_1__8_/right_bottom_grid_pin_41_ cbx_2__8_/bottom_grid_pin_4_
+ cbx_2__8_/bottom_grid_pin_5_ cbx_2__8_/bottom_grid_pin_6_ cbx_2__8_/bottom_grid_pin_7_
+ cbx_2__8_/bottom_grid_pin_8_ cbx_2__8_/bottom_grid_pin_9_ grid_clb
Xsb_7__5_ sb_7__5_/Test_en_N_out sb_7__5_/Test_en_S_in VGND VPWR sb_7__5_/bottom_left_grid_pin_42_
+ sb_7__5_/bottom_left_grid_pin_43_ sb_7__5_/bottom_left_grid_pin_44_ sb_7__5_/bottom_left_grid_pin_45_
+ sb_7__5_/bottom_left_grid_pin_46_ sb_7__5_/bottom_left_grid_pin_47_ sb_7__5_/bottom_left_grid_pin_48_
+ sb_7__5_/bottom_left_grid_pin_49_ sb_7__5_/ccff_head sb_7__5_/ccff_tail sb_7__5_/chanx_left_in[0]
+ sb_7__5_/chanx_left_in[10] sb_7__5_/chanx_left_in[11] sb_7__5_/chanx_left_in[12]
+ sb_7__5_/chanx_left_in[13] sb_7__5_/chanx_left_in[14] sb_7__5_/chanx_left_in[15]
+ sb_7__5_/chanx_left_in[16] sb_7__5_/chanx_left_in[17] sb_7__5_/chanx_left_in[18]
+ sb_7__5_/chanx_left_in[19] sb_7__5_/chanx_left_in[1] sb_7__5_/chanx_left_in[2] sb_7__5_/chanx_left_in[3]
+ sb_7__5_/chanx_left_in[4] sb_7__5_/chanx_left_in[5] sb_7__5_/chanx_left_in[6] sb_7__5_/chanx_left_in[7]
+ sb_7__5_/chanx_left_in[8] sb_7__5_/chanx_left_in[9] sb_7__5_/chanx_left_out[0] sb_7__5_/chanx_left_out[10]
+ sb_7__5_/chanx_left_out[11] sb_7__5_/chanx_left_out[12] sb_7__5_/chanx_left_out[13]
+ sb_7__5_/chanx_left_out[14] sb_7__5_/chanx_left_out[15] sb_7__5_/chanx_left_out[16]
+ sb_7__5_/chanx_left_out[17] sb_7__5_/chanx_left_out[18] sb_7__5_/chanx_left_out[19]
+ sb_7__5_/chanx_left_out[1] sb_7__5_/chanx_left_out[2] sb_7__5_/chanx_left_out[3]
+ sb_7__5_/chanx_left_out[4] sb_7__5_/chanx_left_out[5] sb_7__5_/chanx_left_out[6]
+ sb_7__5_/chanx_left_out[7] sb_7__5_/chanx_left_out[8] sb_7__5_/chanx_left_out[9]
+ sb_7__5_/chanx_right_in[0] sb_7__5_/chanx_right_in[10] sb_7__5_/chanx_right_in[11]
+ sb_7__5_/chanx_right_in[12] sb_7__5_/chanx_right_in[13] sb_7__5_/chanx_right_in[14]
+ sb_7__5_/chanx_right_in[15] sb_7__5_/chanx_right_in[16] sb_7__5_/chanx_right_in[17]
+ sb_7__5_/chanx_right_in[18] sb_7__5_/chanx_right_in[19] sb_7__5_/chanx_right_in[1]
+ sb_7__5_/chanx_right_in[2] sb_7__5_/chanx_right_in[3] sb_7__5_/chanx_right_in[4]
+ sb_7__5_/chanx_right_in[5] sb_7__5_/chanx_right_in[6] sb_7__5_/chanx_right_in[7]
+ sb_7__5_/chanx_right_in[8] sb_7__5_/chanx_right_in[9] cbx_8__5_/chanx_left_in[0]
+ cbx_8__5_/chanx_left_in[10] cbx_8__5_/chanx_left_in[11] cbx_8__5_/chanx_left_in[12]
+ cbx_8__5_/chanx_left_in[13] cbx_8__5_/chanx_left_in[14] cbx_8__5_/chanx_left_in[15]
+ cbx_8__5_/chanx_left_in[16] cbx_8__5_/chanx_left_in[17] cbx_8__5_/chanx_left_in[18]
+ cbx_8__5_/chanx_left_in[19] cbx_8__5_/chanx_left_in[1] cbx_8__5_/chanx_left_in[2]
+ cbx_8__5_/chanx_left_in[3] cbx_8__5_/chanx_left_in[4] cbx_8__5_/chanx_left_in[5]
+ cbx_8__5_/chanx_left_in[6] cbx_8__5_/chanx_left_in[7] cbx_8__5_/chanx_left_in[8]
+ cbx_8__5_/chanx_left_in[9] cby_7__5_/chany_top_out[0] cby_7__5_/chany_top_out[10]
+ cby_7__5_/chany_top_out[11] cby_7__5_/chany_top_out[12] cby_7__5_/chany_top_out[13]
+ cby_7__5_/chany_top_out[14] cby_7__5_/chany_top_out[15] cby_7__5_/chany_top_out[16]
+ cby_7__5_/chany_top_out[17] cby_7__5_/chany_top_out[18] cby_7__5_/chany_top_out[19]
+ cby_7__5_/chany_top_out[1] cby_7__5_/chany_top_out[2] cby_7__5_/chany_top_out[3]
+ cby_7__5_/chany_top_out[4] cby_7__5_/chany_top_out[5] cby_7__5_/chany_top_out[6]
+ cby_7__5_/chany_top_out[7] cby_7__5_/chany_top_out[8] cby_7__5_/chany_top_out[9]
+ cby_7__5_/chany_top_in[0] cby_7__5_/chany_top_in[10] cby_7__5_/chany_top_in[11]
+ cby_7__5_/chany_top_in[12] cby_7__5_/chany_top_in[13] cby_7__5_/chany_top_in[14]
+ cby_7__5_/chany_top_in[15] cby_7__5_/chany_top_in[16] cby_7__5_/chany_top_in[17]
+ cby_7__5_/chany_top_in[18] cby_7__5_/chany_top_in[19] cby_7__5_/chany_top_in[1]
+ cby_7__5_/chany_top_in[2] cby_7__5_/chany_top_in[3] cby_7__5_/chany_top_in[4] cby_7__5_/chany_top_in[5]
+ cby_7__5_/chany_top_in[6] cby_7__5_/chany_top_in[7] cby_7__5_/chany_top_in[8] cby_7__5_/chany_top_in[9]
+ sb_7__5_/chany_top_in[0] sb_7__5_/chany_top_in[10] sb_7__5_/chany_top_in[11] sb_7__5_/chany_top_in[12]
+ sb_7__5_/chany_top_in[13] sb_7__5_/chany_top_in[14] sb_7__5_/chany_top_in[15] sb_7__5_/chany_top_in[16]
+ sb_7__5_/chany_top_in[17] sb_7__5_/chany_top_in[18] sb_7__5_/chany_top_in[19] sb_7__5_/chany_top_in[1]
+ sb_7__5_/chany_top_in[2] sb_7__5_/chany_top_in[3] sb_7__5_/chany_top_in[4] sb_7__5_/chany_top_in[5]
+ sb_7__5_/chany_top_in[6] sb_7__5_/chany_top_in[7] sb_7__5_/chany_top_in[8] sb_7__5_/chany_top_in[9]
+ sb_7__5_/chany_top_out[0] sb_7__5_/chany_top_out[10] sb_7__5_/chany_top_out[11]
+ sb_7__5_/chany_top_out[12] sb_7__5_/chany_top_out[13] sb_7__5_/chany_top_out[14]
+ sb_7__5_/chany_top_out[15] sb_7__5_/chany_top_out[16] sb_7__5_/chany_top_out[17]
+ sb_7__5_/chany_top_out[18] sb_7__5_/chany_top_out[19] sb_7__5_/chany_top_out[1]
+ sb_7__5_/chany_top_out[2] sb_7__5_/chany_top_out[3] sb_7__5_/chany_top_out[4] sb_7__5_/chany_top_out[5]
+ sb_7__5_/chany_top_out[6] sb_7__5_/chany_top_out[7] sb_7__5_/chany_top_out[8] sb_7__5_/chany_top_out[9]
+ sb_7__5_/clk_1_E_out sb_7__5_/clk_1_N_in sb_7__5_/clk_1_W_out sb_7__5_/clk_2_E_out
+ sb_7__5_/clk_2_N_in sb_7__5_/clk_2_N_out sb_7__5_/clk_2_S_out sb_7__5_/clk_2_W_out
+ sb_7__5_/clk_3_E_out sb_7__5_/clk_3_N_in sb_7__5_/clk_3_N_out sb_7__5_/clk_3_S_out
+ sb_7__5_/clk_3_W_out sb_7__5_/left_bottom_grid_pin_34_ sb_7__5_/left_bottom_grid_pin_35_
+ sb_7__5_/left_bottom_grid_pin_36_ sb_7__5_/left_bottom_grid_pin_37_ sb_7__5_/left_bottom_grid_pin_38_
+ sb_7__5_/left_bottom_grid_pin_39_ sb_7__5_/left_bottom_grid_pin_40_ sb_7__5_/left_bottom_grid_pin_41_
+ sb_7__5_/prog_clk_0_N_in sb_7__5_/prog_clk_1_E_out sb_7__5_/prog_clk_1_N_in sb_7__5_/prog_clk_1_W_out
+ sb_7__5_/prog_clk_2_E_out sb_7__5_/prog_clk_2_N_in sb_7__5_/prog_clk_2_N_out sb_7__5_/prog_clk_2_S_out
+ sb_7__5_/prog_clk_2_W_out sb_7__5_/prog_clk_3_E_out sb_7__5_/prog_clk_3_N_in sb_7__5_/prog_clk_3_N_out
+ sb_7__5_/prog_clk_3_S_out sb_7__5_/prog_clk_3_W_out sb_7__5_/right_bottom_grid_pin_34_
+ sb_7__5_/right_bottom_grid_pin_35_ sb_7__5_/right_bottom_grid_pin_36_ sb_7__5_/right_bottom_grid_pin_37_
+ sb_7__5_/right_bottom_grid_pin_38_ sb_7__5_/right_bottom_grid_pin_39_ sb_7__5_/right_bottom_grid_pin_40_
+ sb_7__5_/right_bottom_grid_pin_41_ sb_7__5_/top_left_grid_pin_42_ sb_7__5_/top_left_grid_pin_43_
+ sb_7__5_/top_left_grid_pin_44_ sb_7__5_/top_left_grid_pin_45_ sb_7__5_/top_left_grid_pin_46_
+ sb_7__5_/top_left_grid_pin_47_ sb_7__5_/top_left_grid_pin_48_ sb_7__5_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_4__2_ sb_4__2_/Test_en_N_out sb_4__2_/Test_en_S_in VGND VPWR sb_4__2_/bottom_left_grid_pin_42_
+ sb_4__2_/bottom_left_grid_pin_43_ sb_4__2_/bottom_left_grid_pin_44_ sb_4__2_/bottom_left_grid_pin_45_
+ sb_4__2_/bottom_left_grid_pin_46_ sb_4__2_/bottom_left_grid_pin_47_ sb_4__2_/bottom_left_grid_pin_48_
+ sb_4__2_/bottom_left_grid_pin_49_ sb_4__2_/ccff_head sb_4__2_/ccff_tail sb_4__2_/chanx_left_in[0]
+ sb_4__2_/chanx_left_in[10] sb_4__2_/chanx_left_in[11] sb_4__2_/chanx_left_in[12]
+ sb_4__2_/chanx_left_in[13] sb_4__2_/chanx_left_in[14] sb_4__2_/chanx_left_in[15]
+ sb_4__2_/chanx_left_in[16] sb_4__2_/chanx_left_in[17] sb_4__2_/chanx_left_in[18]
+ sb_4__2_/chanx_left_in[19] sb_4__2_/chanx_left_in[1] sb_4__2_/chanx_left_in[2] sb_4__2_/chanx_left_in[3]
+ sb_4__2_/chanx_left_in[4] sb_4__2_/chanx_left_in[5] sb_4__2_/chanx_left_in[6] sb_4__2_/chanx_left_in[7]
+ sb_4__2_/chanx_left_in[8] sb_4__2_/chanx_left_in[9] sb_4__2_/chanx_left_out[0] sb_4__2_/chanx_left_out[10]
+ sb_4__2_/chanx_left_out[11] sb_4__2_/chanx_left_out[12] sb_4__2_/chanx_left_out[13]
+ sb_4__2_/chanx_left_out[14] sb_4__2_/chanx_left_out[15] sb_4__2_/chanx_left_out[16]
+ sb_4__2_/chanx_left_out[17] sb_4__2_/chanx_left_out[18] sb_4__2_/chanx_left_out[19]
+ sb_4__2_/chanx_left_out[1] sb_4__2_/chanx_left_out[2] sb_4__2_/chanx_left_out[3]
+ sb_4__2_/chanx_left_out[4] sb_4__2_/chanx_left_out[5] sb_4__2_/chanx_left_out[6]
+ sb_4__2_/chanx_left_out[7] sb_4__2_/chanx_left_out[8] sb_4__2_/chanx_left_out[9]
+ sb_4__2_/chanx_right_in[0] sb_4__2_/chanx_right_in[10] sb_4__2_/chanx_right_in[11]
+ sb_4__2_/chanx_right_in[12] sb_4__2_/chanx_right_in[13] sb_4__2_/chanx_right_in[14]
+ sb_4__2_/chanx_right_in[15] sb_4__2_/chanx_right_in[16] sb_4__2_/chanx_right_in[17]
+ sb_4__2_/chanx_right_in[18] sb_4__2_/chanx_right_in[19] sb_4__2_/chanx_right_in[1]
+ sb_4__2_/chanx_right_in[2] sb_4__2_/chanx_right_in[3] sb_4__2_/chanx_right_in[4]
+ sb_4__2_/chanx_right_in[5] sb_4__2_/chanx_right_in[6] sb_4__2_/chanx_right_in[7]
+ sb_4__2_/chanx_right_in[8] sb_4__2_/chanx_right_in[9] cbx_5__2_/chanx_left_in[0]
+ cbx_5__2_/chanx_left_in[10] cbx_5__2_/chanx_left_in[11] cbx_5__2_/chanx_left_in[12]
+ cbx_5__2_/chanx_left_in[13] cbx_5__2_/chanx_left_in[14] cbx_5__2_/chanx_left_in[15]
+ cbx_5__2_/chanx_left_in[16] cbx_5__2_/chanx_left_in[17] cbx_5__2_/chanx_left_in[18]
+ cbx_5__2_/chanx_left_in[19] cbx_5__2_/chanx_left_in[1] cbx_5__2_/chanx_left_in[2]
+ cbx_5__2_/chanx_left_in[3] cbx_5__2_/chanx_left_in[4] cbx_5__2_/chanx_left_in[5]
+ cbx_5__2_/chanx_left_in[6] cbx_5__2_/chanx_left_in[7] cbx_5__2_/chanx_left_in[8]
+ cbx_5__2_/chanx_left_in[9] cby_4__2_/chany_top_out[0] cby_4__2_/chany_top_out[10]
+ cby_4__2_/chany_top_out[11] cby_4__2_/chany_top_out[12] cby_4__2_/chany_top_out[13]
+ cby_4__2_/chany_top_out[14] cby_4__2_/chany_top_out[15] cby_4__2_/chany_top_out[16]
+ cby_4__2_/chany_top_out[17] cby_4__2_/chany_top_out[18] cby_4__2_/chany_top_out[19]
+ cby_4__2_/chany_top_out[1] cby_4__2_/chany_top_out[2] cby_4__2_/chany_top_out[3]
+ cby_4__2_/chany_top_out[4] cby_4__2_/chany_top_out[5] cby_4__2_/chany_top_out[6]
+ cby_4__2_/chany_top_out[7] cby_4__2_/chany_top_out[8] cby_4__2_/chany_top_out[9]
+ cby_4__2_/chany_top_in[0] cby_4__2_/chany_top_in[10] cby_4__2_/chany_top_in[11]
+ cby_4__2_/chany_top_in[12] cby_4__2_/chany_top_in[13] cby_4__2_/chany_top_in[14]
+ cby_4__2_/chany_top_in[15] cby_4__2_/chany_top_in[16] cby_4__2_/chany_top_in[17]
+ cby_4__2_/chany_top_in[18] cby_4__2_/chany_top_in[19] cby_4__2_/chany_top_in[1]
+ cby_4__2_/chany_top_in[2] cby_4__2_/chany_top_in[3] cby_4__2_/chany_top_in[4] cby_4__2_/chany_top_in[5]
+ cby_4__2_/chany_top_in[6] cby_4__2_/chany_top_in[7] cby_4__2_/chany_top_in[8] cby_4__2_/chany_top_in[9]
+ sb_4__2_/chany_top_in[0] sb_4__2_/chany_top_in[10] sb_4__2_/chany_top_in[11] sb_4__2_/chany_top_in[12]
+ sb_4__2_/chany_top_in[13] sb_4__2_/chany_top_in[14] sb_4__2_/chany_top_in[15] sb_4__2_/chany_top_in[16]
+ sb_4__2_/chany_top_in[17] sb_4__2_/chany_top_in[18] sb_4__2_/chany_top_in[19] sb_4__2_/chany_top_in[1]
+ sb_4__2_/chany_top_in[2] sb_4__2_/chany_top_in[3] sb_4__2_/chany_top_in[4] sb_4__2_/chany_top_in[5]
+ sb_4__2_/chany_top_in[6] sb_4__2_/chany_top_in[7] sb_4__2_/chany_top_in[8] sb_4__2_/chany_top_in[9]
+ sb_4__2_/chany_top_out[0] sb_4__2_/chany_top_out[10] sb_4__2_/chany_top_out[11]
+ sb_4__2_/chany_top_out[12] sb_4__2_/chany_top_out[13] sb_4__2_/chany_top_out[14]
+ sb_4__2_/chany_top_out[15] sb_4__2_/chany_top_out[16] sb_4__2_/chany_top_out[17]
+ sb_4__2_/chany_top_out[18] sb_4__2_/chany_top_out[19] sb_4__2_/chany_top_out[1]
+ sb_4__2_/chany_top_out[2] sb_4__2_/chany_top_out[3] sb_4__2_/chany_top_out[4] sb_4__2_/chany_top_out[5]
+ sb_4__2_/chany_top_out[6] sb_4__2_/chany_top_out[7] sb_4__2_/chany_top_out[8] sb_4__2_/chany_top_out[9]
+ sb_4__2_/clk_1_E_out sb_4__2_/clk_1_N_in sb_4__2_/clk_1_W_out sb_4__2_/clk_2_E_out
+ sb_4__2_/clk_2_N_in sb_4__2_/clk_2_N_out sb_4__2_/clk_2_S_out sb_4__2_/clk_2_W_out
+ sb_4__2_/clk_3_E_out sb_4__2_/clk_3_N_in sb_4__2_/clk_3_N_out sb_4__2_/clk_3_S_out
+ sb_4__2_/clk_3_W_out sb_4__2_/left_bottom_grid_pin_34_ sb_4__2_/left_bottom_grid_pin_35_
+ sb_4__2_/left_bottom_grid_pin_36_ sb_4__2_/left_bottom_grid_pin_37_ sb_4__2_/left_bottom_grid_pin_38_
+ sb_4__2_/left_bottom_grid_pin_39_ sb_4__2_/left_bottom_grid_pin_40_ sb_4__2_/left_bottom_grid_pin_41_
+ sb_4__2_/prog_clk_0_N_in sb_4__2_/prog_clk_1_E_out sb_4__2_/prog_clk_1_N_in sb_4__2_/prog_clk_1_W_out
+ sb_4__2_/prog_clk_2_E_out sb_4__2_/prog_clk_2_N_in sb_4__2_/prog_clk_2_N_out sb_4__2_/prog_clk_2_S_out
+ sb_4__2_/prog_clk_2_W_out sb_4__2_/prog_clk_3_E_out sb_4__2_/prog_clk_3_N_in sb_4__2_/prog_clk_3_N_out
+ sb_4__2_/prog_clk_3_S_out sb_4__2_/prog_clk_3_W_out sb_4__2_/right_bottom_grid_pin_34_
+ sb_4__2_/right_bottom_grid_pin_35_ sb_4__2_/right_bottom_grid_pin_36_ sb_4__2_/right_bottom_grid_pin_37_
+ sb_4__2_/right_bottom_grid_pin_38_ sb_4__2_/right_bottom_grid_pin_39_ sb_4__2_/right_bottom_grid_pin_40_
+ sb_4__2_/right_bottom_grid_pin_41_ sb_4__2_/top_left_grid_pin_42_ sb_4__2_/top_left_grid_pin_43_
+ sb_4__2_/top_left_grid_pin_44_ sb_4__2_/top_left_grid_pin_45_ sb_4__2_/top_left_grid_pin_46_
+ sb_4__2_/top_left_grid_pin_47_ sb_4__2_/top_left_grid_pin_48_ sb_4__2_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_3__6_ cby_3__6_/Test_en_W_in cby_3__6_/Test_en_E_out cby_3__6_/Test_en_N_out
+ cby_3__6_/Test_en_W_in cby_3__6_/Test_en_W_in cby_3__6_/Test_en_W_out VGND VPWR
+ cby_3__6_/ccff_head cby_3__6_/ccff_tail sb_3__5_/chany_top_out[0] sb_3__5_/chany_top_out[10]
+ sb_3__5_/chany_top_out[11] sb_3__5_/chany_top_out[12] sb_3__5_/chany_top_out[13]
+ sb_3__5_/chany_top_out[14] sb_3__5_/chany_top_out[15] sb_3__5_/chany_top_out[16]
+ sb_3__5_/chany_top_out[17] sb_3__5_/chany_top_out[18] sb_3__5_/chany_top_out[19]
+ sb_3__5_/chany_top_out[1] sb_3__5_/chany_top_out[2] sb_3__5_/chany_top_out[3] sb_3__5_/chany_top_out[4]
+ sb_3__5_/chany_top_out[5] sb_3__5_/chany_top_out[6] sb_3__5_/chany_top_out[7] sb_3__5_/chany_top_out[8]
+ sb_3__5_/chany_top_out[9] sb_3__5_/chany_top_in[0] sb_3__5_/chany_top_in[10] sb_3__5_/chany_top_in[11]
+ sb_3__5_/chany_top_in[12] sb_3__5_/chany_top_in[13] sb_3__5_/chany_top_in[14] sb_3__5_/chany_top_in[15]
+ sb_3__5_/chany_top_in[16] sb_3__5_/chany_top_in[17] sb_3__5_/chany_top_in[18] sb_3__5_/chany_top_in[19]
+ sb_3__5_/chany_top_in[1] sb_3__5_/chany_top_in[2] sb_3__5_/chany_top_in[3] sb_3__5_/chany_top_in[4]
+ sb_3__5_/chany_top_in[5] sb_3__5_/chany_top_in[6] sb_3__5_/chany_top_in[7] sb_3__5_/chany_top_in[8]
+ sb_3__5_/chany_top_in[9] cby_3__6_/chany_top_in[0] cby_3__6_/chany_top_in[10] cby_3__6_/chany_top_in[11]
+ cby_3__6_/chany_top_in[12] cby_3__6_/chany_top_in[13] cby_3__6_/chany_top_in[14]
+ cby_3__6_/chany_top_in[15] cby_3__6_/chany_top_in[16] cby_3__6_/chany_top_in[17]
+ cby_3__6_/chany_top_in[18] cby_3__6_/chany_top_in[19] cby_3__6_/chany_top_in[1]
+ cby_3__6_/chany_top_in[2] cby_3__6_/chany_top_in[3] cby_3__6_/chany_top_in[4] cby_3__6_/chany_top_in[5]
+ cby_3__6_/chany_top_in[6] cby_3__6_/chany_top_in[7] cby_3__6_/chany_top_in[8] cby_3__6_/chany_top_in[9]
+ cby_3__6_/chany_top_out[0] cby_3__6_/chany_top_out[10] cby_3__6_/chany_top_out[11]
+ cby_3__6_/chany_top_out[12] cby_3__6_/chany_top_out[13] cby_3__6_/chany_top_out[14]
+ cby_3__6_/chany_top_out[15] cby_3__6_/chany_top_out[16] cby_3__6_/chany_top_out[17]
+ cby_3__6_/chany_top_out[18] cby_3__6_/chany_top_out[19] cby_3__6_/chany_top_out[1]
+ cby_3__6_/chany_top_out[2] cby_3__6_/chany_top_out[3] cby_3__6_/chany_top_out[4]
+ cby_3__6_/chany_top_out[5] cby_3__6_/chany_top_out[6] cby_3__6_/chany_top_out[7]
+ cby_3__6_/chany_top_out[8] cby_3__6_/chany_top_out[9] cby_3__6_/clk_2_N_out sb_3__6_/clk_2_S_out
+ sb_3__5_/clk_1_N_in cby_3__6_/clk_3_N_out cby_3__6_/clk_3_S_in cby_3__6_/clk_3_S_out
+ cby_3__6_/left_grid_pin_16_ cby_3__6_/left_grid_pin_17_ cby_3__6_/left_grid_pin_18_
+ cby_3__6_/left_grid_pin_19_ cby_3__6_/left_grid_pin_20_ cby_3__6_/left_grid_pin_21_
+ cby_3__6_/left_grid_pin_22_ cby_3__6_/left_grid_pin_23_ cby_3__6_/left_grid_pin_24_
+ cby_3__6_/left_grid_pin_25_ cby_3__6_/left_grid_pin_26_ cby_3__6_/left_grid_pin_27_
+ cby_3__6_/left_grid_pin_28_ cby_3__6_/left_grid_pin_29_ cby_3__6_/left_grid_pin_30_
+ cby_3__6_/left_grid_pin_31_ cby_3__6_/prog_clk_0_N_out sb_3__5_/prog_clk_0_N_in
+ cby_3__6_/prog_clk_0_W_in cby_3__6_/prog_clk_2_N_out sb_3__6_/prog_clk_2_S_out sb_3__5_/prog_clk_1_N_in
+ cby_3__6_/prog_clk_3_N_out cby_3__6_/prog_clk_3_S_in cby_3__6_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_3__7_ cbx_3__7_/REGIN_FEEDTHROUGH cbx_3__7_/REGOUT_FEEDTHROUGH cbx_3__7_/SC_IN_BOT
+ cbx_3__7_/SC_IN_TOP cbx_3__7_/SC_OUT_BOT cbx_3__7_/SC_OUT_TOP VGND VPWR cbx_3__7_/bottom_grid_pin_0_
+ cbx_3__7_/bottom_grid_pin_10_ cbx_3__7_/bottom_grid_pin_11_ cbx_3__7_/bottom_grid_pin_12_
+ cbx_3__7_/bottom_grid_pin_13_ cbx_3__7_/bottom_grid_pin_14_ cbx_3__7_/bottom_grid_pin_15_
+ cbx_3__7_/bottom_grid_pin_1_ cbx_3__7_/bottom_grid_pin_2_ cbx_3__7_/bottom_grid_pin_3_
+ cbx_3__7_/bottom_grid_pin_4_ cbx_3__7_/bottom_grid_pin_5_ cbx_3__7_/bottom_grid_pin_6_
+ cbx_3__7_/bottom_grid_pin_7_ cbx_3__7_/bottom_grid_pin_8_ cbx_3__7_/bottom_grid_pin_9_
+ sb_3__7_/ccff_tail sb_2__7_/ccff_head cbx_3__7_/chanx_left_in[0] cbx_3__7_/chanx_left_in[10]
+ cbx_3__7_/chanx_left_in[11] cbx_3__7_/chanx_left_in[12] cbx_3__7_/chanx_left_in[13]
+ cbx_3__7_/chanx_left_in[14] cbx_3__7_/chanx_left_in[15] cbx_3__7_/chanx_left_in[16]
+ cbx_3__7_/chanx_left_in[17] cbx_3__7_/chanx_left_in[18] cbx_3__7_/chanx_left_in[19]
+ cbx_3__7_/chanx_left_in[1] cbx_3__7_/chanx_left_in[2] cbx_3__7_/chanx_left_in[3]
+ cbx_3__7_/chanx_left_in[4] cbx_3__7_/chanx_left_in[5] cbx_3__7_/chanx_left_in[6]
+ cbx_3__7_/chanx_left_in[7] cbx_3__7_/chanx_left_in[8] cbx_3__7_/chanx_left_in[9]
+ sb_2__7_/chanx_right_in[0] sb_2__7_/chanx_right_in[10] sb_2__7_/chanx_right_in[11]
+ sb_2__7_/chanx_right_in[12] sb_2__7_/chanx_right_in[13] sb_2__7_/chanx_right_in[14]
+ sb_2__7_/chanx_right_in[15] sb_2__7_/chanx_right_in[16] sb_2__7_/chanx_right_in[17]
+ sb_2__7_/chanx_right_in[18] sb_2__7_/chanx_right_in[19] sb_2__7_/chanx_right_in[1]
+ sb_2__7_/chanx_right_in[2] sb_2__7_/chanx_right_in[3] sb_2__7_/chanx_right_in[4]
+ sb_2__7_/chanx_right_in[5] sb_2__7_/chanx_right_in[6] sb_2__7_/chanx_right_in[7]
+ sb_2__7_/chanx_right_in[8] sb_2__7_/chanx_right_in[9] sb_3__7_/chanx_left_out[0]
+ sb_3__7_/chanx_left_out[10] sb_3__7_/chanx_left_out[11] sb_3__7_/chanx_left_out[12]
+ sb_3__7_/chanx_left_out[13] sb_3__7_/chanx_left_out[14] sb_3__7_/chanx_left_out[15]
+ sb_3__7_/chanx_left_out[16] sb_3__7_/chanx_left_out[17] sb_3__7_/chanx_left_out[18]
+ sb_3__7_/chanx_left_out[19] sb_3__7_/chanx_left_out[1] sb_3__7_/chanx_left_out[2]
+ sb_3__7_/chanx_left_out[3] sb_3__7_/chanx_left_out[4] sb_3__7_/chanx_left_out[5]
+ sb_3__7_/chanx_left_out[6] sb_3__7_/chanx_left_out[7] sb_3__7_/chanx_left_out[8]
+ sb_3__7_/chanx_left_out[9] sb_3__7_/chanx_left_in[0] sb_3__7_/chanx_left_in[10]
+ sb_3__7_/chanx_left_in[11] sb_3__7_/chanx_left_in[12] sb_3__7_/chanx_left_in[13]
+ sb_3__7_/chanx_left_in[14] sb_3__7_/chanx_left_in[15] sb_3__7_/chanx_left_in[16]
+ sb_3__7_/chanx_left_in[17] sb_3__7_/chanx_left_in[18] sb_3__7_/chanx_left_in[19]
+ sb_3__7_/chanx_left_in[1] sb_3__7_/chanx_left_in[2] sb_3__7_/chanx_left_in[3] sb_3__7_/chanx_left_in[4]
+ sb_3__7_/chanx_left_in[5] sb_3__7_/chanx_left_in[6] sb_3__7_/chanx_left_in[7] sb_3__7_/chanx_left_in[8]
+ sb_3__7_/chanx_left_in[9] cbx_3__7_/clk_1_N_out cbx_3__7_/clk_1_S_out sb_3__7_/clk_1_W_out
+ cbx_3__7_/clk_2_E_out cbx_3__7_/clk_2_W_in cbx_3__7_/clk_2_W_out cbx_3__7_/clk_3_E_out
+ cbx_3__7_/clk_3_W_in cbx_3__7_/clk_3_W_out cbx_3__7_/prog_clk_0_N_in cbx_3__7_/prog_clk_0_W_out
+ cbx_3__7_/prog_clk_1_N_out cbx_3__7_/prog_clk_1_S_out sb_3__7_/prog_clk_1_W_out
+ cbx_3__7_/prog_clk_2_E_out cbx_3__7_/prog_clk_2_W_in cbx_3__7_/prog_clk_2_W_out
+ cbx_3__7_/prog_clk_3_E_out cbx_3__7_/prog_clk_3_W_in cbx_3__7_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_7__4_ sb_7__4_/Test_en_N_out sb_7__4_/Test_en_S_in VGND VPWR sb_7__4_/bottom_left_grid_pin_42_
+ sb_7__4_/bottom_left_grid_pin_43_ sb_7__4_/bottom_left_grid_pin_44_ sb_7__4_/bottom_left_grid_pin_45_
+ sb_7__4_/bottom_left_grid_pin_46_ sb_7__4_/bottom_left_grid_pin_47_ sb_7__4_/bottom_left_grid_pin_48_
+ sb_7__4_/bottom_left_grid_pin_49_ sb_7__4_/ccff_head sb_7__4_/ccff_tail sb_7__4_/chanx_left_in[0]
+ sb_7__4_/chanx_left_in[10] sb_7__4_/chanx_left_in[11] sb_7__4_/chanx_left_in[12]
+ sb_7__4_/chanx_left_in[13] sb_7__4_/chanx_left_in[14] sb_7__4_/chanx_left_in[15]
+ sb_7__4_/chanx_left_in[16] sb_7__4_/chanx_left_in[17] sb_7__4_/chanx_left_in[18]
+ sb_7__4_/chanx_left_in[19] sb_7__4_/chanx_left_in[1] sb_7__4_/chanx_left_in[2] sb_7__4_/chanx_left_in[3]
+ sb_7__4_/chanx_left_in[4] sb_7__4_/chanx_left_in[5] sb_7__4_/chanx_left_in[6] sb_7__4_/chanx_left_in[7]
+ sb_7__4_/chanx_left_in[8] sb_7__4_/chanx_left_in[9] sb_7__4_/chanx_left_out[0] sb_7__4_/chanx_left_out[10]
+ sb_7__4_/chanx_left_out[11] sb_7__4_/chanx_left_out[12] sb_7__4_/chanx_left_out[13]
+ sb_7__4_/chanx_left_out[14] sb_7__4_/chanx_left_out[15] sb_7__4_/chanx_left_out[16]
+ sb_7__4_/chanx_left_out[17] sb_7__4_/chanx_left_out[18] sb_7__4_/chanx_left_out[19]
+ sb_7__4_/chanx_left_out[1] sb_7__4_/chanx_left_out[2] sb_7__4_/chanx_left_out[3]
+ sb_7__4_/chanx_left_out[4] sb_7__4_/chanx_left_out[5] sb_7__4_/chanx_left_out[6]
+ sb_7__4_/chanx_left_out[7] sb_7__4_/chanx_left_out[8] sb_7__4_/chanx_left_out[9]
+ sb_7__4_/chanx_right_in[0] sb_7__4_/chanx_right_in[10] sb_7__4_/chanx_right_in[11]
+ sb_7__4_/chanx_right_in[12] sb_7__4_/chanx_right_in[13] sb_7__4_/chanx_right_in[14]
+ sb_7__4_/chanx_right_in[15] sb_7__4_/chanx_right_in[16] sb_7__4_/chanx_right_in[17]
+ sb_7__4_/chanx_right_in[18] sb_7__4_/chanx_right_in[19] sb_7__4_/chanx_right_in[1]
+ sb_7__4_/chanx_right_in[2] sb_7__4_/chanx_right_in[3] sb_7__4_/chanx_right_in[4]
+ sb_7__4_/chanx_right_in[5] sb_7__4_/chanx_right_in[6] sb_7__4_/chanx_right_in[7]
+ sb_7__4_/chanx_right_in[8] sb_7__4_/chanx_right_in[9] cbx_8__4_/chanx_left_in[0]
+ cbx_8__4_/chanx_left_in[10] cbx_8__4_/chanx_left_in[11] cbx_8__4_/chanx_left_in[12]
+ cbx_8__4_/chanx_left_in[13] cbx_8__4_/chanx_left_in[14] cbx_8__4_/chanx_left_in[15]
+ cbx_8__4_/chanx_left_in[16] cbx_8__4_/chanx_left_in[17] cbx_8__4_/chanx_left_in[18]
+ cbx_8__4_/chanx_left_in[19] cbx_8__4_/chanx_left_in[1] cbx_8__4_/chanx_left_in[2]
+ cbx_8__4_/chanx_left_in[3] cbx_8__4_/chanx_left_in[4] cbx_8__4_/chanx_left_in[5]
+ cbx_8__4_/chanx_left_in[6] cbx_8__4_/chanx_left_in[7] cbx_8__4_/chanx_left_in[8]
+ cbx_8__4_/chanx_left_in[9] cby_7__4_/chany_top_out[0] cby_7__4_/chany_top_out[10]
+ cby_7__4_/chany_top_out[11] cby_7__4_/chany_top_out[12] cby_7__4_/chany_top_out[13]
+ cby_7__4_/chany_top_out[14] cby_7__4_/chany_top_out[15] cby_7__4_/chany_top_out[16]
+ cby_7__4_/chany_top_out[17] cby_7__4_/chany_top_out[18] cby_7__4_/chany_top_out[19]
+ cby_7__4_/chany_top_out[1] cby_7__4_/chany_top_out[2] cby_7__4_/chany_top_out[3]
+ cby_7__4_/chany_top_out[4] cby_7__4_/chany_top_out[5] cby_7__4_/chany_top_out[6]
+ cby_7__4_/chany_top_out[7] cby_7__4_/chany_top_out[8] cby_7__4_/chany_top_out[9]
+ cby_7__4_/chany_top_in[0] cby_7__4_/chany_top_in[10] cby_7__4_/chany_top_in[11]
+ cby_7__4_/chany_top_in[12] cby_7__4_/chany_top_in[13] cby_7__4_/chany_top_in[14]
+ cby_7__4_/chany_top_in[15] cby_7__4_/chany_top_in[16] cby_7__4_/chany_top_in[17]
+ cby_7__4_/chany_top_in[18] cby_7__4_/chany_top_in[19] cby_7__4_/chany_top_in[1]
+ cby_7__4_/chany_top_in[2] cby_7__4_/chany_top_in[3] cby_7__4_/chany_top_in[4] cby_7__4_/chany_top_in[5]
+ cby_7__4_/chany_top_in[6] cby_7__4_/chany_top_in[7] cby_7__4_/chany_top_in[8] cby_7__4_/chany_top_in[9]
+ sb_7__4_/chany_top_in[0] sb_7__4_/chany_top_in[10] sb_7__4_/chany_top_in[11] sb_7__4_/chany_top_in[12]
+ sb_7__4_/chany_top_in[13] sb_7__4_/chany_top_in[14] sb_7__4_/chany_top_in[15] sb_7__4_/chany_top_in[16]
+ sb_7__4_/chany_top_in[17] sb_7__4_/chany_top_in[18] sb_7__4_/chany_top_in[19] sb_7__4_/chany_top_in[1]
+ sb_7__4_/chany_top_in[2] sb_7__4_/chany_top_in[3] sb_7__4_/chany_top_in[4] sb_7__4_/chany_top_in[5]
+ sb_7__4_/chany_top_in[6] sb_7__4_/chany_top_in[7] sb_7__4_/chany_top_in[8] sb_7__4_/chany_top_in[9]
+ sb_7__4_/chany_top_out[0] sb_7__4_/chany_top_out[10] sb_7__4_/chany_top_out[11]
+ sb_7__4_/chany_top_out[12] sb_7__4_/chany_top_out[13] sb_7__4_/chany_top_out[14]
+ sb_7__4_/chany_top_out[15] sb_7__4_/chany_top_out[16] sb_7__4_/chany_top_out[17]
+ sb_7__4_/chany_top_out[18] sb_7__4_/chany_top_out[19] sb_7__4_/chany_top_out[1]
+ sb_7__4_/chany_top_out[2] sb_7__4_/chany_top_out[3] sb_7__4_/chany_top_out[4] sb_7__4_/chany_top_out[5]
+ sb_7__4_/chany_top_out[6] sb_7__4_/chany_top_out[7] sb_7__4_/chany_top_out[8] sb_7__4_/chany_top_out[9]
+ sb_7__4_/clk_1_E_out sb_7__4_/clk_1_N_in sb_7__4_/clk_1_W_out sb_7__4_/clk_2_E_out
+ sb_7__4_/clk_2_N_in sb_7__4_/clk_2_N_out sb_7__4_/clk_2_S_out sb_7__4_/clk_2_W_out
+ sb_7__4_/clk_3_E_out sb_7__4_/clk_3_N_in sb_7__4_/clk_3_N_out sb_7__4_/clk_3_S_out
+ sb_7__4_/clk_3_W_out sb_7__4_/left_bottom_grid_pin_34_ sb_7__4_/left_bottom_grid_pin_35_
+ sb_7__4_/left_bottom_grid_pin_36_ sb_7__4_/left_bottom_grid_pin_37_ sb_7__4_/left_bottom_grid_pin_38_
+ sb_7__4_/left_bottom_grid_pin_39_ sb_7__4_/left_bottom_grid_pin_40_ sb_7__4_/left_bottom_grid_pin_41_
+ sb_7__4_/prog_clk_0_N_in sb_7__4_/prog_clk_1_E_out sb_7__4_/prog_clk_1_N_in sb_7__4_/prog_clk_1_W_out
+ sb_7__4_/prog_clk_2_E_out sb_7__4_/prog_clk_2_N_in sb_7__4_/prog_clk_2_N_out sb_7__4_/prog_clk_2_S_out
+ sb_7__4_/prog_clk_2_W_out sb_7__4_/prog_clk_3_E_out sb_7__4_/prog_clk_3_N_in sb_7__4_/prog_clk_3_N_out
+ sb_7__4_/prog_clk_3_S_out sb_7__4_/prog_clk_3_W_out sb_7__4_/right_bottom_grid_pin_34_
+ sb_7__4_/right_bottom_grid_pin_35_ sb_7__4_/right_bottom_grid_pin_36_ sb_7__4_/right_bottom_grid_pin_37_
+ sb_7__4_/right_bottom_grid_pin_38_ sb_7__4_/right_bottom_grid_pin_39_ sb_7__4_/right_bottom_grid_pin_40_
+ sb_7__4_/right_bottom_grid_pin_41_ sb_7__4_/top_left_grid_pin_42_ sb_7__4_/top_left_grid_pin_43_
+ sb_7__4_/top_left_grid_pin_44_ sb_7__4_/top_left_grid_pin_45_ sb_7__4_/top_left_grid_pin_46_
+ sb_7__4_/top_left_grid_pin_47_ sb_7__4_/top_left_grid_pin_48_ sb_7__4_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_0__3_ IO_ISOL_N VGND VPWR sb_0__3_/ccff_tail cby_0__3_/ccff_tail sb_0__2_/chany_top_out[0]
+ sb_0__2_/chany_top_out[10] sb_0__2_/chany_top_out[11] sb_0__2_/chany_top_out[12]
+ sb_0__2_/chany_top_out[13] sb_0__2_/chany_top_out[14] sb_0__2_/chany_top_out[15]
+ sb_0__2_/chany_top_out[16] sb_0__2_/chany_top_out[17] sb_0__2_/chany_top_out[18]
+ sb_0__2_/chany_top_out[19] sb_0__2_/chany_top_out[1] sb_0__2_/chany_top_out[2] sb_0__2_/chany_top_out[3]
+ sb_0__2_/chany_top_out[4] sb_0__2_/chany_top_out[5] sb_0__2_/chany_top_out[6] sb_0__2_/chany_top_out[7]
+ sb_0__2_/chany_top_out[8] sb_0__2_/chany_top_out[9] sb_0__2_/chany_top_in[0] sb_0__2_/chany_top_in[10]
+ sb_0__2_/chany_top_in[11] sb_0__2_/chany_top_in[12] sb_0__2_/chany_top_in[13] sb_0__2_/chany_top_in[14]
+ sb_0__2_/chany_top_in[15] sb_0__2_/chany_top_in[16] sb_0__2_/chany_top_in[17] sb_0__2_/chany_top_in[18]
+ sb_0__2_/chany_top_in[19] sb_0__2_/chany_top_in[1] sb_0__2_/chany_top_in[2] sb_0__2_/chany_top_in[3]
+ sb_0__2_/chany_top_in[4] sb_0__2_/chany_top_in[5] sb_0__2_/chany_top_in[6] sb_0__2_/chany_top_in[7]
+ sb_0__2_/chany_top_in[8] sb_0__2_/chany_top_in[9] cby_0__3_/chany_top_in[0] cby_0__3_/chany_top_in[10]
+ cby_0__3_/chany_top_in[11] cby_0__3_/chany_top_in[12] cby_0__3_/chany_top_in[13]
+ cby_0__3_/chany_top_in[14] cby_0__3_/chany_top_in[15] cby_0__3_/chany_top_in[16]
+ cby_0__3_/chany_top_in[17] cby_0__3_/chany_top_in[18] cby_0__3_/chany_top_in[19]
+ cby_0__3_/chany_top_in[1] cby_0__3_/chany_top_in[2] cby_0__3_/chany_top_in[3] cby_0__3_/chany_top_in[4]
+ cby_0__3_/chany_top_in[5] cby_0__3_/chany_top_in[6] cby_0__3_/chany_top_in[7] cby_0__3_/chany_top_in[8]
+ cby_0__3_/chany_top_in[9] cby_0__3_/chany_top_out[0] cby_0__3_/chany_top_out[10]
+ cby_0__3_/chany_top_out[11] cby_0__3_/chany_top_out[12] cby_0__3_/chany_top_out[13]
+ cby_0__3_/chany_top_out[14] cby_0__3_/chany_top_out[15] cby_0__3_/chany_top_out[16]
+ cby_0__3_/chany_top_out[17] cby_0__3_/chany_top_out[18] cby_0__3_/chany_top_out[19]
+ cby_0__3_/chany_top_out[1] cby_0__3_/chany_top_out[2] cby_0__3_/chany_top_out[3]
+ cby_0__3_/chany_top_out[4] cby_0__3_/chany_top_out[5] cby_0__3_/chany_top_out[6]
+ cby_0__3_/chany_top_out[7] cby_0__3_/chany_top_out[8] cby_0__3_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
+ cby_0__3_/left_grid_pin_0_ cby_0__3_/prog_clk_0_E_in cby_0__3_/left_grid_pin_0_
+ sb_0__2_/top_left_grid_pin_1_ sb_0__3_/bottom_left_grid_pin_1_ cby_0__1_
Xgrid_clb_2__7_ cbx_2__6_/SC_OUT_TOP grid_clb_2__7_/SC_OUT_BOT cbx_2__7_/SC_IN_BOT
+ cby_2__7_/Test_en_W_out grid_clb_2__7_/Test_en_E_out cby_2__7_/Test_en_W_out cby_1__7_/Test_en_W_in
+ VGND VPWR cbx_2__6_/REGIN_FEEDTHROUGH grid_clb_2__7_/bottom_width_0_height_0__pin_51_
+ cby_1__7_/ccff_tail cby_2__7_/ccff_head cbx_2__7_/clk_1_S_out cbx_2__7_/clk_1_S_out
+ cby_2__7_/prog_clk_0_W_in cbx_2__7_/prog_clk_1_S_out grid_clb_2__7_/prog_clk_0_N_out
+ cbx_2__7_/prog_clk_1_S_out cbx_2__6_/prog_clk_0_N_in grid_clb_2__7_/prog_clk_0_W_out
+ cby_2__7_/left_grid_pin_16_ cby_2__7_/left_grid_pin_17_ cby_2__7_/left_grid_pin_18_
+ cby_2__7_/left_grid_pin_19_ cby_2__7_/left_grid_pin_20_ cby_2__7_/left_grid_pin_21_
+ cby_2__7_/left_grid_pin_22_ cby_2__7_/left_grid_pin_23_ cby_2__7_/left_grid_pin_24_
+ cby_2__7_/left_grid_pin_25_ cby_2__7_/left_grid_pin_26_ cby_2__7_/left_grid_pin_27_
+ cby_2__7_/left_grid_pin_28_ cby_2__7_/left_grid_pin_29_ cby_2__7_/left_grid_pin_30_
+ cby_2__7_/left_grid_pin_31_ sb_2__6_/top_left_grid_pin_42_ sb_2__7_/bottom_left_grid_pin_42_
+ sb_2__6_/top_left_grid_pin_43_ sb_2__7_/bottom_left_grid_pin_43_ sb_2__6_/top_left_grid_pin_44_
+ sb_2__7_/bottom_left_grid_pin_44_ sb_2__6_/top_left_grid_pin_45_ sb_2__7_/bottom_left_grid_pin_45_
+ sb_2__6_/top_left_grid_pin_46_ sb_2__7_/bottom_left_grid_pin_46_ sb_2__6_/top_left_grid_pin_47_
+ sb_2__7_/bottom_left_grid_pin_47_ sb_2__6_/top_left_grid_pin_48_ sb_2__7_/bottom_left_grid_pin_48_
+ sb_2__6_/top_left_grid_pin_49_ sb_2__7_/bottom_left_grid_pin_49_ cbx_2__7_/bottom_grid_pin_0_
+ cbx_2__7_/bottom_grid_pin_10_ cbx_2__7_/bottom_grid_pin_11_ cbx_2__7_/bottom_grid_pin_12_
+ cbx_2__7_/bottom_grid_pin_13_ cbx_2__7_/bottom_grid_pin_14_ cbx_2__7_/bottom_grid_pin_15_
+ cbx_2__7_/bottom_grid_pin_1_ cbx_2__7_/bottom_grid_pin_2_ cbx_2__7_/REGOUT_FEEDTHROUGH
+ grid_clb_2__7_/top_width_0_height_0__pin_33_ sb_2__7_/left_bottom_grid_pin_34_ sb_1__7_/right_bottom_grid_pin_34_
+ sb_2__7_/left_bottom_grid_pin_35_ sb_1__7_/right_bottom_grid_pin_35_ sb_2__7_/left_bottom_grid_pin_36_
+ sb_1__7_/right_bottom_grid_pin_36_ sb_2__7_/left_bottom_grid_pin_37_ sb_1__7_/right_bottom_grid_pin_37_
+ sb_2__7_/left_bottom_grid_pin_38_ sb_1__7_/right_bottom_grid_pin_38_ sb_2__7_/left_bottom_grid_pin_39_
+ sb_1__7_/right_bottom_grid_pin_39_ cbx_2__7_/bottom_grid_pin_3_ sb_2__7_/left_bottom_grid_pin_40_
+ sb_1__7_/right_bottom_grid_pin_40_ sb_2__7_/left_bottom_grid_pin_41_ sb_1__7_/right_bottom_grid_pin_41_
+ cbx_2__7_/bottom_grid_pin_4_ cbx_2__7_/bottom_grid_pin_5_ cbx_2__7_/bottom_grid_pin_6_
+ cbx_2__7_/bottom_grid_pin_7_ cbx_2__7_/bottom_grid_pin_8_ cbx_2__7_/bottom_grid_pin_9_
+ grid_clb
Xsb_4__1_ sb_4__1_/Test_en_N_out sb_4__1_/Test_en_S_in VGND VPWR sb_4__1_/bottom_left_grid_pin_42_
+ sb_4__1_/bottom_left_grid_pin_43_ sb_4__1_/bottom_left_grid_pin_44_ sb_4__1_/bottom_left_grid_pin_45_
+ sb_4__1_/bottom_left_grid_pin_46_ sb_4__1_/bottom_left_grid_pin_47_ sb_4__1_/bottom_left_grid_pin_48_
+ sb_4__1_/bottom_left_grid_pin_49_ sb_4__1_/ccff_head sb_4__1_/ccff_tail sb_4__1_/chanx_left_in[0]
+ sb_4__1_/chanx_left_in[10] sb_4__1_/chanx_left_in[11] sb_4__1_/chanx_left_in[12]
+ sb_4__1_/chanx_left_in[13] sb_4__1_/chanx_left_in[14] sb_4__1_/chanx_left_in[15]
+ sb_4__1_/chanx_left_in[16] sb_4__1_/chanx_left_in[17] sb_4__1_/chanx_left_in[18]
+ sb_4__1_/chanx_left_in[19] sb_4__1_/chanx_left_in[1] sb_4__1_/chanx_left_in[2] sb_4__1_/chanx_left_in[3]
+ sb_4__1_/chanx_left_in[4] sb_4__1_/chanx_left_in[5] sb_4__1_/chanx_left_in[6] sb_4__1_/chanx_left_in[7]
+ sb_4__1_/chanx_left_in[8] sb_4__1_/chanx_left_in[9] sb_4__1_/chanx_left_out[0] sb_4__1_/chanx_left_out[10]
+ sb_4__1_/chanx_left_out[11] sb_4__1_/chanx_left_out[12] sb_4__1_/chanx_left_out[13]
+ sb_4__1_/chanx_left_out[14] sb_4__1_/chanx_left_out[15] sb_4__1_/chanx_left_out[16]
+ sb_4__1_/chanx_left_out[17] sb_4__1_/chanx_left_out[18] sb_4__1_/chanx_left_out[19]
+ sb_4__1_/chanx_left_out[1] sb_4__1_/chanx_left_out[2] sb_4__1_/chanx_left_out[3]
+ sb_4__1_/chanx_left_out[4] sb_4__1_/chanx_left_out[5] sb_4__1_/chanx_left_out[6]
+ sb_4__1_/chanx_left_out[7] sb_4__1_/chanx_left_out[8] sb_4__1_/chanx_left_out[9]
+ sb_4__1_/chanx_right_in[0] sb_4__1_/chanx_right_in[10] sb_4__1_/chanx_right_in[11]
+ sb_4__1_/chanx_right_in[12] sb_4__1_/chanx_right_in[13] sb_4__1_/chanx_right_in[14]
+ sb_4__1_/chanx_right_in[15] sb_4__1_/chanx_right_in[16] sb_4__1_/chanx_right_in[17]
+ sb_4__1_/chanx_right_in[18] sb_4__1_/chanx_right_in[19] sb_4__1_/chanx_right_in[1]
+ sb_4__1_/chanx_right_in[2] sb_4__1_/chanx_right_in[3] sb_4__1_/chanx_right_in[4]
+ sb_4__1_/chanx_right_in[5] sb_4__1_/chanx_right_in[6] sb_4__1_/chanx_right_in[7]
+ sb_4__1_/chanx_right_in[8] sb_4__1_/chanx_right_in[9] cbx_5__1_/chanx_left_in[0]
+ cbx_5__1_/chanx_left_in[10] cbx_5__1_/chanx_left_in[11] cbx_5__1_/chanx_left_in[12]
+ cbx_5__1_/chanx_left_in[13] cbx_5__1_/chanx_left_in[14] cbx_5__1_/chanx_left_in[15]
+ cbx_5__1_/chanx_left_in[16] cbx_5__1_/chanx_left_in[17] cbx_5__1_/chanx_left_in[18]
+ cbx_5__1_/chanx_left_in[19] cbx_5__1_/chanx_left_in[1] cbx_5__1_/chanx_left_in[2]
+ cbx_5__1_/chanx_left_in[3] cbx_5__1_/chanx_left_in[4] cbx_5__1_/chanx_left_in[5]
+ cbx_5__1_/chanx_left_in[6] cbx_5__1_/chanx_left_in[7] cbx_5__1_/chanx_left_in[8]
+ cbx_5__1_/chanx_left_in[9] cby_4__1_/chany_top_out[0] cby_4__1_/chany_top_out[10]
+ cby_4__1_/chany_top_out[11] cby_4__1_/chany_top_out[12] cby_4__1_/chany_top_out[13]
+ cby_4__1_/chany_top_out[14] cby_4__1_/chany_top_out[15] cby_4__1_/chany_top_out[16]
+ cby_4__1_/chany_top_out[17] cby_4__1_/chany_top_out[18] cby_4__1_/chany_top_out[19]
+ cby_4__1_/chany_top_out[1] cby_4__1_/chany_top_out[2] cby_4__1_/chany_top_out[3]
+ cby_4__1_/chany_top_out[4] cby_4__1_/chany_top_out[5] cby_4__1_/chany_top_out[6]
+ cby_4__1_/chany_top_out[7] cby_4__1_/chany_top_out[8] cby_4__1_/chany_top_out[9]
+ cby_4__1_/chany_top_in[0] cby_4__1_/chany_top_in[10] cby_4__1_/chany_top_in[11]
+ cby_4__1_/chany_top_in[12] cby_4__1_/chany_top_in[13] cby_4__1_/chany_top_in[14]
+ cby_4__1_/chany_top_in[15] cby_4__1_/chany_top_in[16] cby_4__1_/chany_top_in[17]
+ cby_4__1_/chany_top_in[18] cby_4__1_/chany_top_in[19] cby_4__1_/chany_top_in[1]
+ cby_4__1_/chany_top_in[2] cby_4__1_/chany_top_in[3] cby_4__1_/chany_top_in[4] cby_4__1_/chany_top_in[5]
+ cby_4__1_/chany_top_in[6] cby_4__1_/chany_top_in[7] cby_4__1_/chany_top_in[8] cby_4__1_/chany_top_in[9]
+ sb_4__1_/chany_top_in[0] sb_4__1_/chany_top_in[10] sb_4__1_/chany_top_in[11] sb_4__1_/chany_top_in[12]
+ sb_4__1_/chany_top_in[13] sb_4__1_/chany_top_in[14] sb_4__1_/chany_top_in[15] sb_4__1_/chany_top_in[16]
+ sb_4__1_/chany_top_in[17] sb_4__1_/chany_top_in[18] sb_4__1_/chany_top_in[19] sb_4__1_/chany_top_in[1]
+ sb_4__1_/chany_top_in[2] sb_4__1_/chany_top_in[3] sb_4__1_/chany_top_in[4] sb_4__1_/chany_top_in[5]
+ sb_4__1_/chany_top_in[6] sb_4__1_/chany_top_in[7] sb_4__1_/chany_top_in[8] sb_4__1_/chany_top_in[9]
+ sb_4__1_/chany_top_out[0] sb_4__1_/chany_top_out[10] sb_4__1_/chany_top_out[11]
+ sb_4__1_/chany_top_out[12] sb_4__1_/chany_top_out[13] sb_4__1_/chany_top_out[14]
+ sb_4__1_/chany_top_out[15] sb_4__1_/chany_top_out[16] sb_4__1_/chany_top_out[17]
+ sb_4__1_/chany_top_out[18] sb_4__1_/chany_top_out[19] sb_4__1_/chany_top_out[1]
+ sb_4__1_/chany_top_out[2] sb_4__1_/chany_top_out[3] sb_4__1_/chany_top_out[4] sb_4__1_/chany_top_out[5]
+ sb_4__1_/chany_top_out[6] sb_4__1_/chany_top_out[7] sb_4__1_/chany_top_out[8] sb_4__1_/chany_top_out[9]
+ sb_4__1_/clk_1_E_out sb_4__1_/clk_1_N_in sb_4__1_/clk_1_W_out sb_4__1_/clk_2_E_out
+ sb_4__1_/clk_2_N_in sb_4__1_/clk_2_N_out sb_4__1_/clk_2_S_out sb_4__1_/clk_2_W_out
+ sb_4__1_/clk_3_E_out sb_4__1_/clk_3_N_in sb_4__1_/clk_3_N_out sb_4__1_/clk_3_S_out
+ sb_4__1_/clk_3_W_out sb_4__1_/left_bottom_grid_pin_34_ sb_4__1_/left_bottom_grid_pin_35_
+ sb_4__1_/left_bottom_grid_pin_36_ sb_4__1_/left_bottom_grid_pin_37_ sb_4__1_/left_bottom_grid_pin_38_
+ sb_4__1_/left_bottom_grid_pin_39_ sb_4__1_/left_bottom_grid_pin_40_ sb_4__1_/left_bottom_grid_pin_41_
+ sb_4__1_/prog_clk_0_N_in sb_4__1_/prog_clk_1_E_out sb_4__1_/prog_clk_1_N_in sb_4__1_/prog_clk_1_W_out
+ sb_4__1_/prog_clk_2_E_out sb_4__1_/prog_clk_2_N_in sb_4__1_/prog_clk_2_N_out sb_4__1_/prog_clk_2_S_out
+ sb_4__1_/prog_clk_2_W_out sb_4__1_/prog_clk_3_E_out sb_4__1_/prog_clk_3_N_in sb_4__1_/prog_clk_3_N_out
+ sb_4__1_/prog_clk_3_S_out sb_4__1_/prog_clk_3_W_out sb_4__1_/right_bottom_grid_pin_34_
+ sb_4__1_/right_bottom_grid_pin_35_ sb_4__1_/right_bottom_grid_pin_36_ sb_4__1_/right_bottom_grid_pin_37_
+ sb_4__1_/right_bottom_grid_pin_38_ sb_4__1_/right_bottom_grid_pin_39_ sb_4__1_/right_bottom_grid_pin_40_
+ sb_4__1_/right_bottom_grid_pin_41_ sb_4__1_/top_left_grid_pin_42_ sb_4__1_/top_left_grid_pin_43_
+ sb_4__1_/top_left_grid_pin_44_ sb_4__1_/top_left_grid_pin_45_ sb_4__1_/top_left_grid_pin_46_
+ sb_4__1_/top_left_grid_pin_47_ sb_4__1_/top_left_grid_pin_48_ sb_4__1_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_6__8_ cby_6__8_/Test_en_W_in cby_6__8_/Test_en_E_out cby_6__8_/Test_en_N_out
+ cby_6__8_/Test_en_W_in cby_6__8_/Test_en_W_in cby_6__8_/Test_en_W_out VGND VPWR
+ cby_6__8_/ccff_head cby_6__8_/ccff_tail sb_6__7_/chany_top_out[0] sb_6__7_/chany_top_out[10]
+ sb_6__7_/chany_top_out[11] sb_6__7_/chany_top_out[12] sb_6__7_/chany_top_out[13]
+ sb_6__7_/chany_top_out[14] sb_6__7_/chany_top_out[15] sb_6__7_/chany_top_out[16]
+ sb_6__7_/chany_top_out[17] sb_6__7_/chany_top_out[18] sb_6__7_/chany_top_out[19]
+ sb_6__7_/chany_top_out[1] sb_6__7_/chany_top_out[2] sb_6__7_/chany_top_out[3] sb_6__7_/chany_top_out[4]
+ sb_6__7_/chany_top_out[5] sb_6__7_/chany_top_out[6] sb_6__7_/chany_top_out[7] sb_6__7_/chany_top_out[8]
+ sb_6__7_/chany_top_out[9] sb_6__7_/chany_top_in[0] sb_6__7_/chany_top_in[10] sb_6__7_/chany_top_in[11]
+ sb_6__7_/chany_top_in[12] sb_6__7_/chany_top_in[13] sb_6__7_/chany_top_in[14] sb_6__7_/chany_top_in[15]
+ sb_6__7_/chany_top_in[16] sb_6__7_/chany_top_in[17] sb_6__7_/chany_top_in[18] sb_6__7_/chany_top_in[19]
+ sb_6__7_/chany_top_in[1] sb_6__7_/chany_top_in[2] sb_6__7_/chany_top_in[3] sb_6__7_/chany_top_in[4]
+ sb_6__7_/chany_top_in[5] sb_6__7_/chany_top_in[6] sb_6__7_/chany_top_in[7] sb_6__7_/chany_top_in[8]
+ sb_6__7_/chany_top_in[9] cby_6__8_/chany_top_in[0] cby_6__8_/chany_top_in[10] cby_6__8_/chany_top_in[11]
+ cby_6__8_/chany_top_in[12] cby_6__8_/chany_top_in[13] cby_6__8_/chany_top_in[14]
+ cby_6__8_/chany_top_in[15] cby_6__8_/chany_top_in[16] cby_6__8_/chany_top_in[17]
+ cby_6__8_/chany_top_in[18] cby_6__8_/chany_top_in[19] cby_6__8_/chany_top_in[1]
+ cby_6__8_/chany_top_in[2] cby_6__8_/chany_top_in[3] cby_6__8_/chany_top_in[4] cby_6__8_/chany_top_in[5]
+ cby_6__8_/chany_top_in[6] cby_6__8_/chany_top_in[7] cby_6__8_/chany_top_in[8] cby_6__8_/chany_top_in[9]
+ cby_6__8_/chany_top_out[0] cby_6__8_/chany_top_out[10] cby_6__8_/chany_top_out[11]
+ cby_6__8_/chany_top_out[12] cby_6__8_/chany_top_out[13] cby_6__8_/chany_top_out[14]
+ cby_6__8_/chany_top_out[15] cby_6__8_/chany_top_out[16] cby_6__8_/chany_top_out[17]
+ cby_6__8_/chany_top_out[18] cby_6__8_/chany_top_out[19] cby_6__8_/chany_top_out[1]
+ cby_6__8_/chany_top_out[2] cby_6__8_/chany_top_out[3] cby_6__8_/chany_top_out[4]
+ cby_6__8_/chany_top_out[5] cby_6__8_/chany_top_out[6] cby_6__8_/chany_top_out[7]
+ cby_6__8_/chany_top_out[8] cby_6__8_/chany_top_out[9] cby_6__8_/clk_2_N_out cby_6__8_/clk_2_S_in
+ cby_6__8_/clk_2_S_out cby_6__8_/clk_3_N_out cby_6__8_/clk_3_S_in cby_6__8_/clk_3_S_out
+ cby_6__8_/left_grid_pin_16_ cby_6__8_/left_grid_pin_17_ cby_6__8_/left_grid_pin_18_
+ cby_6__8_/left_grid_pin_19_ cby_6__8_/left_grid_pin_20_ cby_6__8_/left_grid_pin_21_
+ cby_6__8_/left_grid_pin_22_ cby_6__8_/left_grid_pin_23_ cby_6__8_/left_grid_pin_24_
+ cby_6__8_/left_grid_pin_25_ cby_6__8_/left_grid_pin_26_ cby_6__8_/left_grid_pin_27_
+ cby_6__8_/left_grid_pin_28_ cby_6__8_/left_grid_pin_29_ cby_6__8_/left_grid_pin_30_
+ cby_6__8_/left_grid_pin_31_ sb_6__8_/prog_clk_0_S_in sb_6__7_/prog_clk_0_N_in cby_6__8_/prog_clk_0_W_in
+ cby_6__8_/prog_clk_2_N_out cby_6__8_/prog_clk_2_S_in cby_6__8_/prog_clk_2_S_out
+ cby_6__8_/prog_clk_3_N_out cby_6__8_/prog_clk_3_S_in cby_6__8_/prog_clk_3_S_out
+ cby_1__1_
Xcby_3__5_ cby_3__5_/Test_en_W_in cby_3__5_/Test_en_E_out cby_3__5_/Test_en_N_out
+ cby_3__5_/Test_en_W_in cby_3__5_/Test_en_W_in cby_3__5_/Test_en_W_out VGND VPWR
+ cby_3__5_/ccff_head cby_3__5_/ccff_tail sb_3__4_/chany_top_out[0] sb_3__4_/chany_top_out[10]
+ sb_3__4_/chany_top_out[11] sb_3__4_/chany_top_out[12] sb_3__4_/chany_top_out[13]
+ sb_3__4_/chany_top_out[14] sb_3__4_/chany_top_out[15] sb_3__4_/chany_top_out[16]
+ sb_3__4_/chany_top_out[17] sb_3__4_/chany_top_out[18] sb_3__4_/chany_top_out[19]
+ sb_3__4_/chany_top_out[1] sb_3__4_/chany_top_out[2] sb_3__4_/chany_top_out[3] sb_3__4_/chany_top_out[4]
+ sb_3__4_/chany_top_out[5] sb_3__4_/chany_top_out[6] sb_3__4_/chany_top_out[7] sb_3__4_/chany_top_out[8]
+ sb_3__4_/chany_top_out[9] sb_3__4_/chany_top_in[0] sb_3__4_/chany_top_in[10] sb_3__4_/chany_top_in[11]
+ sb_3__4_/chany_top_in[12] sb_3__4_/chany_top_in[13] sb_3__4_/chany_top_in[14] sb_3__4_/chany_top_in[15]
+ sb_3__4_/chany_top_in[16] sb_3__4_/chany_top_in[17] sb_3__4_/chany_top_in[18] sb_3__4_/chany_top_in[19]
+ sb_3__4_/chany_top_in[1] sb_3__4_/chany_top_in[2] sb_3__4_/chany_top_in[3] sb_3__4_/chany_top_in[4]
+ sb_3__4_/chany_top_in[5] sb_3__4_/chany_top_in[6] sb_3__4_/chany_top_in[7] sb_3__4_/chany_top_in[8]
+ sb_3__4_/chany_top_in[9] cby_3__5_/chany_top_in[0] cby_3__5_/chany_top_in[10] cby_3__5_/chany_top_in[11]
+ cby_3__5_/chany_top_in[12] cby_3__5_/chany_top_in[13] cby_3__5_/chany_top_in[14]
+ cby_3__5_/chany_top_in[15] cby_3__5_/chany_top_in[16] cby_3__5_/chany_top_in[17]
+ cby_3__5_/chany_top_in[18] cby_3__5_/chany_top_in[19] cby_3__5_/chany_top_in[1]
+ cby_3__5_/chany_top_in[2] cby_3__5_/chany_top_in[3] cby_3__5_/chany_top_in[4] cby_3__5_/chany_top_in[5]
+ cby_3__5_/chany_top_in[6] cby_3__5_/chany_top_in[7] cby_3__5_/chany_top_in[8] cby_3__5_/chany_top_in[9]
+ cby_3__5_/chany_top_out[0] cby_3__5_/chany_top_out[10] cby_3__5_/chany_top_out[11]
+ cby_3__5_/chany_top_out[12] cby_3__5_/chany_top_out[13] cby_3__5_/chany_top_out[14]
+ cby_3__5_/chany_top_out[15] cby_3__5_/chany_top_out[16] cby_3__5_/chany_top_out[17]
+ cby_3__5_/chany_top_out[18] cby_3__5_/chany_top_out[19] cby_3__5_/chany_top_out[1]
+ cby_3__5_/chany_top_out[2] cby_3__5_/chany_top_out[3] cby_3__5_/chany_top_out[4]
+ cby_3__5_/chany_top_out[5] cby_3__5_/chany_top_out[6] cby_3__5_/chany_top_out[7]
+ cby_3__5_/chany_top_out[8] cby_3__5_/chany_top_out[9] cby_3__5_/clk_2_N_out cby_3__5_/clk_2_S_in
+ cby_3__5_/clk_2_S_out cby_3__5_/clk_3_N_out cby_3__5_/clk_3_S_in cby_3__5_/clk_3_S_out
+ cby_3__5_/left_grid_pin_16_ cby_3__5_/left_grid_pin_17_ cby_3__5_/left_grid_pin_18_
+ cby_3__5_/left_grid_pin_19_ cby_3__5_/left_grid_pin_20_ cby_3__5_/left_grid_pin_21_
+ cby_3__5_/left_grid_pin_22_ cby_3__5_/left_grid_pin_23_ cby_3__5_/left_grid_pin_24_
+ cby_3__5_/left_grid_pin_25_ cby_3__5_/left_grid_pin_26_ cby_3__5_/left_grid_pin_27_
+ cby_3__5_/left_grid_pin_28_ cby_3__5_/left_grid_pin_29_ cby_3__5_/left_grid_pin_30_
+ cby_3__5_/left_grid_pin_31_ cby_3__5_/prog_clk_0_N_out sb_3__4_/prog_clk_0_N_in
+ cby_3__5_/prog_clk_0_W_in cby_3__5_/prog_clk_2_N_out cby_3__5_/prog_clk_2_S_in cby_3__5_/prog_clk_2_S_out
+ cby_3__5_/prog_clk_3_N_out cby_3__5_/prog_clk_3_S_in cby_3__5_/prog_clk_3_S_out
+ cby_1__1_
Xcby_0__2_ IO_ISOL_N VGND VPWR sb_0__2_/ccff_tail cby_0__2_/ccff_tail sb_0__1_/chany_top_out[0]
+ sb_0__1_/chany_top_out[10] sb_0__1_/chany_top_out[11] sb_0__1_/chany_top_out[12]
+ sb_0__1_/chany_top_out[13] sb_0__1_/chany_top_out[14] sb_0__1_/chany_top_out[15]
+ sb_0__1_/chany_top_out[16] sb_0__1_/chany_top_out[17] sb_0__1_/chany_top_out[18]
+ sb_0__1_/chany_top_out[19] sb_0__1_/chany_top_out[1] sb_0__1_/chany_top_out[2] sb_0__1_/chany_top_out[3]
+ sb_0__1_/chany_top_out[4] sb_0__1_/chany_top_out[5] sb_0__1_/chany_top_out[6] sb_0__1_/chany_top_out[7]
+ sb_0__1_/chany_top_out[8] sb_0__1_/chany_top_out[9] sb_0__1_/chany_top_in[0] sb_0__1_/chany_top_in[10]
+ sb_0__1_/chany_top_in[11] sb_0__1_/chany_top_in[12] sb_0__1_/chany_top_in[13] sb_0__1_/chany_top_in[14]
+ sb_0__1_/chany_top_in[15] sb_0__1_/chany_top_in[16] sb_0__1_/chany_top_in[17] sb_0__1_/chany_top_in[18]
+ sb_0__1_/chany_top_in[19] sb_0__1_/chany_top_in[1] sb_0__1_/chany_top_in[2] sb_0__1_/chany_top_in[3]
+ sb_0__1_/chany_top_in[4] sb_0__1_/chany_top_in[5] sb_0__1_/chany_top_in[6] sb_0__1_/chany_top_in[7]
+ sb_0__1_/chany_top_in[8] sb_0__1_/chany_top_in[9] cby_0__2_/chany_top_in[0] cby_0__2_/chany_top_in[10]
+ cby_0__2_/chany_top_in[11] cby_0__2_/chany_top_in[12] cby_0__2_/chany_top_in[13]
+ cby_0__2_/chany_top_in[14] cby_0__2_/chany_top_in[15] cby_0__2_/chany_top_in[16]
+ cby_0__2_/chany_top_in[17] cby_0__2_/chany_top_in[18] cby_0__2_/chany_top_in[19]
+ cby_0__2_/chany_top_in[1] cby_0__2_/chany_top_in[2] cby_0__2_/chany_top_in[3] cby_0__2_/chany_top_in[4]
+ cby_0__2_/chany_top_in[5] cby_0__2_/chany_top_in[6] cby_0__2_/chany_top_in[7] cby_0__2_/chany_top_in[8]
+ cby_0__2_/chany_top_in[9] cby_0__2_/chany_top_out[0] cby_0__2_/chany_top_out[10]
+ cby_0__2_/chany_top_out[11] cby_0__2_/chany_top_out[12] cby_0__2_/chany_top_out[13]
+ cby_0__2_/chany_top_out[14] cby_0__2_/chany_top_out[15] cby_0__2_/chany_top_out[16]
+ cby_0__2_/chany_top_out[17] cby_0__2_/chany_top_out[18] cby_0__2_/chany_top_out[19]
+ cby_0__2_/chany_top_out[1] cby_0__2_/chany_top_out[2] cby_0__2_/chany_top_out[3]
+ cby_0__2_/chany_top_out[4] cby_0__2_/chany_top_out[5] cby_0__2_/chany_top_out[6]
+ cby_0__2_/chany_top_out[7] cby_0__2_/chany_top_out[8] cby_0__2_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
+ cby_0__2_/left_grid_pin_0_ cby_0__2_/prog_clk_0_E_in cby_0__2_/left_grid_pin_0_
+ sb_0__1_/top_left_grid_pin_1_ sb_0__2_/bottom_left_grid_pin_1_ cby_0__1_
Xcbx_3__6_ cbx_3__6_/REGIN_FEEDTHROUGH cbx_3__6_/REGOUT_FEEDTHROUGH cbx_3__6_/SC_IN_BOT
+ cbx_3__6_/SC_IN_TOP cbx_3__6_/SC_OUT_BOT cbx_3__6_/SC_OUT_TOP VGND VPWR cbx_3__6_/bottom_grid_pin_0_
+ cbx_3__6_/bottom_grid_pin_10_ cbx_3__6_/bottom_grid_pin_11_ cbx_3__6_/bottom_grid_pin_12_
+ cbx_3__6_/bottom_grid_pin_13_ cbx_3__6_/bottom_grid_pin_14_ cbx_3__6_/bottom_grid_pin_15_
+ cbx_3__6_/bottom_grid_pin_1_ cbx_3__6_/bottom_grid_pin_2_ cbx_3__6_/bottom_grid_pin_3_
+ cbx_3__6_/bottom_grid_pin_4_ cbx_3__6_/bottom_grid_pin_5_ cbx_3__6_/bottom_grid_pin_6_
+ cbx_3__6_/bottom_grid_pin_7_ cbx_3__6_/bottom_grid_pin_8_ cbx_3__6_/bottom_grid_pin_9_
+ sb_3__6_/ccff_tail sb_2__6_/ccff_head cbx_3__6_/chanx_left_in[0] cbx_3__6_/chanx_left_in[10]
+ cbx_3__6_/chanx_left_in[11] cbx_3__6_/chanx_left_in[12] cbx_3__6_/chanx_left_in[13]
+ cbx_3__6_/chanx_left_in[14] cbx_3__6_/chanx_left_in[15] cbx_3__6_/chanx_left_in[16]
+ cbx_3__6_/chanx_left_in[17] cbx_3__6_/chanx_left_in[18] cbx_3__6_/chanx_left_in[19]
+ cbx_3__6_/chanx_left_in[1] cbx_3__6_/chanx_left_in[2] cbx_3__6_/chanx_left_in[3]
+ cbx_3__6_/chanx_left_in[4] cbx_3__6_/chanx_left_in[5] cbx_3__6_/chanx_left_in[6]
+ cbx_3__6_/chanx_left_in[7] cbx_3__6_/chanx_left_in[8] cbx_3__6_/chanx_left_in[9]
+ sb_2__6_/chanx_right_in[0] sb_2__6_/chanx_right_in[10] sb_2__6_/chanx_right_in[11]
+ sb_2__6_/chanx_right_in[12] sb_2__6_/chanx_right_in[13] sb_2__6_/chanx_right_in[14]
+ sb_2__6_/chanx_right_in[15] sb_2__6_/chanx_right_in[16] sb_2__6_/chanx_right_in[17]
+ sb_2__6_/chanx_right_in[18] sb_2__6_/chanx_right_in[19] sb_2__6_/chanx_right_in[1]
+ sb_2__6_/chanx_right_in[2] sb_2__6_/chanx_right_in[3] sb_2__6_/chanx_right_in[4]
+ sb_2__6_/chanx_right_in[5] sb_2__6_/chanx_right_in[6] sb_2__6_/chanx_right_in[7]
+ sb_2__6_/chanx_right_in[8] sb_2__6_/chanx_right_in[9] sb_3__6_/chanx_left_out[0]
+ sb_3__6_/chanx_left_out[10] sb_3__6_/chanx_left_out[11] sb_3__6_/chanx_left_out[12]
+ sb_3__6_/chanx_left_out[13] sb_3__6_/chanx_left_out[14] sb_3__6_/chanx_left_out[15]
+ sb_3__6_/chanx_left_out[16] sb_3__6_/chanx_left_out[17] sb_3__6_/chanx_left_out[18]
+ sb_3__6_/chanx_left_out[19] sb_3__6_/chanx_left_out[1] sb_3__6_/chanx_left_out[2]
+ sb_3__6_/chanx_left_out[3] sb_3__6_/chanx_left_out[4] sb_3__6_/chanx_left_out[5]
+ sb_3__6_/chanx_left_out[6] sb_3__6_/chanx_left_out[7] sb_3__6_/chanx_left_out[8]
+ sb_3__6_/chanx_left_out[9] sb_3__6_/chanx_left_in[0] sb_3__6_/chanx_left_in[10]
+ sb_3__6_/chanx_left_in[11] sb_3__6_/chanx_left_in[12] sb_3__6_/chanx_left_in[13]
+ sb_3__6_/chanx_left_in[14] sb_3__6_/chanx_left_in[15] sb_3__6_/chanx_left_in[16]
+ sb_3__6_/chanx_left_in[17] sb_3__6_/chanx_left_in[18] sb_3__6_/chanx_left_in[19]
+ sb_3__6_/chanx_left_in[1] sb_3__6_/chanx_left_in[2] sb_3__6_/chanx_left_in[3] sb_3__6_/chanx_left_in[4]
+ sb_3__6_/chanx_left_in[5] sb_3__6_/chanx_left_in[6] sb_3__6_/chanx_left_in[7] sb_3__6_/chanx_left_in[8]
+ sb_3__6_/chanx_left_in[9] cbx_3__6_/clk_1_N_out cbx_3__6_/clk_1_S_out cbx_3__6_/clk_1_W_in
+ sb_3__6_/clk_2_N_in sb_2__6_/clk_2_E_out cbx_3__6_/clk_2_W_out cbx_3__6_/clk_3_E_out
+ cbx_3__6_/clk_3_W_in cbx_3__6_/clk_3_W_out cbx_3__6_/prog_clk_0_N_in cbx_3__6_/prog_clk_0_W_out
+ cbx_3__6_/prog_clk_1_N_out cbx_3__6_/prog_clk_1_S_out cbx_3__6_/prog_clk_1_W_in
+ sb_3__6_/prog_clk_2_N_in sb_2__6_/prog_clk_2_E_out cbx_3__6_/prog_clk_2_W_out cbx_3__6_/prog_clk_3_E_out
+ cbx_3__6_/prog_clk_3_W_in cbx_3__6_/prog_clk_3_W_out cbx_1__1_
Xgrid_clb_2__6_ cbx_2__5_/SC_OUT_TOP grid_clb_2__6_/SC_OUT_BOT cbx_2__6_/SC_IN_BOT
+ cby_2__6_/Test_en_W_out grid_clb_2__6_/Test_en_E_out cby_2__6_/Test_en_W_out cby_1__6_/Test_en_W_in
+ VGND VPWR cbx_2__5_/REGIN_FEEDTHROUGH grid_clb_2__6_/bottom_width_0_height_0__pin_51_
+ cby_1__6_/ccff_tail cby_2__6_/ccff_head cbx_2__5_/clk_1_N_out cbx_2__5_/clk_1_N_out
+ cby_2__6_/prog_clk_0_W_in cbx_2__5_/prog_clk_1_N_out grid_clb_2__6_/prog_clk_0_N_out
+ cbx_2__5_/prog_clk_1_N_out cbx_2__5_/prog_clk_0_N_in grid_clb_2__6_/prog_clk_0_W_out
+ cby_2__6_/left_grid_pin_16_ cby_2__6_/left_grid_pin_17_ cby_2__6_/left_grid_pin_18_
+ cby_2__6_/left_grid_pin_19_ cby_2__6_/left_grid_pin_20_ cby_2__6_/left_grid_pin_21_
+ cby_2__6_/left_grid_pin_22_ cby_2__6_/left_grid_pin_23_ cby_2__6_/left_grid_pin_24_
+ cby_2__6_/left_grid_pin_25_ cby_2__6_/left_grid_pin_26_ cby_2__6_/left_grid_pin_27_
+ cby_2__6_/left_grid_pin_28_ cby_2__6_/left_grid_pin_29_ cby_2__6_/left_grid_pin_30_
+ cby_2__6_/left_grid_pin_31_ sb_2__5_/top_left_grid_pin_42_ sb_2__6_/bottom_left_grid_pin_42_
+ sb_2__5_/top_left_grid_pin_43_ sb_2__6_/bottom_left_grid_pin_43_ sb_2__5_/top_left_grid_pin_44_
+ sb_2__6_/bottom_left_grid_pin_44_ sb_2__5_/top_left_grid_pin_45_ sb_2__6_/bottom_left_grid_pin_45_
+ sb_2__5_/top_left_grid_pin_46_ sb_2__6_/bottom_left_grid_pin_46_ sb_2__5_/top_left_grid_pin_47_
+ sb_2__6_/bottom_left_grid_pin_47_ sb_2__5_/top_left_grid_pin_48_ sb_2__6_/bottom_left_grid_pin_48_
+ sb_2__5_/top_left_grid_pin_49_ sb_2__6_/bottom_left_grid_pin_49_ cbx_2__6_/bottom_grid_pin_0_
+ cbx_2__6_/bottom_grid_pin_10_ cbx_2__6_/bottom_grid_pin_11_ cbx_2__6_/bottom_grid_pin_12_
+ cbx_2__6_/bottom_grid_pin_13_ cbx_2__6_/bottom_grid_pin_14_ cbx_2__6_/bottom_grid_pin_15_
+ cbx_2__6_/bottom_grid_pin_1_ cbx_2__6_/bottom_grid_pin_2_ cbx_2__6_/REGOUT_FEEDTHROUGH
+ grid_clb_2__6_/top_width_0_height_0__pin_33_ sb_2__6_/left_bottom_grid_pin_34_ sb_1__6_/right_bottom_grid_pin_34_
+ sb_2__6_/left_bottom_grid_pin_35_ sb_1__6_/right_bottom_grid_pin_35_ sb_2__6_/left_bottom_grid_pin_36_
+ sb_1__6_/right_bottom_grid_pin_36_ sb_2__6_/left_bottom_grid_pin_37_ sb_1__6_/right_bottom_grid_pin_37_
+ sb_2__6_/left_bottom_grid_pin_38_ sb_1__6_/right_bottom_grid_pin_38_ sb_2__6_/left_bottom_grid_pin_39_
+ sb_1__6_/right_bottom_grid_pin_39_ cbx_2__6_/bottom_grid_pin_3_ sb_2__6_/left_bottom_grid_pin_40_
+ sb_1__6_/right_bottom_grid_pin_40_ sb_2__6_/left_bottom_grid_pin_41_ sb_1__6_/right_bottom_grid_pin_41_
+ cbx_2__6_/bottom_grid_pin_4_ cbx_2__6_/bottom_grid_pin_5_ cbx_2__6_/bottom_grid_pin_6_
+ cbx_2__6_/bottom_grid_pin_7_ cbx_2__6_/bottom_grid_pin_8_ cbx_2__6_/bottom_grid_pin_9_
+ grid_clb
Xsb_7__3_ sb_7__3_/Test_en_N_out sb_7__3_/Test_en_S_in VGND VPWR sb_7__3_/bottom_left_grid_pin_42_
+ sb_7__3_/bottom_left_grid_pin_43_ sb_7__3_/bottom_left_grid_pin_44_ sb_7__3_/bottom_left_grid_pin_45_
+ sb_7__3_/bottom_left_grid_pin_46_ sb_7__3_/bottom_left_grid_pin_47_ sb_7__3_/bottom_left_grid_pin_48_
+ sb_7__3_/bottom_left_grid_pin_49_ sb_7__3_/ccff_head sb_7__3_/ccff_tail sb_7__3_/chanx_left_in[0]
+ sb_7__3_/chanx_left_in[10] sb_7__3_/chanx_left_in[11] sb_7__3_/chanx_left_in[12]
+ sb_7__3_/chanx_left_in[13] sb_7__3_/chanx_left_in[14] sb_7__3_/chanx_left_in[15]
+ sb_7__3_/chanx_left_in[16] sb_7__3_/chanx_left_in[17] sb_7__3_/chanx_left_in[18]
+ sb_7__3_/chanx_left_in[19] sb_7__3_/chanx_left_in[1] sb_7__3_/chanx_left_in[2] sb_7__3_/chanx_left_in[3]
+ sb_7__3_/chanx_left_in[4] sb_7__3_/chanx_left_in[5] sb_7__3_/chanx_left_in[6] sb_7__3_/chanx_left_in[7]
+ sb_7__3_/chanx_left_in[8] sb_7__3_/chanx_left_in[9] sb_7__3_/chanx_left_out[0] sb_7__3_/chanx_left_out[10]
+ sb_7__3_/chanx_left_out[11] sb_7__3_/chanx_left_out[12] sb_7__3_/chanx_left_out[13]
+ sb_7__3_/chanx_left_out[14] sb_7__3_/chanx_left_out[15] sb_7__3_/chanx_left_out[16]
+ sb_7__3_/chanx_left_out[17] sb_7__3_/chanx_left_out[18] sb_7__3_/chanx_left_out[19]
+ sb_7__3_/chanx_left_out[1] sb_7__3_/chanx_left_out[2] sb_7__3_/chanx_left_out[3]
+ sb_7__3_/chanx_left_out[4] sb_7__3_/chanx_left_out[5] sb_7__3_/chanx_left_out[6]
+ sb_7__3_/chanx_left_out[7] sb_7__3_/chanx_left_out[8] sb_7__3_/chanx_left_out[9]
+ sb_7__3_/chanx_right_in[0] sb_7__3_/chanx_right_in[10] sb_7__3_/chanx_right_in[11]
+ sb_7__3_/chanx_right_in[12] sb_7__3_/chanx_right_in[13] sb_7__3_/chanx_right_in[14]
+ sb_7__3_/chanx_right_in[15] sb_7__3_/chanx_right_in[16] sb_7__3_/chanx_right_in[17]
+ sb_7__3_/chanx_right_in[18] sb_7__3_/chanx_right_in[19] sb_7__3_/chanx_right_in[1]
+ sb_7__3_/chanx_right_in[2] sb_7__3_/chanx_right_in[3] sb_7__3_/chanx_right_in[4]
+ sb_7__3_/chanx_right_in[5] sb_7__3_/chanx_right_in[6] sb_7__3_/chanx_right_in[7]
+ sb_7__3_/chanx_right_in[8] sb_7__3_/chanx_right_in[9] cbx_8__3_/chanx_left_in[0]
+ cbx_8__3_/chanx_left_in[10] cbx_8__3_/chanx_left_in[11] cbx_8__3_/chanx_left_in[12]
+ cbx_8__3_/chanx_left_in[13] cbx_8__3_/chanx_left_in[14] cbx_8__3_/chanx_left_in[15]
+ cbx_8__3_/chanx_left_in[16] cbx_8__3_/chanx_left_in[17] cbx_8__3_/chanx_left_in[18]
+ cbx_8__3_/chanx_left_in[19] cbx_8__3_/chanx_left_in[1] cbx_8__3_/chanx_left_in[2]
+ cbx_8__3_/chanx_left_in[3] cbx_8__3_/chanx_left_in[4] cbx_8__3_/chanx_left_in[5]
+ cbx_8__3_/chanx_left_in[6] cbx_8__3_/chanx_left_in[7] cbx_8__3_/chanx_left_in[8]
+ cbx_8__3_/chanx_left_in[9] cby_7__3_/chany_top_out[0] cby_7__3_/chany_top_out[10]
+ cby_7__3_/chany_top_out[11] cby_7__3_/chany_top_out[12] cby_7__3_/chany_top_out[13]
+ cby_7__3_/chany_top_out[14] cby_7__3_/chany_top_out[15] cby_7__3_/chany_top_out[16]
+ cby_7__3_/chany_top_out[17] cby_7__3_/chany_top_out[18] cby_7__3_/chany_top_out[19]
+ cby_7__3_/chany_top_out[1] cby_7__3_/chany_top_out[2] cby_7__3_/chany_top_out[3]
+ cby_7__3_/chany_top_out[4] cby_7__3_/chany_top_out[5] cby_7__3_/chany_top_out[6]
+ cby_7__3_/chany_top_out[7] cby_7__3_/chany_top_out[8] cby_7__3_/chany_top_out[9]
+ cby_7__3_/chany_top_in[0] cby_7__3_/chany_top_in[10] cby_7__3_/chany_top_in[11]
+ cby_7__3_/chany_top_in[12] cby_7__3_/chany_top_in[13] cby_7__3_/chany_top_in[14]
+ cby_7__3_/chany_top_in[15] cby_7__3_/chany_top_in[16] cby_7__3_/chany_top_in[17]
+ cby_7__3_/chany_top_in[18] cby_7__3_/chany_top_in[19] cby_7__3_/chany_top_in[1]
+ cby_7__3_/chany_top_in[2] cby_7__3_/chany_top_in[3] cby_7__3_/chany_top_in[4] cby_7__3_/chany_top_in[5]
+ cby_7__3_/chany_top_in[6] cby_7__3_/chany_top_in[7] cby_7__3_/chany_top_in[8] cby_7__3_/chany_top_in[9]
+ sb_7__3_/chany_top_in[0] sb_7__3_/chany_top_in[10] sb_7__3_/chany_top_in[11] sb_7__3_/chany_top_in[12]
+ sb_7__3_/chany_top_in[13] sb_7__3_/chany_top_in[14] sb_7__3_/chany_top_in[15] sb_7__3_/chany_top_in[16]
+ sb_7__3_/chany_top_in[17] sb_7__3_/chany_top_in[18] sb_7__3_/chany_top_in[19] sb_7__3_/chany_top_in[1]
+ sb_7__3_/chany_top_in[2] sb_7__3_/chany_top_in[3] sb_7__3_/chany_top_in[4] sb_7__3_/chany_top_in[5]
+ sb_7__3_/chany_top_in[6] sb_7__3_/chany_top_in[7] sb_7__3_/chany_top_in[8] sb_7__3_/chany_top_in[9]
+ sb_7__3_/chany_top_out[0] sb_7__3_/chany_top_out[10] sb_7__3_/chany_top_out[11]
+ sb_7__3_/chany_top_out[12] sb_7__3_/chany_top_out[13] sb_7__3_/chany_top_out[14]
+ sb_7__3_/chany_top_out[15] sb_7__3_/chany_top_out[16] sb_7__3_/chany_top_out[17]
+ sb_7__3_/chany_top_out[18] sb_7__3_/chany_top_out[19] sb_7__3_/chany_top_out[1]
+ sb_7__3_/chany_top_out[2] sb_7__3_/chany_top_out[3] sb_7__3_/chany_top_out[4] sb_7__3_/chany_top_out[5]
+ sb_7__3_/chany_top_out[6] sb_7__3_/chany_top_out[7] sb_7__3_/chany_top_out[8] sb_7__3_/chany_top_out[9]
+ sb_7__3_/clk_1_E_out sb_7__3_/clk_1_N_in sb_7__3_/clk_1_W_out sb_7__3_/clk_2_E_out
+ sb_7__3_/clk_2_N_in sb_7__3_/clk_2_N_out sb_7__3_/clk_2_S_out sb_7__3_/clk_2_W_out
+ sb_7__3_/clk_3_E_out sb_7__3_/clk_3_N_in sb_7__3_/clk_3_N_out sb_7__3_/clk_3_S_out
+ sb_7__3_/clk_3_W_out sb_7__3_/left_bottom_grid_pin_34_ sb_7__3_/left_bottom_grid_pin_35_
+ sb_7__3_/left_bottom_grid_pin_36_ sb_7__3_/left_bottom_grid_pin_37_ sb_7__3_/left_bottom_grid_pin_38_
+ sb_7__3_/left_bottom_grid_pin_39_ sb_7__3_/left_bottom_grid_pin_40_ sb_7__3_/left_bottom_grid_pin_41_
+ sb_7__3_/prog_clk_0_N_in sb_7__3_/prog_clk_1_E_out sb_7__3_/prog_clk_1_N_in sb_7__3_/prog_clk_1_W_out
+ sb_7__3_/prog_clk_2_E_out sb_7__3_/prog_clk_2_N_in sb_7__3_/prog_clk_2_N_out sb_7__3_/prog_clk_2_S_out
+ sb_7__3_/prog_clk_2_W_out sb_7__3_/prog_clk_3_E_out sb_7__3_/prog_clk_3_N_in sb_7__3_/prog_clk_3_N_out
+ sb_7__3_/prog_clk_3_S_out sb_7__3_/prog_clk_3_W_out sb_7__3_/right_bottom_grid_pin_34_
+ sb_7__3_/right_bottom_grid_pin_35_ sb_7__3_/right_bottom_grid_pin_36_ sb_7__3_/right_bottom_grid_pin_37_
+ sb_7__3_/right_bottom_grid_pin_38_ sb_7__3_/right_bottom_grid_pin_39_ sb_7__3_/right_bottom_grid_pin_40_
+ sb_7__3_/right_bottom_grid_pin_41_ sb_7__3_/top_left_grid_pin_42_ sb_7__3_/top_left_grid_pin_43_
+ sb_7__3_/top_left_grid_pin_44_ sb_7__3_/top_left_grid_pin_45_ sb_7__3_/top_left_grid_pin_46_
+ sb_7__3_/top_left_grid_pin_47_ sb_7__3_/top_left_grid_pin_48_ sb_7__3_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_4__0_ sb_4__0_/SC_IN_TOP sb_4__0_/SC_OUT_TOP sb_4__0_/Test_en_N_out Test_en VGND
+ VPWR sb_4__0_/ccff_head sb_4__0_/ccff_tail sb_4__0_/chanx_left_in[0] sb_4__0_/chanx_left_in[10]
+ sb_4__0_/chanx_left_in[11] sb_4__0_/chanx_left_in[12] sb_4__0_/chanx_left_in[13]
+ sb_4__0_/chanx_left_in[14] sb_4__0_/chanx_left_in[15] sb_4__0_/chanx_left_in[16]
+ sb_4__0_/chanx_left_in[17] sb_4__0_/chanx_left_in[18] sb_4__0_/chanx_left_in[19]
+ sb_4__0_/chanx_left_in[1] sb_4__0_/chanx_left_in[2] sb_4__0_/chanx_left_in[3] sb_4__0_/chanx_left_in[4]
+ sb_4__0_/chanx_left_in[5] sb_4__0_/chanx_left_in[6] sb_4__0_/chanx_left_in[7] sb_4__0_/chanx_left_in[8]
+ sb_4__0_/chanx_left_in[9] sb_4__0_/chanx_left_out[0] sb_4__0_/chanx_left_out[10]
+ sb_4__0_/chanx_left_out[11] sb_4__0_/chanx_left_out[12] sb_4__0_/chanx_left_out[13]
+ sb_4__0_/chanx_left_out[14] sb_4__0_/chanx_left_out[15] sb_4__0_/chanx_left_out[16]
+ sb_4__0_/chanx_left_out[17] sb_4__0_/chanx_left_out[18] sb_4__0_/chanx_left_out[19]
+ sb_4__0_/chanx_left_out[1] sb_4__0_/chanx_left_out[2] sb_4__0_/chanx_left_out[3]
+ sb_4__0_/chanx_left_out[4] sb_4__0_/chanx_left_out[5] sb_4__0_/chanx_left_out[6]
+ sb_4__0_/chanx_left_out[7] sb_4__0_/chanx_left_out[8] sb_4__0_/chanx_left_out[9]
+ sb_4__0_/chanx_right_in[0] sb_4__0_/chanx_right_in[10] sb_4__0_/chanx_right_in[11]
+ sb_4__0_/chanx_right_in[12] sb_4__0_/chanx_right_in[13] sb_4__0_/chanx_right_in[14]
+ sb_4__0_/chanx_right_in[15] sb_4__0_/chanx_right_in[16] sb_4__0_/chanx_right_in[17]
+ sb_4__0_/chanx_right_in[18] sb_4__0_/chanx_right_in[19] sb_4__0_/chanx_right_in[1]
+ sb_4__0_/chanx_right_in[2] sb_4__0_/chanx_right_in[3] sb_4__0_/chanx_right_in[4]
+ sb_4__0_/chanx_right_in[5] sb_4__0_/chanx_right_in[6] sb_4__0_/chanx_right_in[7]
+ sb_4__0_/chanx_right_in[8] sb_4__0_/chanx_right_in[9] cbx_5__0_/chanx_left_in[0]
+ cbx_5__0_/chanx_left_in[10] cbx_5__0_/chanx_left_in[11] cbx_5__0_/chanx_left_in[12]
+ cbx_5__0_/chanx_left_in[13] cbx_5__0_/chanx_left_in[14] cbx_5__0_/chanx_left_in[15]
+ cbx_5__0_/chanx_left_in[16] cbx_5__0_/chanx_left_in[17] cbx_5__0_/chanx_left_in[18]
+ cbx_5__0_/chanx_left_in[19] cbx_5__0_/chanx_left_in[1] cbx_5__0_/chanx_left_in[2]
+ cbx_5__0_/chanx_left_in[3] cbx_5__0_/chanx_left_in[4] cbx_5__0_/chanx_left_in[5]
+ cbx_5__0_/chanx_left_in[6] cbx_5__0_/chanx_left_in[7] cbx_5__0_/chanx_left_in[8]
+ cbx_5__0_/chanx_left_in[9] sb_4__0_/chany_top_in[0] sb_4__0_/chany_top_in[10] sb_4__0_/chany_top_in[11]
+ sb_4__0_/chany_top_in[12] sb_4__0_/chany_top_in[13] sb_4__0_/chany_top_in[14] sb_4__0_/chany_top_in[15]
+ sb_4__0_/chany_top_in[16] sb_4__0_/chany_top_in[17] sb_4__0_/chany_top_in[18] sb_4__0_/chany_top_in[19]
+ sb_4__0_/chany_top_in[1] sb_4__0_/chany_top_in[2] sb_4__0_/chany_top_in[3] sb_4__0_/chany_top_in[4]
+ sb_4__0_/chany_top_in[5] sb_4__0_/chany_top_in[6] sb_4__0_/chany_top_in[7] sb_4__0_/chany_top_in[8]
+ sb_4__0_/chany_top_in[9] sb_4__0_/chany_top_out[0] sb_4__0_/chany_top_out[10] sb_4__0_/chany_top_out[11]
+ sb_4__0_/chany_top_out[12] sb_4__0_/chany_top_out[13] sb_4__0_/chany_top_out[14]
+ sb_4__0_/chany_top_out[15] sb_4__0_/chany_top_out[16] sb_4__0_/chany_top_out[17]
+ sb_4__0_/chany_top_out[18] sb_4__0_/chany_top_out[19] sb_4__0_/chany_top_out[1]
+ sb_4__0_/chany_top_out[2] sb_4__0_/chany_top_out[3] sb_4__0_/chany_top_out[4] sb_4__0_/chany_top_out[5]
+ sb_4__0_/chany_top_out[6] sb_4__0_/chany_top_out[7] sb_4__0_/chany_top_out[8] sb_4__0_/chany_top_out[9]
+ sb_4__0_/clk_3_N_out clk sb_4__0_/left_bottom_grid_pin_11_ sb_4__0_/left_bottom_grid_pin_13_
+ sb_4__0_/left_bottom_grid_pin_15_ sb_4__0_/left_bottom_grid_pin_17_ sb_4__0_/left_bottom_grid_pin_1_
+ sb_4__0_/left_bottom_grid_pin_3_ sb_4__0_/left_bottom_grid_pin_5_ sb_4__0_/left_bottom_grid_pin_7_
+ sb_4__0_/left_bottom_grid_pin_9_ sb_4__0_/prog_clk_0_N_in sb_4__0_/prog_clk_3_N_out
+ prog_clk sb_4__0_/right_bottom_grid_pin_11_ sb_4__0_/right_bottom_grid_pin_13_ sb_4__0_/right_bottom_grid_pin_15_
+ sb_4__0_/right_bottom_grid_pin_17_ sb_4__0_/right_bottom_grid_pin_1_ sb_4__0_/right_bottom_grid_pin_3_
+ sb_4__0_/right_bottom_grid_pin_5_ sb_4__0_/right_bottom_grid_pin_7_ sb_4__0_/right_bottom_grid_pin_9_
+ sb_4__0_/top_left_grid_pin_42_ sb_4__0_/top_left_grid_pin_43_ sb_4__0_/top_left_grid_pin_44_
+ sb_4__0_/top_left_grid_pin_45_ sb_4__0_/top_left_grid_pin_46_ sb_4__0_/top_left_grid_pin_47_
+ sb_4__0_/top_left_grid_pin_48_ sb_4__0_/top_left_grid_pin_49_ sb_1__0_
Xsb_0__8_ sc_head sb_0__8_/SC_OUT_BOT VGND VPWR sb_0__8_/bottom_left_grid_pin_1_ sb_0__8_/ccff_head
+ sb_0__8_/ccff_tail sb_0__8_/chanx_right_in[0] sb_0__8_/chanx_right_in[10] sb_0__8_/chanx_right_in[11]
+ sb_0__8_/chanx_right_in[12] sb_0__8_/chanx_right_in[13] sb_0__8_/chanx_right_in[14]
+ sb_0__8_/chanx_right_in[15] sb_0__8_/chanx_right_in[16] sb_0__8_/chanx_right_in[17]
+ sb_0__8_/chanx_right_in[18] sb_0__8_/chanx_right_in[19] sb_0__8_/chanx_right_in[1]
+ sb_0__8_/chanx_right_in[2] sb_0__8_/chanx_right_in[3] sb_0__8_/chanx_right_in[4]
+ sb_0__8_/chanx_right_in[5] sb_0__8_/chanx_right_in[6] sb_0__8_/chanx_right_in[7]
+ sb_0__8_/chanx_right_in[8] sb_0__8_/chanx_right_in[9] cbx_1__8_/chanx_left_in[0]
+ cbx_1__8_/chanx_left_in[10] cbx_1__8_/chanx_left_in[11] cbx_1__8_/chanx_left_in[12]
+ cbx_1__8_/chanx_left_in[13] cbx_1__8_/chanx_left_in[14] cbx_1__8_/chanx_left_in[15]
+ cbx_1__8_/chanx_left_in[16] cbx_1__8_/chanx_left_in[17] cbx_1__8_/chanx_left_in[18]
+ cbx_1__8_/chanx_left_in[19] cbx_1__8_/chanx_left_in[1] cbx_1__8_/chanx_left_in[2]
+ cbx_1__8_/chanx_left_in[3] cbx_1__8_/chanx_left_in[4] cbx_1__8_/chanx_left_in[5]
+ cbx_1__8_/chanx_left_in[6] cbx_1__8_/chanx_left_in[7] cbx_1__8_/chanx_left_in[8]
+ cbx_1__8_/chanx_left_in[9] cby_0__8_/chany_top_out[0] cby_0__8_/chany_top_out[10]
+ cby_0__8_/chany_top_out[11] cby_0__8_/chany_top_out[12] cby_0__8_/chany_top_out[13]
+ cby_0__8_/chany_top_out[14] cby_0__8_/chany_top_out[15] cby_0__8_/chany_top_out[16]
+ cby_0__8_/chany_top_out[17] cby_0__8_/chany_top_out[18] cby_0__8_/chany_top_out[19]
+ cby_0__8_/chany_top_out[1] cby_0__8_/chany_top_out[2] cby_0__8_/chany_top_out[3]
+ cby_0__8_/chany_top_out[4] cby_0__8_/chany_top_out[5] cby_0__8_/chany_top_out[6]
+ cby_0__8_/chany_top_out[7] cby_0__8_/chany_top_out[8] cby_0__8_/chany_top_out[9]
+ cby_0__8_/chany_top_in[0] cby_0__8_/chany_top_in[10] cby_0__8_/chany_top_in[11]
+ cby_0__8_/chany_top_in[12] cby_0__8_/chany_top_in[13] cby_0__8_/chany_top_in[14]
+ cby_0__8_/chany_top_in[15] cby_0__8_/chany_top_in[16] cby_0__8_/chany_top_in[17]
+ cby_0__8_/chany_top_in[18] cby_0__8_/chany_top_in[19] cby_0__8_/chany_top_in[1]
+ cby_0__8_/chany_top_in[2] cby_0__8_/chany_top_in[3] cby_0__8_/chany_top_in[4] cby_0__8_/chany_top_in[5]
+ cby_0__8_/chany_top_in[6] cby_0__8_/chany_top_in[7] cby_0__8_/chany_top_in[8] cby_0__8_/chany_top_in[9]
+ sb_0__8_/prog_clk_0_E_in sb_0__8_/right_bottom_grid_pin_34_ sb_0__8_/right_bottom_grid_pin_35_
+ sb_0__8_/right_bottom_grid_pin_36_ sb_0__8_/right_bottom_grid_pin_37_ sb_0__8_/right_bottom_grid_pin_38_
+ sb_0__8_/right_bottom_grid_pin_39_ sb_0__8_/right_bottom_grid_pin_40_ sb_0__8_/right_bottom_grid_pin_41_
+ sb_0__8_/right_top_grid_pin_1_ sb_0__2_
Xcby_6__7_ cby_6__7_/Test_en_W_in cby_6__7_/Test_en_E_out cby_6__7_/Test_en_N_out
+ cby_6__7_/Test_en_W_in cby_6__7_/Test_en_W_in cby_6__7_/Test_en_W_out VGND VPWR
+ cby_6__7_/ccff_head cby_6__7_/ccff_tail sb_6__6_/chany_top_out[0] sb_6__6_/chany_top_out[10]
+ sb_6__6_/chany_top_out[11] sb_6__6_/chany_top_out[12] sb_6__6_/chany_top_out[13]
+ sb_6__6_/chany_top_out[14] sb_6__6_/chany_top_out[15] sb_6__6_/chany_top_out[16]
+ sb_6__6_/chany_top_out[17] sb_6__6_/chany_top_out[18] sb_6__6_/chany_top_out[19]
+ sb_6__6_/chany_top_out[1] sb_6__6_/chany_top_out[2] sb_6__6_/chany_top_out[3] sb_6__6_/chany_top_out[4]
+ sb_6__6_/chany_top_out[5] sb_6__6_/chany_top_out[6] sb_6__6_/chany_top_out[7] sb_6__6_/chany_top_out[8]
+ sb_6__6_/chany_top_out[9] sb_6__6_/chany_top_in[0] sb_6__6_/chany_top_in[10] sb_6__6_/chany_top_in[11]
+ sb_6__6_/chany_top_in[12] sb_6__6_/chany_top_in[13] sb_6__6_/chany_top_in[14] sb_6__6_/chany_top_in[15]
+ sb_6__6_/chany_top_in[16] sb_6__6_/chany_top_in[17] sb_6__6_/chany_top_in[18] sb_6__6_/chany_top_in[19]
+ sb_6__6_/chany_top_in[1] sb_6__6_/chany_top_in[2] sb_6__6_/chany_top_in[3] sb_6__6_/chany_top_in[4]
+ sb_6__6_/chany_top_in[5] sb_6__6_/chany_top_in[6] sb_6__6_/chany_top_in[7] sb_6__6_/chany_top_in[8]
+ sb_6__6_/chany_top_in[9] cby_6__7_/chany_top_in[0] cby_6__7_/chany_top_in[10] cby_6__7_/chany_top_in[11]
+ cby_6__7_/chany_top_in[12] cby_6__7_/chany_top_in[13] cby_6__7_/chany_top_in[14]
+ cby_6__7_/chany_top_in[15] cby_6__7_/chany_top_in[16] cby_6__7_/chany_top_in[17]
+ cby_6__7_/chany_top_in[18] cby_6__7_/chany_top_in[19] cby_6__7_/chany_top_in[1]
+ cby_6__7_/chany_top_in[2] cby_6__7_/chany_top_in[3] cby_6__7_/chany_top_in[4] cby_6__7_/chany_top_in[5]
+ cby_6__7_/chany_top_in[6] cby_6__7_/chany_top_in[7] cby_6__7_/chany_top_in[8] cby_6__7_/chany_top_in[9]
+ cby_6__7_/chany_top_out[0] cby_6__7_/chany_top_out[10] cby_6__7_/chany_top_out[11]
+ cby_6__7_/chany_top_out[12] cby_6__7_/chany_top_out[13] cby_6__7_/chany_top_out[14]
+ cby_6__7_/chany_top_out[15] cby_6__7_/chany_top_out[16] cby_6__7_/chany_top_out[17]
+ cby_6__7_/chany_top_out[18] cby_6__7_/chany_top_out[19] cby_6__7_/chany_top_out[1]
+ cby_6__7_/chany_top_out[2] cby_6__7_/chany_top_out[3] cby_6__7_/chany_top_out[4]
+ cby_6__7_/chany_top_out[5] cby_6__7_/chany_top_out[6] cby_6__7_/chany_top_out[7]
+ cby_6__7_/chany_top_out[8] cby_6__7_/chany_top_out[9] cby_6__7_/clk_2_N_out cby_6__7_/clk_2_S_in
+ cby_6__7_/clk_2_S_out cby_6__7_/clk_3_N_out cby_6__7_/clk_3_S_in cby_6__7_/clk_3_S_out
+ cby_6__7_/left_grid_pin_16_ cby_6__7_/left_grid_pin_17_ cby_6__7_/left_grid_pin_18_
+ cby_6__7_/left_grid_pin_19_ cby_6__7_/left_grid_pin_20_ cby_6__7_/left_grid_pin_21_
+ cby_6__7_/left_grid_pin_22_ cby_6__7_/left_grid_pin_23_ cby_6__7_/left_grid_pin_24_
+ cby_6__7_/left_grid_pin_25_ cby_6__7_/left_grid_pin_26_ cby_6__7_/left_grid_pin_27_
+ cby_6__7_/left_grid_pin_28_ cby_6__7_/left_grid_pin_29_ cby_6__7_/left_grid_pin_30_
+ cby_6__7_/left_grid_pin_31_ cby_6__7_/prog_clk_0_N_out sb_6__6_/prog_clk_0_N_in
+ cby_6__7_/prog_clk_0_W_in cby_6__7_/prog_clk_2_N_out cby_6__7_/prog_clk_2_S_in cby_6__7_/prog_clk_2_S_out
+ cby_6__7_/prog_clk_3_N_out cby_6__7_/prog_clk_3_S_in cby_6__7_/prog_clk_3_S_out
+ cby_1__1_
Xcby_3__4_ cby_3__4_/Test_en_W_in cby_3__4_/Test_en_E_out cby_3__4_/Test_en_N_out
+ cby_3__4_/Test_en_W_in cby_3__4_/Test_en_W_in cby_3__4_/Test_en_W_out VGND VPWR
+ cby_3__4_/ccff_head cby_3__4_/ccff_tail sb_3__3_/chany_top_out[0] sb_3__3_/chany_top_out[10]
+ sb_3__3_/chany_top_out[11] sb_3__3_/chany_top_out[12] sb_3__3_/chany_top_out[13]
+ sb_3__3_/chany_top_out[14] sb_3__3_/chany_top_out[15] sb_3__3_/chany_top_out[16]
+ sb_3__3_/chany_top_out[17] sb_3__3_/chany_top_out[18] sb_3__3_/chany_top_out[19]
+ sb_3__3_/chany_top_out[1] sb_3__3_/chany_top_out[2] sb_3__3_/chany_top_out[3] sb_3__3_/chany_top_out[4]
+ sb_3__3_/chany_top_out[5] sb_3__3_/chany_top_out[6] sb_3__3_/chany_top_out[7] sb_3__3_/chany_top_out[8]
+ sb_3__3_/chany_top_out[9] sb_3__3_/chany_top_in[0] sb_3__3_/chany_top_in[10] sb_3__3_/chany_top_in[11]
+ sb_3__3_/chany_top_in[12] sb_3__3_/chany_top_in[13] sb_3__3_/chany_top_in[14] sb_3__3_/chany_top_in[15]
+ sb_3__3_/chany_top_in[16] sb_3__3_/chany_top_in[17] sb_3__3_/chany_top_in[18] sb_3__3_/chany_top_in[19]
+ sb_3__3_/chany_top_in[1] sb_3__3_/chany_top_in[2] sb_3__3_/chany_top_in[3] sb_3__3_/chany_top_in[4]
+ sb_3__3_/chany_top_in[5] sb_3__3_/chany_top_in[6] sb_3__3_/chany_top_in[7] sb_3__3_/chany_top_in[8]
+ sb_3__3_/chany_top_in[9] cby_3__4_/chany_top_in[0] cby_3__4_/chany_top_in[10] cby_3__4_/chany_top_in[11]
+ cby_3__4_/chany_top_in[12] cby_3__4_/chany_top_in[13] cby_3__4_/chany_top_in[14]
+ cby_3__4_/chany_top_in[15] cby_3__4_/chany_top_in[16] cby_3__4_/chany_top_in[17]
+ cby_3__4_/chany_top_in[18] cby_3__4_/chany_top_in[19] cby_3__4_/chany_top_in[1]
+ cby_3__4_/chany_top_in[2] cby_3__4_/chany_top_in[3] cby_3__4_/chany_top_in[4] cby_3__4_/chany_top_in[5]
+ cby_3__4_/chany_top_in[6] cby_3__4_/chany_top_in[7] cby_3__4_/chany_top_in[8] cby_3__4_/chany_top_in[9]
+ cby_3__4_/chany_top_out[0] cby_3__4_/chany_top_out[10] cby_3__4_/chany_top_out[11]
+ cby_3__4_/chany_top_out[12] cby_3__4_/chany_top_out[13] cby_3__4_/chany_top_out[14]
+ cby_3__4_/chany_top_out[15] cby_3__4_/chany_top_out[16] cby_3__4_/chany_top_out[17]
+ cby_3__4_/chany_top_out[18] cby_3__4_/chany_top_out[19] cby_3__4_/chany_top_out[1]
+ cby_3__4_/chany_top_out[2] cby_3__4_/chany_top_out[3] cby_3__4_/chany_top_out[4]
+ cby_3__4_/chany_top_out[5] cby_3__4_/chany_top_out[6] cby_3__4_/chany_top_out[7]
+ cby_3__4_/chany_top_out[8] cby_3__4_/chany_top_out[9] cby_3__4_/clk_2_N_out cby_3__4_/clk_2_S_in
+ cby_3__4_/clk_2_S_out cby_3__4_/clk_3_N_out cby_3__4_/clk_3_S_in cby_3__4_/clk_3_S_out
+ cby_3__4_/left_grid_pin_16_ cby_3__4_/left_grid_pin_17_ cby_3__4_/left_grid_pin_18_
+ cby_3__4_/left_grid_pin_19_ cby_3__4_/left_grid_pin_20_ cby_3__4_/left_grid_pin_21_
+ cby_3__4_/left_grid_pin_22_ cby_3__4_/left_grid_pin_23_ cby_3__4_/left_grid_pin_24_
+ cby_3__4_/left_grid_pin_25_ cby_3__4_/left_grid_pin_26_ cby_3__4_/left_grid_pin_27_
+ cby_3__4_/left_grid_pin_28_ cby_3__4_/left_grid_pin_29_ cby_3__4_/left_grid_pin_30_
+ cby_3__4_/left_grid_pin_31_ cby_3__4_/prog_clk_0_N_out sb_3__3_/prog_clk_0_N_in
+ cby_3__4_/prog_clk_0_W_in cby_3__4_/prog_clk_2_N_out cby_3__4_/prog_clk_2_S_in cby_3__4_/prog_clk_2_S_out
+ cby_3__4_/prog_clk_3_N_out cby_3__4_/prog_clk_3_S_in cby_3__4_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_6__8_ IO_ISOL_N cbx_6__8_/SC_IN_BOT cbx_6__8_/SC_IN_TOP cbx_6__8_/SC_OUT_BOT
+ sb_6__8_/SC_IN_BOT VGND VPWR cbx_6__8_/bottom_grid_pin_0_ cbx_6__8_/bottom_grid_pin_10_
+ cbx_6__8_/bottom_grid_pin_11_ cbx_6__8_/bottom_grid_pin_12_ cbx_6__8_/bottom_grid_pin_13_
+ cbx_6__8_/bottom_grid_pin_14_ cbx_6__8_/bottom_grid_pin_15_ cbx_6__8_/bottom_grid_pin_1_
+ cbx_6__8_/bottom_grid_pin_2_ cbx_6__8_/bottom_grid_pin_3_ cbx_6__8_/bottom_grid_pin_4_
+ cbx_6__8_/bottom_grid_pin_5_ cbx_6__8_/bottom_grid_pin_6_ cbx_6__8_/bottom_grid_pin_7_
+ cbx_6__8_/bottom_grid_pin_8_ cbx_6__8_/bottom_grid_pin_9_ cbx_6__8_/top_grid_pin_0_
+ sb_6__8_/left_top_grid_pin_1_ sb_5__8_/right_top_grid_pin_1_ sb_6__8_/ccff_tail
+ sb_5__8_/ccff_head cbx_6__8_/chanx_left_in[0] cbx_6__8_/chanx_left_in[10] cbx_6__8_/chanx_left_in[11]
+ cbx_6__8_/chanx_left_in[12] cbx_6__8_/chanx_left_in[13] cbx_6__8_/chanx_left_in[14]
+ cbx_6__8_/chanx_left_in[15] cbx_6__8_/chanx_left_in[16] cbx_6__8_/chanx_left_in[17]
+ cbx_6__8_/chanx_left_in[18] cbx_6__8_/chanx_left_in[19] cbx_6__8_/chanx_left_in[1]
+ cbx_6__8_/chanx_left_in[2] cbx_6__8_/chanx_left_in[3] cbx_6__8_/chanx_left_in[4]
+ cbx_6__8_/chanx_left_in[5] cbx_6__8_/chanx_left_in[6] cbx_6__8_/chanx_left_in[7]
+ cbx_6__8_/chanx_left_in[8] cbx_6__8_/chanx_left_in[9] sb_5__8_/chanx_right_in[0]
+ sb_5__8_/chanx_right_in[10] sb_5__8_/chanx_right_in[11] sb_5__8_/chanx_right_in[12]
+ sb_5__8_/chanx_right_in[13] sb_5__8_/chanx_right_in[14] sb_5__8_/chanx_right_in[15]
+ sb_5__8_/chanx_right_in[16] sb_5__8_/chanx_right_in[17] sb_5__8_/chanx_right_in[18]
+ sb_5__8_/chanx_right_in[19] sb_5__8_/chanx_right_in[1] sb_5__8_/chanx_right_in[2]
+ sb_5__8_/chanx_right_in[3] sb_5__8_/chanx_right_in[4] sb_5__8_/chanx_right_in[5]
+ sb_5__8_/chanx_right_in[6] sb_5__8_/chanx_right_in[7] sb_5__8_/chanx_right_in[8]
+ sb_5__8_/chanx_right_in[9] sb_6__8_/chanx_left_out[0] sb_6__8_/chanx_left_out[10]
+ sb_6__8_/chanx_left_out[11] sb_6__8_/chanx_left_out[12] sb_6__8_/chanx_left_out[13]
+ sb_6__8_/chanx_left_out[14] sb_6__8_/chanx_left_out[15] sb_6__8_/chanx_left_out[16]
+ sb_6__8_/chanx_left_out[17] sb_6__8_/chanx_left_out[18] sb_6__8_/chanx_left_out[19]
+ sb_6__8_/chanx_left_out[1] sb_6__8_/chanx_left_out[2] sb_6__8_/chanx_left_out[3]
+ sb_6__8_/chanx_left_out[4] sb_6__8_/chanx_left_out[5] sb_6__8_/chanx_left_out[6]
+ sb_6__8_/chanx_left_out[7] sb_6__8_/chanx_left_out[8] sb_6__8_/chanx_left_out[9]
+ sb_6__8_/chanx_left_in[0] sb_6__8_/chanx_left_in[10] sb_6__8_/chanx_left_in[11]
+ sb_6__8_/chanx_left_in[12] sb_6__8_/chanx_left_in[13] sb_6__8_/chanx_left_in[14]
+ sb_6__8_/chanx_left_in[15] sb_6__8_/chanx_left_in[16] sb_6__8_/chanx_left_in[17]
+ sb_6__8_/chanx_left_in[18] sb_6__8_/chanx_left_in[19] sb_6__8_/chanx_left_in[1]
+ sb_6__8_/chanx_left_in[2] sb_6__8_/chanx_left_in[3] sb_6__8_/chanx_left_in[4] sb_6__8_/chanx_left_in[5]
+ sb_6__8_/chanx_left_in[6] sb_6__8_/chanx_left_in[7] sb_6__8_/chanx_left_in[8] sb_6__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
+ cbx_6__8_/prog_clk_0_S_in cbx_6__8_/prog_clk_0_W_out cbx_6__8_/top_grid_pin_0_ cbx_1__2_
Xgrid_clb_5__8_ cbx_5__8_/SC_OUT_BOT cbx_5__7_/SC_IN_TOP grid_clb_5__8_/SC_OUT_TOP
+ cby_4__8_/Test_en_E_out cby_5__8_/Test_en_W_in cby_4__8_/Test_en_E_out grid_clb_5__8_/Test_en_W_out
+ VGND VPWR cbx_5__7_/REGIN_FEEDTHROUGH grid_clb_5__8_/bottom_width_0_height_0__pin_51_
+ cby_4__8_/ccff_tail cby_5__8_/ccff_head cbx_5__7_/clk_1_N_out cbx_5__7_/clk_1_N_out
+ cby_5__8_/prog_clk_0_W_in cbx_5__7_/prog_clk_1_N_out cbx_5__8_/prog_clk_0_S_in cbx_5__7_/prog_clk_1_N_out
+ cbx_5__7_/prog_clk_0_N_in grid_clb_5__8_/prog_clk_0_W_out cby_5__8_/left_grid_pin_16_
+ cby_5__8_/left_grid_pin_17_ cby_5__8_/left_grid_pin_18_ cby_5__8_/left_grid_pin_19_
+ cby_5__8_/left_grid_pin_20_ cby_5__8_/left_grid_pin_21_ cby_5__8_/left_grid_pin_22_
+ cby_5__8_/left_grid_pin_23_ cby_5__8_/left_grid_pin_24_ cby_5__8_/left_grid_pin_25_
+ cby_5__8_/left_grid_pin_26_ cby_5__8_/left_grid_pin_27_ cby_5__8_/left_grid_pin_28_
+ cby_5__8_/left_grid_pin_29_ cby_5__8_/left_grid_pin_30_ cby_5__8_/left_grid_pin_31_
+ sb_5__7_/top_left_grid_pin_42_ sb_5__8_/bottom_left_grid_pin_42_ sb_5__7_/top_left_grid_pin_43_
+ sb_5__8_/bottom_left_grid_pin_43_ sb_5__7_/top_left_grid_pin_44_ sb_5__8_/bottom_left_grid_pin_44_
+ sb_5__7_/top_left_grid_pin_45_ sb_5__8_/bottom_left_grid_pin_45_ sb_5__7_/top_left_grid_pin_46_
+ sb_5__8_/bottom_left_grid_pin_46_ sb_5__7_/top_left_grid_pin_47_ sb_5__8_/bottom_left_grid_pin_47_
+ sb_5__7_/top_left_grid_pin_48_ sb_5__8_/bottom_left_grid_pin_48_ sb_5__7_/top_left_grid_pin_49_
+ sb_5__8_/bottom_left_grid_pin_49_ cbx_5__8_/bottom_grid_pin_0_ cbx_5__8_/bottom_grid_pin_10_
+ cbx_5__8_/bottom_grid_pin_11_ cbx_5__8_/bottom_grid_pin_12_ cbx_5__8_/bottom_grid_pin_13_
+ cbx_5__8_/bottom_grid_pin_14_ cbx_5__8_/bottom_grid_pin_15_ cbx_5__8_/bottom_grid_pin_1_
+ cbx_5__8_/bottom_grid_pin_2_ tie_array/x[4] grid_clb_5__8_/top_width_0_height_0__pin_33_
+ sb_5__8_/left_bottom_grid_pin_34_ sb_4__8_/right_bottom_grid_pin_34_ sb_5__8_/left_bottom_grid_pin_35_
+ sb_4__8_/right_bottom_grid_pin_35_ sb_5__8_/left_bottom_grid_pin_36_ sb_4__8_/right_bottom_grid_pin_36_
+ sb_5__8_/left_bottom_grid_pin_37_ sb_4__8_/right_bottom_grid_pin_37_ sb_5__8_/left_bottom_grid_pin_38_
+ sb_4__8_/right_bottom_grid_pin_38_ sb_5__8_/left_bottom_grid_pin_39_ sb_4__8_/right_bottom_grid_pin_39_
+ cbx_5__8_/bottom_grid_pin_3_ sb_5__8_/left_bottom_grid_pin_40_ sb_4__8_/right_bottom_grid_pin_40_
+ sb_5__8_/left_bottom_grid_pin_41_ sb_4__8_/right_bottom_grid_pin_41_ cbx_5__8_/bottom_grid_pin_4_
+ cbx_5__8_/bottom_grid_pin_5_ cbx_5__8_/bottom_grid_pin_6_ cbx_5__8_/bottom_grid_pin_7_
+ cbx_5__8_/bottom_grid_pin_8_ cbx_5__8_/bottom_grid_pin_9_ grid_clb
Xcbx_3__5_ cbx_3__5_/REGIN_FEEDTHROUGH cbx_3__5_/REGOUT_FEEDTHROUGH cbx_3__5_/SC_IN_BOT
+ cbx_3__5_/SC_IN_TOP cbx_3__5_/SC_OUT_BOT cbx_3__5_/SC_OUT_TOP VGND VPWR cbx_3__5_/bottom_grid_pin_0_
+ cbx_3__5_/bottom_grid_pin_10_ cbx_3__5_/bottom_grid_pin_11_ cbx_3__5_/bottom_grid_pin_12_
+ cbx_3__5_/bottom_grid_pin_13_ cbx_3__5_/bottom_grid_pin_14_ cbx_3__5_/bottom_grid_pin_15_
+ cbx_3__5_/bottom_grid_pin_1_ cbx_3__5_/bottom_grid_pin_2_ cbx_3__5_/bottom_grid_pin_3_
+ cbx_3__5_/bottom_grid_pin_4_ cbx_3__5_/bottom_grid_pin_5_ cbx_3__5_/bottom_grid_pin_6_
+ cbx_3__5_/bottom_grid_pin_7_ cbx_3__5_/bottom_grid_pin_8_ cbx_3__5_/bottom_grid_pin_9_
+ sb_3__5_/ccff_tail sb_2__5_/ccff_head cbx_3__5_/chanx_left_in[0] cbx_3__5_/chanx_left_in[10]
+ cbx_3__5_/chanx_left_in[11] cbx_3__5_/chanx_left_in[12] cbx_3__5_/chanx_left_in[13]
+ cbx_3__5_/chanx_left_in[14] cbx_3__5_/chanx_left_in[15] cbx_3__5_/chanx_left_in[16]
+ cbx_3__5_/chanx_left_in[17] cbx_3__5_/chanx_left_in[18] cbx_3__5_/chanx_left_in[19]
+ cbx_3__5_/chanx_left_in[1] cbx_3__5_/chanx_left_in[2] cbx_3__5_/chanx_left_in[3]
+ cbx_3__5_/chanx_left_in[4] cbx_3__5_/chanx_left_in[5] cbx_3__5_/chanx_left_in[6]
+ cbx_3__5_/chanx_left_in[7] cbx_3__5_/chanx_left_in[8] cbx_3__5_/chanx_left_in[9]
+ sb_2__5_/chanx_right_in[0] sb_2__5_/chanx_right_in[10] sb_2__5_/chanx_right_in[11]
+ sb_2__5_/chanx_right_in[12] sb_2__5_/chanx_right_in[13] sb_2__5_/chanx_right_in[14]
+ sb_2__5_/chanx_right_in[15] sb_2__5_/chanx_right_in[16] sb_2__5_/chanx_right_in[17]
+ sb_2__5_/chanx_right_in[18] sb_2__5_/chanx_right_in[19] sb_2__5_/chanx_right_in[1]
+ sb_2__5_/chanx_right_in[2] sb_2__5_/chanx_right_in[3] sb_2__5_/chanx_right_in[4]
+ sb_2__5_/chanx_right_in[5] sb_2__5_/chanx_right_in[6] sb_2__5_/chanx_right_in[7]
+ sb_2__5_/chanx_right_in[8] sb_2__5_/chanx_right_in[9] sb_3__5_/chanx_left_out[0]
+ sb_3__5_/chanx_left_out[10] sb_3__5_/chanx_left_out[11] sb_3__5_/chanx_left_out[12]
+ sb_3__5_/chanx_left_out[13] sb_3__5_/chanx_left_out[14] sb_3__5_/chanx_left_out[15]
+ sb_3__5_/chanx_left_out[16] sb_3__5_/chanx_left_out[17] sb_3__5_/chanx_left_out[18]
+ sb_3__5_/chanx_left_out[19] sb_3__5_/chanx_left_out[1] sb_3__5_/chanx_left_out[2]
+ sb_3__5_/chanx_left_out[3] sb_3__5_/chanx_left_out[4] sb_3__5_/chanx_left_out[5]
+ sb_3__5_/chanx_left_out[6] sb_3__5_/chanx_left_out[7] sb_3__5_/chanx_left_out[8]
+ sb_3__5_/chanx_left_out[9] sb_3__5_/chanx_left_in[0] sb_3__5_/chanx_left_in[10]
+ sb_3__5_/chanx_left_in[11] sb_3__5_/chanx_left_in[12] sb_3__5_/chanx_left_in[13]
+ sb_3__5_/chanx_left_in[14] sb_3__5_/chanx_left_in[15] sb_3__5_/chanx_left_in[16]
+ sb_3__5_/chanx_left_in[17] sb_3__5_/chanx_left_in[18] sb_3__5_/chanx_left_in[19]
+ sb_3__5_/chanx_left_in[1] sb_3__5_/chanx_left_in[2] sb_3__5_/chanx_left_in[3] sb_3__5_/chanx_left_in[4]
+ sb_3__5_/chanx_left_in[5] sb_3__5_/chanx_left_in[6] sb_3__5_/chanx_left_in[7] sb_3__5_/chanx_left_in[8]
+ sb_3__5_/chanx_left_in[9] cbx_3__5_/clk_1_N_out cbx_3__5_/clk_1_S_out sb_3__5_/clk_1_W_out
+ cbx_3__5_/clk_2_E_out cbx_3__5_/clk_2_W_in cbx_3__5_/clk_2_W_out cbx_3__5_/clk_3_E_out
+ cbx_3__5_/clk_3_W_in cbx_3__5_/clk_3_W_out cbx_3__5_/prog_clk_0_N_in cbx_3__5_/prog_clk_0_W_out
+ cbx_3__5_/prog_clk_1_N_out cbx_3__5_/prog_clk_1_S_out sb_3__5_/prog_clk_1_W_out
+ cbx_3__5_/prog_clk_2_E_out cbx_3__5_/prog_clk_2_W_in cbx_3__5_/prog_clk_2_W_out
+ cbx_3__5_/prog_clk_3_E_out cbx_3__5_/prog_clk_3_W_in cbx_3__5_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_0__1_ IO_ISOL_N VGND VPWR sb_0__1_/ccff_tail cby_0__1_/ccff_tail sb_0__0_/chany_top_out[0]
+ sb_0__0_/chany_top_out[10] sb_0__0_/chany_top_out[11] sb_0__0_/chany_top_out[12]
+ sb_0__0_/chany_top_out[13] sb_0__0_/chany_top_out[14] sb_0__0_/chany_top_out[15]
+ sb_0__0_/chany_top_out[16] sb_0__0_/chany_top_out[17] sb_0__0_/chany_top_out[18]
+ sb_0__0_/chany_top_out[19] sb_0__0_/chany_top_out[1] sb_0__0_/chany_top_out[2] sb_0__0_/chany_top_out[3]
+ sb_0__0_/chany_top_out[4] sb_0__0_/chany_top_out[5] sb_0__0_/chany_top_out[6] sb_0__0_/chany_top_out[7]
+ sb_0__0_/chany_top_out[8] sb_0__0_/chany_top_out[9] sb_0__0_/chany_top_in[0] sb_0__0_/chany_top_in[10]
+ sb_0__0_/chany_top_in[11] sb_0__0_/chany_top_in[12] sb_0__0_/chany_top_in[13] sb_0__0_/chany_top_in[14]
+ sb_0__0_/chany_top_in[15] sb_0__0_/chany_top_in[16] sb_0__0_/chany_top_in[17] sb_0__0_/chany_top_in[18]
+ sb_0__0_/chany_top_in[19] sb_0__0_/chany_top_in[1] sb_0__0_/chany_top_in[2] sb_0__0_/chany_top_in[3]
+ sb_0__0_/chany_top_in[4] sb_0__0_/chany_top_in[5] sb_0__0_/chany_top_in[6] sb_0__0_/chany_top_in[7]
+ sb_0__0_/chany_top_in[8] sb_0__0_/chany_top_in[9] cby_0__1_/chany_top_in[0] cby_0__1_/chany_top_in[10]
+ cby_0__1_/chany_top_in[11] cby_0__1_/chany_top_in[12] cby_0__1_/chany_top_in[13]
+ cby_0__1_/chany_top_in[14] cby_0__1_/chany_top_in[15] cby_0__1_/chany_top_in[16]
+ cby_0__1_/chany_top_in[17] cby_0__1_/chany_top_in[18] cby_0__1_/chany_top_in[19]
+ cby_0__1_/chany_top_in[1] cby_0__1_/chany_top_in[2] cby_0__1_/chany_top_in[3] cby_0__1_/chany_top_in[4]
+ cby_0__1_/chany_top_in[5] cby_0__1_/chany_top_in[6] cby_0__1_/chany_top_in[7] cby_0__1_/chany_top_in[8]
+ cby_0__1_/chany_top_in[9] cby_0__1_/chany_top_out[0] cby_0__1_/chany_top_out[10]
+ cby_0__1_/chany_top_out[11] cby_0__1_/chany_top_out[12] cby_0__1_/chany_top_out[13]
+ cby_0__1_/chany_top_out[14] cby_0__1_/chany_top_out[15] cby_0__1_/chany_top_out[16]
+ cby_0__1_/chany_top_out[17] cby_0__1_/chany_top_out[18] cby_0__1_/chany_top_out[19]
+ cby_0__1_/chany_top_out[1] cby_0__1_/chany_top_out[2] cby_0__1_/chany_top_out[3]
+ cby_0__1_/chany_top_out[4] cby_0__1_/chany_top_out[5] cby_0__1_/chany_top_out[6]
+ cby_0__1_/chany_top_out[7] cby_0__1_/chany_top_out[8] cby_0__1_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
+ cby_0__1_/left_grid_pin_0_ cby_0__1_/prog_clk_0_E_in cby_0__1_/left_grid_pin_0_
+ sb_0__0_/top_left_grid_pin_1_ sb_0__1_/bottom_left_grid_pin_1_ cby_0__1_
Xsb_7__2_ sb_7__2_/Test_en_N_out sb_7__2_/Test_en_S_in VGND VPWR sb_7__2_/bottom_left_grid_pin_42_
+ sb_7__2_/bottom_left_grid_pin_43_ sb_7__2_/bottom_left_grid_pin_44_ sb_7__2_/bottom_left_grid_pin_45_
+ sb_7__2_/bottom_left_grid_pin_46_ sb_7__2_/bottom_left_grid_pin_47_ sb_7__2_/bottom_left_grid_pin_48_
+ sb_7__2_/bottom_left_grid_pin_49_ sb_7__2_/ccff_head sb_7__2_/ccff_tail sb_7__2_/chanx_left_in[0]
+ sb_7__2_/chanx_left_in[10] sb_7__2_/chanx_left_in[11] sb_7__2_/chanx_left_in[12]
+ sb_7__2_/chanx_left_in[13] sb_7__2_/chanx_left_in[14] sb_7__2_/chanx_left_in[15]
+ sb_7__2_/chanx_left_in[16] sb_7__2_/chanx_left_in[17] sb_7__2_/chanx_left_in[18]
+ sb_7__2_/chanx_left_in[19] sb_7__2_/chanx_left_in[1] sb_7__2_/chanx_left_in[2] sb_7__2_/chanx_left_in[3]
+ sb_7__2_/chanx_left_in[4] sb_7__2_/chanx_left_in[5] sb_7__2_/chanx_left_in[6] sb_7__2_/chanx_left_in[7]
+ sb_7__2_/chanx_left_in[8] sb_7__2_/chanx_left_in[9] sb_7__2_/chanx_left_out[0] sb_7__2_/chanx_left_out[10]
+ sb_7__2_/chanx_left_out[11] sb_7__2_/chanx_left_out[12] sb_7__2_/chanx_left_out[13]
+ sb_7__2_/chanx_left_out[14] sb_7__2_/chanx_left_out[15] sb_7__2_/chanx_left_out[16]
+ sb_7__2_/chanx_left_out[17] sb_7__2_/chanx_left_out[18] sb_7__2_/chanx_left_out[19]
+ sb_7__2_/chanx_left_out[1] sb_7__2_/chanx_left_out[2] sb_7__2_/chanx_left_out[3]
+ sb_7__2_/chanx_left_out[4] sb_7__2_/chanx_left_out[5] sb_7__2_/chanx_left_out[6]
+ sb_7__2_/chanx_left_out[7] sb_7__2_/chanx_left_out[8] sb_7__2_/chanx_left_out[9]
+ sb_7__2_/chanx_right_in[0] sb_7__2_/chanx_right_in[10] sb_7__2_/chanx_right_in[11]
+ sb_7__2_/chanx_right_in[12] sb_7__2_/chanx_right_in[13] sb_7__2_/chanx_right_in[14]
+ sb_7__2_/chanx_right_in[15] sb_7__2_/chanx_right_in[16] sb_7__2_/chanx_right_in[17]
+ sb_7__2_/chanx_right_in[18] sb_7__2_/chanx_right_in[19] sb_7__2_/chanx_right_in[1]
+ sb_7__2_/chanx_right_in[2] sb_7__2_/chanx_right_in[3] sb_7__2_/chanx_right_in[4]
+ sb_7__2_/chanx_right_in[5] sb_7__2_/chanx_right_in[6] sb_7__2_/chanx_right_in[7]
+ sb_7__2_/chanx_right_in[8] sb_7__2_/chanx_right_in[9] cbx_8__2_/chanx_left_in[0]
+ cbx_8__2_/chanx_left_in[10] cbx_8__2_/chanx_left_in[11] cbx_8__2_/chanx_left_in[12]
+ cbx_8__2_/chanx_left_in[13] cbx_8__2_/chanx_left_in[14] cbx_8__2_/chanx_left_in[15]
+ cbx_8__2_/chanx_left_in[16] cbx_8__2_/chanx_left_in[17] cbx_8__2_/chanx_left_in[18]
+ cbx_8__2_/chanx_left_in[19] cbx_8__2_/chanx_left_in[1] cbx_8__2_/chanx_left_in[2]
+ cbx_8__2_/chanx_left_in[3] cbx_8__2_/chanx_left_in[4] cbx_8__2_/chanx_left_in[5]
+ cbx_8__2_/chanx_left_in[6] cbx_8__2_/chanx_left_in[7] cbx_8__2_/chanx_left_in[8]
+ cbx_8__2_/chanx_left_in[9] cby_7__2_/chany_top_out[0] cby_7__2_/chany_top_out[10]
+ cby_7__2_/chany_top_out[11] cby_7__2_/chany_top_out[12] cby_7__2_/chany_top_out[13]
+ cby_7__2_/chany_top_out[14] cby_7__2_/chany_top_out[15] cby_7__2_/chany_top_out[16]
+ cby_7__2_/chany_top_out[17] cby_7__2_/chany_top_out[18] cby_7__2_/chany_top_out[19]
+ cby_7__2_/chany_top_out[1] cby_7__2_/chany_top_out[2] cby_7__2_/chany_top_out[3]
+ cby_7__2_/chany_top_out[4] cby_7__2_/chany_top_out[5] cby_7__2_/chany_top_out[6]
+ cby_7__2_/chany_top_out[7] cby_7__2_/chany_top_out[8] cby_7__2_/chany_top_out[9]
+ cby_7__2_/chany_top_in[0] cby_7__2_/chany_top_in[10] cby_7__2_/chany_top_in[11]
+ cby_7__2_/chany_top_in[12] cby_7__2_/chany_top_in[13] cby_7__2_/chany_top_in[14]
+ cby_7__2_/chany_top_in[15] cby_7__2_/chany_top_in[16] cby_7__2_/chany_top_in[17]
+ cby_7__2_/chany_top_in[18] cby_7__2_/chany_top_in[19] cby_7__2_/chany_top_in[1]
+ cby_7__2_/chany_top_in[2] cby_7__2_/chany_top_in[3] cby_7__2_/chany_top_in[4] cby_7__2_/chany_top_in[5]
+ cby_7__2_/chany_top_in[6] cby_7__2_/chany_top_in[7] cby_7__2_/chany_top_in[8] cby_7__2_/chany_top_in[9]
+ sb_7__2_/chany_top_in[0] sb_7__2_/chany_top_in[10] sb_7__2_/chany_top_in[11] sb_7__2_/chany_top_in[12]
+ sb_7__2_/chany_top_in[13] sb_7__2_/chany_top_in[14] sb_7__2_/chany_top_in[15] sb_7__2_/chany_top_in[16]
+ sb_7__2_/chany_top_in[17] sb_7__2_/chany_top_in[18] sb_7__2_/chany_top_in[19] sb_7__2_/chany_top_in[1]
+ sb_7__2_/chany_top_in[2] sb_7__2_/chany_top_in[3] sb_7__2_/chany_top_in[4] sb_7__2_/chany_top_in[5]
+ sb_7__2_/chany_top_in[6] sb_7__2_/chany_top_in[7] sb_7__2_/chany_top_in[8] sb_7__2_/chany_top_in[9]
+ sb_7__2_/chany_top_out[0] sb_7__2_/chany_top_out[10] sb_7__2_/chany_top_out[11]
+ sb_7__2_/chany_top_out[12] sb_7__2_/chany_top_out[13] sb_7__2_/chany_top_out[14]
+ sb_7__2_/chany_top_out[15] sb_7__2_/chany_top_out[16] sb_7__2_/chany_top_out[17]
+ sb_7__2_/chany_top_out[18] sb_7__2_/chany_top_out[19] sb_7__2_/chany_top_out[1]
+ sb_7__2_/chany_top_out[2] sb_7__2_/chany_top_out[3] sb_7__2_/chany_top_out[4] sb_7__2_/chany_top_out[5]
+ sb_7__2_/chany_top_out[6] sb_7__2_/chany_top_out[7] sb_7__2_/chany_top_out[8] sb_7__2_/chany_top_out[9]
+ sb_7__2_/clk_1_E_out sb_7__2_/clk_1_N_in sb_7__2_/clk_1_W_out sb_7__2_/clk_2_E_out
+ sb_7__2_/clk_2_N_in sb_7__2_/clk_2_N_out sb_7__2_/clk_2_S_out sb_7__2_/clk_2_W_out
+ sb_7__2_/clk_3_E_out sb_7__2_/clk_3_N_in sb_7__2_/clk_3_N_out sb_7__2_/clk_3_S_out
+ sb_7__2_/clk_3_W_out sb_7__2_/left_bottom_grid_pin_34_ sb_7__2_/left_bottom_grid_pin_35_
+ sb_7__2_/left_bottom_grid_pin_36_ sb_7__2_/left_bottom_grid_pin_37_ sb_7__2_/left_bottom_grid_pin_38_
+ sb_7__2_/left_bottom_grid_pin_39_ sb_7__2_/left_bottom_grid_pin_40_ sb_7__2_/left_bottom_grid_pin_41_
+ sb_7__2_/prog_clk_0_N_in sb_7__2_/prog_clk_1_E_out sb_7__2_/prog_clk_1_N_in sb_7__2_/prog_clk_1_W_out
+ sb_7__2_/prog_clk_2_E_out sb_7__2_/prog_clk_2_N_in sb_7__2_/prog_clk_2_N_out sb_7__2_/prog_clk_2_S_out
+ sb_7__2_/prog_clk_2_W_out sb_7__2_/prog_clk_3_E_out sb_7__2_/prog_clk_3_N_in sb_7__2_/prog_clk_3_N_out
+ sb_7__2_/prog_clk_3_S_out sb_7__2_/prog_clk_3_W_out sb_7__2_/right_bottom_grid_pin_34_
+ sb_7__2_/right_bottom_grid_pin_35_ sb_7__2_/right_bottom_grid_pin_36_ sb_7__2_/right_bottom_grid_pin_37_
+ sb_7__2_/right_bottom_grid_pin_38_ sb_7__2_/right_bottom_grid_pin_39_ sb_7__2_/right_bottom_grid_pin_40_
+ sb_7__2_/right_bottom_grid_pin_41_ sb_7__2_/top_left_grid_pin_42_ sb_7__2_/top_left_grid_pin_43_
+ sb_7__2_/top_left_grid_pin_44_ sb_7__2_/top_left_grid_pin_45_ sb_7__2_/top_left_grid_pin_46_
+ sb_7__2_/top_left_grid_pin_47_ sb_7__2_/top_left_grid_pin_48_ sb_7__2_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_0__7_ VGND VPWR sb_0__7_/bottom_left_grid_pin_1_ sb_0__7_/ccff_head sb_0__7_/ccff_tail
+ sb_0__7_/chanx_right_in[0] sb_0__7_/chanx_right_in[10] sb_0__7_/chanx_right_in[11]
+ sb_0__7_/chanx_right_in[12] sb_0__7_/chanx_right_in[13] sb_0__7_/chanx_right_in[14]
+ sb_0__7_/chanx_right_in[15] sb_0__7_/chanx_right_in[16] sb_0__7_/chanx_right_in[17]
+ sb_0__7_/chanx_right_in[18] sb_0__7_/chanx_right_in[19] sb_0__7_/chanx_right_in[1]
+ sb_0__7_/chanx_right_in[2] sb_0__7_/chanx_right_in[3] sb_0__7_/chanx_right_in[4]
+ sb_0__7_/chanx_right_in[5] sb_0__7_/chanx_right_in[6] sb_0__7_/chanx_right_in[7]
+ sb_0__7_/chanx_right_in[8] sb_0__7_/chanx_right_in[9] cbx_1__7_/chanx_left_in[0]
+ cbx_1__7_/chanx_left_in[10] cbx_1__7_/chanx_left_in[11] cbx_1__7_/chanx_left_in[12]
+ cbx_1__7_/chanx_left_in[13] cbx_1__7_/chanx_left_in[14] cbx_1__7_/chanx_left_in[15]
+ cbx_1__7_/chanx_left_in[16] cbx_1__7_/chanx_left_in[17] cbx_1__7_/chanx_left_in[18]
+ cbx_1__7_/chanx_left_in[19] cbx_1__7_/chanx_left_in[1] cbx_1__7_/chanx_left_in[2]
+ cbx_1__7_/chanx_left_in[3] cbx_1__7_/chanx_left_in[4] cbx_1__7_/chanx_left_in[5]
+ cbx_1__7_/chanx_left_in[6] cbx_1__7_/chanx_left_in[7] cbx_1__7_/chanx_left_in[8]
+ cbx_1__7_/chanx_left_in[9] cby_0__7_/chany_top_out[0] cby_0__7_/chany_top_out[10]
+ cby_0__7_/chany_top_out[11] cby_0__7_/chany_top_out[12] cby_0__7_/chany_top_out[13]
+ cby_0__7_/chany_top_out[14] cby_0__7_/chany_top_out[15] cby_0__7_/chany_top_out[16]
+ cby_0__7_/chany_top_out[17] cby_0__7_/chany_top_out[18] cby_0__7_/chany_top_out[19]
+ cby_0__7_/chany_top_out[1] cby_0__7_/chany_top_out[2] cby_0__7_/chany_top_out[3]
+ cby_0__7_/chany_top_out[4] cby_0__7_/chany_top_out[5] cby_0__7_/chany_top_out[6]
+ cby_0__7_/chany_top_out[7] cby_0__7_/chany_top_out[8] cby_0__7_/chany_top_out[9]
+ cby_0__7_/chany_top_in[0] cby_0__7_/chany_top_in[10] cby_0__7_/chany_top_in[11]
+ cby_0__7_/chany_top_in[12] cby_0__7_/chany_top_in[13] cby_0__7_/chany_top_in[14]
+ cby_0__7_/chany_top_in[15] cby_0__7_/chany_top_in[16] cby_0__7_/chany_top_in[17]
+ cby_0__7_/chany_top_in[18] cby_0__7_/chany_top_in[19] cby_0__7_/chany_top_in[1]
+ cby_0__7_/chany_top_in[2] cby_0__7_/chany_top_in[3] cby_0__7_/chany_top_in[4] cby_0__7_/chany_top_in[5]
+ cby_0__7_/chany_top_in[6] cby_0__7_/chany_top_in[7] cby_0__7_/chany_top_in[8] cby_0__7_/chany_top_in[9]
+ sb_0__7_/chany_top_in[0] sb_0__7_/chany_top_in[10] sb_0__7_/chany_top_in[11] sb_0__7_/chany_top_in[12]
+ sb_0__7_/chany_top_in[13] sb_0__7_/chany_top_in[14] sb_0__7_/chany_top_in[15] sb_0__7_/chany_top_in[16]
+ sb_0__7_/chany_top_in[17] sb_0__7_/chany_top_in[18] sb_0__7_/chany_top_in[19] sb_0__7_/chany_top_in[1]
+ sb_0__7_/chany_top_in[2] sb_0__7_/chany_top_in[3] sb_0__7_/chany_top_in[4] sb_0__7_/chany_top_in[5]
+ sb_0__7_/chany_top_in[6] sb_0__7_/chany_top_in[7] sb_0__7_/chany_top_in[8] sb_0__7_/chany_top_in[9]
+ sb_0__7_/chany_top_out[0] sb_0__7_/chany_top_out[10] sb_0__7_/chany_top_out[11]
+ sb_0__7_/chany_top_out[12] sb_0__7_/chany_top_out[13] sb_0__7_/chany_top_out[14]
+ sb_0__7_/chany_top_out[15] sb_0__7_/chany_top_out[16] sb_0__7_/chany_top_out[17]
+ sb_0__7_/chany_top_out[18] sb_0__7_/chany_top_out[19] sb_0__7_/chany_top_out[1]
+ sb_0__7_/chany_top_out[2] sb_0__7_/chany_top_out[3] sb_0__7_/chany_top_out[4] sb_0__7_/chany_top_out[5]
+ sb_0__7_/chany_top_out[6] sb_0__7_/chany_top_out[7] sb_0__7_/chany_top_out[8] sb_0__7_/chany_top_out[9]
+ sb_0__7_/prog_clk_0_E_in sb_0__7_/right_bottom_grid_pin_34_ sb_0__7_/right_bottom_grid_pin_35_
+ sb_0__7_/right_bottom_grid_pin_36_ sb_0__7_/right_bottom_grid_pin_37_ sb_0__7_/right_bottom_grid_pin_38_
+ sb_0__7_/right_bottom_grid_pin_39_ sb_0__7_/right_bottom_grid_pin_40_ sb_0__7_/right_bottom_grid_pin_41_
+ sb_0__7_/top_left_grid_pin_1_ sb_0__1_
Xgrid_clb_2__5_ cbx_2__4_/SC_OUT_TOP grid_clb_2__5_/SC_OUT_BOT cbx_2__5_/SC_IN_BOT
+ cby_2__5_/Test_en_W_out grid_clb_2__5_/Test_en_E_out cby_2__5_/Test_en_W_out cby_1__5_/Test_en_W_in
+ VGND VPWR cbx_2__4_/REGIN_FEEDTHROUGH grid_clb_2__5_/bottom_width_0_height_0__pin_51_
+ cby_1__5_/ccff_tail cby_2__5_/ccff_head cbx_2__5_/clk_1_S_out cbx_2__5_/clk_1_S_out
+ cby_2__5_/prog_clk_0_W_in cbx_2__5_/prog_clk_1_S_out grid_clb_2__5_/prog_clk_0_N_out
+ cbx_2__5_/prog_clk_1_S_out cbx_2__4_/prog_clk_0_N_in grid_clb_2__5_/prog_clk_0_W_out
+ cby_2__5_/left_grid_pin_16_ cby_2__5_/left_grid_pin_17_ cby_2__5_/left_grid_pin_18_
+ cby_2__5_/left_grid_pin_19_ cby_2__5_/left_grid_pin_20_ cby_2__5_/left_grid_pin_21_
+ cby_2__5_/left_grid_pin_22_ cby_2__5_/left_grid_pin_23_ cby_2__5_/left_grid_pin_24_
+ cby_2__5_/left_grid_pin_25_ cby_2__5_/left_grid_pin_26_ cby_2__5_/left_grid_pin_27_
+ cby_2__5_/left_grid_pin_28_ cby_2__5_/left_grid_pin_29_ cby_2__5_/left_grid_pin_30_
+ cby_2__5_/left_grid_pin_31_ sb_2__4_/top_left_grid_pin_42_ sb_2__5_/bottom_left_grid_pin_42_
+ sb_2__4_/top_left_grid_pin_43_ sb_2__5_/bottom_left_grid_pin_43_ sb_2__4_/top_left_grid_pin_44_
+ sb_2__5_/bottom_left_grid_pin_44_ sb_2__4_/top_left_grid_pin_45_ sb_2__5_/bottom_left_grid_pin_45_
+ sb_2__4_/top_left_grid_pin_46_ sb_2__5_/bottom_left_grid_pin_46_ sb_2__4_/top_left_grid_pin_47_
+ sb_2__5_/bottom_left_grid_pin_47_ sb_2__4_/top_left_grid_pin_48_ sb_2__5_/bottom_left_grid_pin_48_
+ sb_2__4_/top_left_grid_pin_49_ sb_2__5_/bottom_left_grid_pin_49_ cbx_2__5_/bottom_grid_pin_0_
+ cbx_2__5_/bottom_grid_pin_10_ cbx_2__5_/bottom_grid_pin_11_ cbx_2__5_/bottom_grid_pin_12_
+ cbx_2__5_/bottom_grid_pin_13_ cbx_2__5_/bottom_grid_pin_14_ cbx_2__5_/bottom_grid_pin_15_
+ cbx_2__5_/bottom_grid_pin_1_ cbx_2__5_/bottom_grid_pin_2_ cbx_2__5_/REGOUT_FEEDTHROUGH
+ grid_clb_2__5_/top_width_0_height_0__pin_33_ sb_2__5_/left_bottom_grid_pin_34_ sb_1__5_/right_bottom_grid_pin_34_
+ sb_2__5_/left_bottom_grid_pin_35_ sb_1__5_/right_bottom_grid_pin_35_ sb_2__5_/left_bottom_grid_pin_36_
+ sb_1__5_/right_bottom_grid_pin_36_ sb_2__5_/left_bottom_grid_pin_37_ sb_1__5_/right_bottom_grid_pin_37_
+ sb_2__5_/left_bottom_grid_pin_38_ sb_1__5_/right_bottom_grid_pin_38_ sb_2__5_/left_bottom_grid_pin_39_
+ sb_1__5_/right_bottom_grid_pin_39_ cbx_2__5_/bottom_grid_pin_3_ sb_2__5_/left_bottom_grid_pin_40_
+ sb_1__5_/right_bottom_grid_pin_40_ sb_2__5_/left_bottom_grid_pin_41_ sb_1__5_/right_bottom_grid_pin_41_
+ cbx_2__5_/bottom_grid_pin_4_ cbx_2__5_/bottom_grid_pin_5_ cbx_2__5_/bottom_grid_pin_6_
+ cbx_2__5_/bottom_grid_pin_7_ cbx_2__5_/bottom_grid_pin_8_ cbx_2__5_/bottom_grid_pin_9_
+ grid_clb
Xcby_6__6_ cby_6__6_/Test_en_W_in cby_6__6_/Test_en_E_out cby_6__6_/Test_en_N_out
+ cby_6__6_/Test_en_W_in cby_6__6_/Test_en_W_in cby_6__6_/Test_en_W_out VGND VPWR
+ cby_6__6_/ccff_head cby_6__6_/ccff_tail sb_6__5_/chany_top_out[0] sb_6__5_/chany_top_out[10]
+ sb_6__5_/chany_top_out[11] sb_6__5_/chany_top_out[12] sb_6__5_/chany_top_out[13]
+ sb_6__5_/chany_top_out[14] sb_6__5_/chany_top_out[15] sb_6__5_/chany_top_out[16]
+ sb_6__5_/chany_top_out[17] sb_6__5_/chany_top_out[18] sb_6__5_/chany_top_out[19]
+ sb_6__5_/chany_top_out[1] sb_6__5_/chany_top_out[2] sb_6__5_/chany_top_out[3] sb_6__5_/chany_top_out[4]
+ sb_6__5_/chany_top_out[5] sb_6__5_/chany_top_out[6] sb_6__5_/chany_top_out[7] sb_6__5_/chany_top_out[8]
+ sb_6__5_/chany_top_out[9] sb_6__5_/chany_top_in[0] sb_6__5_/chany_top_in[10] sb_6__5_/chany_top_in[11]
+ sb_6__5_/chany_top_in[12] sb_6__5_/chany_top_in[13] sb_6__5_/chany_top_in[14] sb_6__5_/chany_top_in[15]
+ sb_6__5_/chany_top_in[16] sb_6__5_/chany_top_in[17] sb_6__5_/chany_top_in[18] sb_6__5_/chany_top_in[19]
+ sb_6__5_/chany_top_in[1] sb_6__5_/chany_top_in[2] sb_6__5_/chany_top_in[3] sb_6__5_/chany_top_in[4]
+ sb_6__5_/chany_top_in[5] sb_6__5_/chany_top_in[6] sb_6__5_/chany_top_in[7] sb_6__5_/chany_top_in[8]
+ sb_6__5_/chany_top_in[9] cby_6__6_/chany_top_in[0] cby_6__6_/chany_top_in[10] cby_6__6_/chany_top_in[11]
+ cby_6__6_/chany_top_in[12] cby_6__6_/chany_top_in[13] cby_6__6_/chany_top_in[14]
+ cby_6__6_/chany_top_in[15] cby_6__6_/chany_top_in[16] cby_6__6_/chany_top_in[17]
+ cby_6__6_/chany_top_in[18] cby_6__6_/chany_top_in[19] cby_6__6_/chany_top_in[1]
+ cby_6__6_/chany_top_in[2] cby_6__6_/chany_top_in[3] cby_6__6_/chany_top_in[4] cby_6__6_/chany_top_in[5]
+ cby_6__6_/chany_top_in[6] cby_6__6_/chany_top_in[7] cby_6__6_/chany_top_in[8] cby_6__6_/chany_top_in[9]
+ cby_6__6_/chany_top_out[0] cby_6__6_/chany_top_out[10] cby_6__6_/chany_top_out[11]
+ cby_6__6_/chany_top_out[12] cby_6__6_/chany_top_out[13] cby_6__6_/chany_top_out[14]
+ cby_6__6_/chany_top_out[15] cby_6__6_/chany_top_out[16] cby_6__6_/chany_top_out[17]
+ cby_6__6_/chany_top_out[18] cby_6__6_/chany_top_out[19] cby_6__6_/chany_top_out[1]
+ cby_6__6_/chany_top_out[2] cby_6__6_/chany_top_out[3] cby_6__6_/chany_top_out[4]
+ cby_6__6_/chany_top_out[5] cby_6__6_/chany_top_out[6] cby_6__6_/chany_top_out[7]
+ cby_6__6_/chany_top_out[8] cby_6__6_/chany_top_out[9] cby_6__6_/clk_2_N_out cby_6__6_/clk_2_S_in
+ cby_6__6_/clk_2_S_out sb_6__6_/clk_2_N_in sb_6__5_/clk_3_N_out cby_6__6_/clk_3_S_out
+ cby_6__6_/left_grid_pin_16_ cby_6__6_/left_grid_pin_17_ cby_6__6_/left_grid_pin_18_
+ cby_6__6_/left_grid_pin_19_ cby_6__6_/left_grid_pin_20_ cby_6__6_/left_grid_pin_21_
+ cby_6__6_/left_grid_pin_22_ cby_6__6_/left_grid_pin_23_ cby_6__6_/left_grid_pin_24_
+ cby_6__6_/left_grid_pin_25_ cby_6__6_/left_grid_pin_26_ cby_6__6_/left_grid_pin_27_
+ cby_6__6_/left_grid_pin_28_ cby_6__6_/left_grid_pin_29_ cby_6__6_/left_grid_pin_30_
+ cby_6__6_/left_grid_pin_31_ cby_6__6_/prog_clk_0_N_out sb_6__5_/prog_clk_0_N_in
+ cby_6__6_/prog_clk_0_W_in cby_6__6_/prog_clk_2_N_out cby_6__6_/prog_clk_2_S_in cby_6__6_/prog_clk_2_S_out
+ sb_6__6_/prog_clk_2_N_in sb_6__5_/prog_clk_3_N_out cby_6__6_/prog_clk_3_S_out cby_1__1_
Xcbx_6__7_ cbx_6__7_/REGIN_FEEDTHROUGH cbx_6__7_/REGOUT_FEEDTHROUGH cbx_6__7_/SC_IN_BOT
+ cbx_6__7_/SC_IN_TOP cbx_6__7_/SC_OUT_BOT cbx_6__7_/SC_OUT_TOP VGND VPWR cbx_6__7_/bottom_grid_pin_0_
+ cbx_6__7_/bottom_grid_pin_10_ cbx_6__7_/bottom_grid_pin_11_ cbx_6__7_/bottom_grid_pin_12_
+ cbx_6__7_/bottom_grid_pin_13_ cbx_6__7_/bottom_grid_pin_14_ cbx_6__7_/bottom_grid_pin_15_
+ cbx_6__7_/bottom_grid_pin_1_ cbx_6__7_/bottom_grid_pin_2_ cbx_6__7_/bottom_grid_pin_3_
+ cbx_6__7_/bottom_grid_pin_4_ cbx_6__7_/bottom_grid_pin_5_ cbx_6__7_/bottom_grid_pin_6_
+ cbx_6__7_/bottom_grid_pin_7_ cbx_6__7_/bottom_grid_pin_8_ cbx_6__7_/bottom_grid_pin_9_
+ sb_6__7_/ccff_tail sb_5__7_/ccff_head cbx_6__7_/chanx_left_in[0] cbx_6__7_/chanx_left_in[10]
+ cbx_6__7_/chanx_left_in[11] cbx_6__7_/chanx_left_in[12] cbx_6__7_/chanx_left_in[13]
+ cbx_6__7_/chanx_left_in[14] cbx_6__7_/chanx_left_in[15] cbx_6__7_/chanx_left_in[16]
+ cbx_6__7_/chanx_left_in[17] cbx_6__7_/chanx_left_in[18] cbx_6__7_/chanx_left_in[19]
+ cbx_6__7_/chanx_left_in[1] cbx_6__7_/chanx_left_in[2] cbx_6__7_/chanx_left_in[3]
+ cbx_6__7_/chanx_left_in[4] cbx_6__7_/chanx_left_in[5] cbx_6__7_/chanx_left_in[6]
+ cbx_6__7_/chanx_left_in[7] cbx_6__7_/chanx_left_in[8] cbx_6__7_/chanx_left_in[9]
+ sb_5__7_/chanx_right_in[0] sb_5__7_/chanx_right_in[10] sb_5__7_/chanx_right_in[11]
+ sb_5__7_/chanx_right_in[12] sb_5__7_/chanx_right_in[13] sb_5__7_/chanx_right_in[14]
+ sb_5__7_/chanx_right_in[15] sb_5__7_/chanx_right_in[16] sb_5__7_/chanx_right_in[17]
+ sb_5__7_/chanx_right_in[18] sb_5__7_/chanx_right_in[19] sb_5__7_/chanx_right_in[1]
+ sb_5__7_/chanx_right_in[2] sb_5__7_/chanx_right_in[3] sb_5__7_/chanx_right_in[4]
+ sb_5__7_/chanx_right_in[5] sb_5__7_/chanx_right_in[6] sb_5__7_/chanx_right_in[7]
+ sb_5__7_/chanx_right_in[8] sb_5__7_/chanx_right_in[9] sb_6__7_/chanx_left_out[0]
+ sb_6__7_/chanx_left_out[10] sb_6__7_/chanx_left_out[11] sb_6__7_/chanx_left_out[12]
+ sb_6__7_/chanx_left_out[13] sb_6__7_/chanx_left_out[14] sb_6__7_/chanx_left_out[15]
+ sb_6__7_/chanx_left_out[16] sb_6__7_/chanx_left_out[17] sb_6__7_/chanx_left_out[18]
+ sb_6__7_/chanx_left_out[19] sb_6__7_/chanx_left_out[1] sb_6__7_/chanx_left_out[2]
+ sb_6__7_/chanx_left_out[3] sb_6__7_/chanx_left_out[4] sb_6__7_/chanx_left_out[5]
+ sb_6__7_/chanx_left_out[6] sb_6__7_/chanx_left_out[7] sb_6__7_/chanx_left_out[8]
+ sb_6__7_/chanx_left_out[9] sb_6__7_/chanx_left_in[0] sb_6__7_/chanx_left_in[10]
+ sb_6__7_/chanx_left_in[11] sb_6__7_/chanx_left_in[12] sb_6__7_/chanx_left_in[13]
+ sb_6__7_/chanx_left_in[14] sb_6__7_/chanx_left_in[15] sb_6__7_/chanx_left_in[16]
+ sb_6__7_/chanx_left_in[17] sb_6__7_/chanx_left_in[18] sb_6__7_/chanx_left_in[19]
+ sb_6__7_/chanx_left_in[1] sb_6__7_/chanx_left_in[2] sb_6__7_/chanx_left_in[3] sb_6__7_/chanx_left_in[4]
+ sb_6__7_/chanx_left_in[5] sb_6__7_/chanx_left_in[6] sb_6__7_/chanx_left_in[7] sb_6__7_/chanx_left_in[8]
+ sb_6__7_/chanx_left_in[9] cbx_6__7_/clk_1_N_out cbx_6__7_/clk_1_S_out sb_5__7_/clk_1_E_out
+ cbx_6__7_/clk_2_E_out cbx_6__7_/clk_2_W_in cbx_6__7_/clk_2_W_out cbx_6__7_/clk_3_E_out
+ cbx_6__7_/clk_3_W_in cbx_6__7_/clk_3_W_out cbx_6__7_/prog_clk_0_N_in cbx_6__7_/prog_clk_0_W_out
+ cbx_6__7_/prog_clk_1_N_out cbx_6__7_/prog_clk_1_S_out sb_5__7_/prog_clk_1_E_out
+ cbx_6__7_/prog_clk_2_E_out cbx_6__7_/prog_clk_2_W_in cbx_6__7_/prog_clk_2_W_out
+ cbx_6__7_/prog_clk_3_E_out cbx_6__7_/prog_clk_3_W_in cbx_6__7_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_3__3_ cby_3__3_/Test_en_W_in cby_3__3_/Test_en_E_out cby_3__3_/Test_en_N_out
+ cby_3__3_/Test_en_W_in cby_3__3_/Test_en_W_in cby_3__3_/Test_en_W_out VGND VPWR
+ cby_3__3_/ccff_head cby_3__3_/ccff_tail sb_3__2_/chany_top_out[0] sb_3__2_/chany_top_out[10]
+ sb_3__2_/chany_top_out[11] sb_3__2_/chany_top_out[12] sb_3__2_/chany_top_out[13]
+ sb_3__2_/chany_top_out[14] sb_3__2_/chany_top_out[15] sb_3__2_/chany_top_out[16]
+ sb_3__2_/chany_top_out[17] sb_3__2_/chany_top_out[18] sb_3__2_/chany_top_out[19]
+ sb_3__2_/chany_top_out[1] sb_3__2_/chany_top_out[2] sb_3__2_/chany_top_out[3] sb_3__2_/chany_top_out[4]
+ sb_3__2_/chany_top_out[5] sb_3__2_/chany_top_out[6] sb_3__2_/chany_top_out[7] sb_3__2_/chany_top_out[8]
+ sb_3__2_/chany_top_out[9] sb_3__2_/chany_top_in[0] sb_3__2_/chany_top_in[10] sb_3__2_/chany_top_in[11]
+ sb_3__2_/chany_top_in[12] sb_3__2_/chany_top_in[13] sb_3__2_/chany_top_in[14] sb_3__2_/chany_top_in[15]
+ sb_3__2_/chany_top_in[16] sb_3__2_/chany_top_in[17] sb_3__2_/chany_top_in[18] sb_3__2_/chany_top_in[19]
+ sb_3__2_/chany_top_in[1] sb_3__2_/chany_top_in[2] sb_3__2_/chany_top_in[3] sb_3__2_/chany_top_in[4]
+ sb_3__2_/chany_top_in[5] sb_3__2_/chany_top_in[6] sb_3__2_/chany_top_in[7] sb_3__2_/chany_top_in[8]
+ sb_3__2_/chany_top_in[9] cby_3__3_/chany_top_in[0] cby_3__3_/chany_top_in[10] cby_3__3_/chany_top_in[11]
+ cby_3__3_/chany_top_in[12] cby_3__3_/chany_top_in[13] cby_3__3_/chany_top_in[14]
+ cby_3__3_/chany_top_in[15] cby_3__3_/chany_top_in[16] cby_3__3_/chany_top_in[17]
+ cby_3__3_/chany_top_in[18] cby_3__3_/chany_top_in[19] cby_3__3_/chany_top_in[1]
+ cby_3__3_/chany_top_in[2] cby_3__3_/chany_top_in[3] cby_3__3_/chany_top_in[4] cby_3__3_/chany_top_in[5]
+ cby_3__3_/chany_top_in[6] cby_3__3_/chany_top_in[7] cby_3__3_/chany_top_in[8] cby_3__3_/chany_top_in[9]
+ cby_3__3_/chany_top_out[0] cby_3__3_/chany_top_out[10] cby_3__3_/chany_top_out[11]
+ cby_3__3_/chany_top_out[12] cby_3__3_/chany_top_out[13] cby_3__3_/chany_top_out[14]
+ cby_3__3_/chany_top_out[15] cby_3__3_/chany_top_out[16] cby_3__3_/chany_top_out[17]
+ cby_3__3_/chany_top_out[18] cby_3__3_/chany_top_out[19] cby_3__3_/chany_top_out[1]
+ cby_3__3_/chany_top_out[2] cby_3__3_/chany_top_out[3] cby_3__3_/chany_top_out[4]
+ cby_3__3_/chany_top_out[5] cby_3__3_/chany_top_out[6] cby_3__3_/chany_top_out[7]
+ cby_3__3_/chany_top_out[8] cby_3__3_/chany_top_out[9] sb_3__3_/clk_1_N_in sb_3__2_/clk_2_N_out
+ cby_3__3_/clk_2_S_out cby_3__3_/clk_3_N_out cby_3__3_/clk_3_S_in cby_3__3_/clk_3_S_out
+ cby_3__3_/left_grid_pin_16_ cby_3__3_/left_grid_pin_17_ cby_3__3_/left_grid_pin_18_
+ cby_3__3_/left_grid_pin_19_ cby_3__3_/left_grid_pin_20_ cby_3__3_/left_grid_pin_21_
+ cby_3__3_/left_grid_pin_22_ cby_3__3_/left_grid_pin_23_ cby_3__3_/left_grid_pin_24_
+ cby_3__3_/left_grid_pin_25_ cby_3__3_/left_grid_pin_26_ cby_3__3_/left_grid_pin_27_
+ cby_3__3_/left_grid_pin_28_ cby_3__3_/left_grid_pin_29_ cby_3__3_/left_grid_pin_30_
+ cby_3__3_/left_grid_pin_31_ cby_3__3_/prog_clk_0_N_out sb_3__2_/prog_clk_0_N_in
+ cby_3__3_/prog_clk_0_W_in sb_3__3_/prog_clk_1_N_in sb_3__2_/prog_clk_2_N_out cby_3__3_/prog_clk_2_S_out
+ cby_3__3_/prog_clk_3_N_out cby_3__3_/prog_clk_3_S_in cby_3__3_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_5__7_ cbx_5__7_/SC_OUT_BOT cbx_5__6_/SC_IN_TOP grid_clb_5__7_/SC_OUT_TOP
+ cby_4__7_/Test_en_E_out cby_5__7_/Test_en_W_in cby_4__7_/Test_en_E_out grid_clb_5__7_/Test_en_W_out
+ VGND VPWR cbx_5__6_/REGIN_FEEDTHROUGH grid_clb_5__7_/bottom_width_0_height_0__pin_51_
+ cby_4__7_/ccff_tail cby_5__7_/ccff_head cbx_5__7_/clk_1_S_out cbx_5__7_/clk_1_S_out
+ cby_5__7_/prog_clk_0_W_in cbx_5__7_/prog_clk_1_S_out grid_clb_5__7_/prog_clk_0_N_out
+ cbx_5__7_/prog_clk_1_S_out cbx_5__6_/prog_clk_0_N_in grid_clb_5__7_/prog_clk_0_W_out
+ cby_5__7_/left_grid_pin_16_ cby_5__7_/left_grid_pin_17_ cby_5__7_/left_grid_pin_18_
+ cby_5__7_/left_grid_pin_19_ cby_5__7_/left_grid_pin_20_ cby_5__7_/left_grid_pin_21_
+ cby_5__7_/left_grid_pin_22_ cby_5__7_/left_grid_pin_23_ cby_5__7_/left_grid_pin_24_
+ cby_5__7_/left_grid_pin_25_ cby_5__7_/left_grid_pin_26_ cby_5__7_/left_grid_pin_27_
+ cby_5__7_/left_grid_pin_28_ cby_5__7_/left_grid_pin_29_ cby_5__7_/left_grid_pin_30_
+ cby_5__7_/left_grid_pin_31_ sb_5__6_/top_left_grid_pin_42_ sb_5__7_/bottom_left_grid_pin_42_
+ sb_5__6_/top_left_grid_pin_43_ sb_5__7_/bottom_left_grid_pin_43_ sb_5__6_/top_left_grid_pin_44_
+ sb_5__7_/bottom_left_grid_pin_44_ sb_5__6_/top_left_grid_pin_45_ sb_5__7_/bottom_left_grid_pin_45_
+ sb_5__6_/top_left_grid_pin_46_ sb_5__7_/bottom_left_grid_pin_46_ sb_5__6_/top_left_grid_pin_47_
+ sb_5__7_/bottom_left_grid_pin_47_ sb_5__6_/top_left_grid_pin_48_ sb_5__7_/bottom_left_grid_pin_48_
+ sb_5__6_/top_left_grid_pin_49_ sb_5__7_/bottom_left_grid_pin_49_ cbx_5__7_/bottom_grid_pin_0_
+ cbx_5__7_/bottom_grid_pin_10_ cbx_5__7_/bottom_grid_pin_11_ cbx_5__7_/bottom_grid_pin_12_
+ cbx_5__7_/bottom_grid_pin_13_ cbx_5__7_/bottom_grid_pin_14_ cbx_5__7_/bottom_grid_pin_15_
+ cbx_5__7_/bottom_grid_pin_1_ cbx_5__7_/bottom_grid_pin_2_ cbx_5__7_/REGOUT_FEEDTHROUGH
+ grid_clb_5__7_/top_width_0_height_0__pin_33_ sb_5__7_/left_bottom_grid_pin_34_ sb_4__7_/right_bottom_grid_pin_34_
+ sb_5__7_/left_bottom_grid_pin_35_ sb_4__7_/right_bottom_grid_pin_35_ sb_5__7_/left_bottom_grid_pin_36_
+ sb_4__7_/right_bottom_grid_pin_36_ sb_5__7_/left_bottom_grid_pin_37_ sb_4__7_/right_bottom_grid_pin_37_
+ sb_5__7_/left_bottom_grid_pin_38_ sb_4__7_/right_bottom_grid_pin_38_ sb_5__7_/left_bottom_grid_pin_39_
+ sb_4__7_/right_bottom_grid_pin_39_ cbx_5__7_/bottom_grid_pin_3_ sb_5__7_/left_bottom_grid_pin_40_
+ sb_4__7_/right_bottom_grid_pin_40_ sb_5__7_/left_bottom_grid_pin_41_ sb_4__7_/right_bottom_grid_pin_41_
+ cbx_5__7_/bottom_grid_pin_4_ cbx_5__7_/bottom_grid_pin_5_ cbx_5__7_/bottom_grid_pin_6_
+ cbx_5__7_/bottom_grid_pin_7_ cbx_5__7_/bottom_grid_pin_8_ cbx_5__7_/bottom_grid_pin_9_
+ grid_clb
Xcbx_3__4_ cbx_3__4_/REGIN_FEEDTHROUGH cbx_3__4_/REGOUT_FEEDTHROUGH cbx_3__4_/SC_IN_BOT
+ cbx_3__4_/SC_IN_TOP cbx_3__4_/SC_OUT_BOT cbx_3__4_/SC_OUT_TOP VGND VPWR cbx_3__4_/bottom_grid_pin_0_
+ cbx_3__4_/bottom_grid_pin_10_ cbx_3__4_/bottom_grid_pin_11_ cbx_3__4_/bottom_grid_pin_12_
+ cbx_3__4_/bottom_grid_pin_13_ cbx_3__4_/bottom_grid_pin_14_ cbx_3__4_/bottom_grid_pin_15_
+ cbx_3__4_/bottom_grid_pin_1_ cbx_3__4_/bottom_grid_pin_2_ cbx_3__4_/bottom_grid_pin_3_
+ cbx_3__4_/bottom_grid_pin_4_ cbx_3__4_/bottom_grid_pin_5_ cbx_3__4_/bottom_grid_pin_6_
+ cbx_3__4_/bottom_grid_pin_7_ cbx_3__4_/bottom_grid_pin_8_ cbx_3__4_/bottom_grid_pin_9_
+ sb_3__4_/ccff_tail sb_2__4_/ccff_head cbx_3__4_/chanx_left_in[0] cbx_3__4_/chanx_left_in[10]
+ cbx_3__4_/chanx_left_in[11] cbx_3__4_/chanx_left_in[12] cbx_3__4_/chanx_left_in[13]
+ cbx_3__4_/chanx_left_in[14] cbx_3__4_/chanx_left_in[15] cbx_3__4_/chanx_left_in[16]
+ cbx_3__4_/chanx_left_in[17] cbx_3__4_/chanx_left_in[18] cbx_3__4_/chanx_left_in[19]
+ cbx_3__4_/chanx_left_in[1] cbx_3__4_/chanx_left_in[2] cbx_3__4_/chanx_left_in[3]
+ cbx_3__4_/chanx_left_in[4] cbx_3__4_/chanx_left_in[5] cbx_3__4_/chanx_left_in[6]
+ cbx_3__4_/chanx_left_in[7] cbx_3__4_/chanx_left_in[8] cbx_3__4_/chanx_left_in[9]
+ sb_2__4_/chanx_right_in[0] sb_2__4_/chanx_right_in[10] sb_2__4_/chanx_right_in[11]
+ sb_2__4_/chanx_right_in[12] sb_2__4_/chanx_right_in[13] sb_2__4_/chanx_right_in[14]
+ sb_2__4_/chanx_right_in[15] sb_2__4_/chanx_right_in[16] sb_2__4_/chanx_right_in[17]
+ sb_2__4_/chanx_right_in[18] sb_2__4_/chanx_right_in[19] sb_2__4_/chanx_right_in[1]
+ sb_2__4_/chanx_right_in[2] sb_2__4_/chanx_right_in[3] sb_2__4_/chanx_right_in[4]
+ sb_2__4_/chanx_right_in[5] sb_2__4_/chanx_right_in[6] sb_2__4_/chanx_right_in[7]
+ sb_2__4_/chanx_right_in[8] sb_2__4_/chanx_right_in[9] sb_3__4_/chanx_left_out[0]
+ sb_3__4_/chanx_left_out[10] sb_3__4_/chanx_left_out[11] sb_3__4_/chanx_left_out[12]
+ sb_3__4_/chanx_left_out[13] sb_3__4_/chanx_left_out[14] sb_3__4_/chanx_left_out[15]
+ sb_3__4_/chanx_left_out[16] sb_3__4_/chanx_left_out[17] sb_3__4_/chanx_left_out[18]
+ sb_3__4_/chanx_left_out[19] sb_3__4_/chanx_left_out[1] sb_3__4_/chanx_left_out[2]
+ sb_3__4_/chanx_left_out[3] sb_3__4_/chanx_left_out[4] sb_3__4_/chanx_left_out[5]
+ sb_3__4_/chanx_left_out[6] sb_3__4_/chanx_left_out[7] sb_3__4_/chanx_left_out[8]
+ sb_3__4_/chanx_left_out[9] sb_3__4_/chanx_left_in[0] sb_3__4_/chanx_left_in[10]
+ sb_3__4_/chanx_left_in[11] sb_3__4_/chanx_left_in[12] sb_3__4_/chanx_left_in[13]
+ sb_3__4_/chanx_left_in[14] sb_3__4_/chanx_left_in[15] sb_3__4_/chanx_left_in[16]
+ sb_3__4_/chanx_left_in[17] sb_3__4_/chanx_left_in[18] sb_3__4_/chanx_left_in[19]
+ sb_3__4_/chanx_left_in[1] sb_3__4_/chanx_left_in[2] sb_3__4_/chanx_left_in[3] sb_3__4_/chanx_left_in[4]
+ sb_3__4_/chanx_left_in[5] sb_3__4_/chanx_left_in[6] sb_3__4_/chanx_left_in[7] sb_3__4_/chanx_left_in[8]
+ sb_3__4_/chanx_left_in[9] cbx_3__4_/clk_1_N_out cbx_3__4_/clk_1_S_out cbx_3__4_/clk_1_W_in
+ cbx_3__4_/clk_2_E_out cbx_3__4_/clk_2_W_in cbx_3__4_/clk_2_W_out cbx_3__4_/clk_3_E_out
+ sb_3__4_/clk_3_W_out sb_2__4_/clk_3_N_in cbx_3__4_/prog_clk_0_N_in cbx_3__4_/prog_clk_0_W_out
+ cbx_3__4_/prog_clk_1_N_out cbx_3__4_/prog_clk_1_S_out cbx_3__4_/prog_clk_1_W_in
+ cbx_3__4_/prog_clk_2_E_out cbx_3__4_/prog_clk_2_W_in cbx_3__4_/prog_clk_2_W_out
+ cbx_3__4_/prog_clk_3_E_out sb_3__4_/prog_clk_3_W_out sb_2__4_/prog_clk_3_N_in cbx_1__1_
Xgrid_clb_2__4_ cbx_2__3_/SC_OUT_TOP grid_clb_2__4_/SC_OUT_BOT cbx_2__4_/SC_IN_BOT
+ cby_2__4_/Test_en_W_out grid_clb_2__4_/Test_en_E_out cby_2__4_/Test_en_W_out cby_1__4_/Test_en_W_in
+ VGND VPWR cbx_2__3_/REGIN_FEEDTHROUGH grid_clb_2__4_/bottom_width_0_height_0__pin_51_
+ cby_1__4_/ccff_tail cby_2__4_/ccff_head cbx_2__3_/clk_1_N_out cbx_2__3_/clk_1_N_out
+ cby_2__4_/prog_clk_0_W_in cbx_2__3_/prog_clk_1_N_out grid_clb_2__4_/prog_clk_0_N_out
+ cbx_2__3_/prog_clk_1_N_out cbx_2__3_/prog_clk_0_N_in grid_clb_2__4_/prog_clk_0_W_out
+ cby_2__4_/left_grid_pin_16_ cby_2__4_/left_grid_pin_17_ cby_2__4_/left_grid_pin_18_
+ cby_2__4_/left_grid_pin_19_ cby_2__4_/left_grid_pin_20_ cby_2__4_/left_grid_pin_21_
+ cby_2__4_/left_grid_pin_22_ cby_2__4_/left_grid_pin_23_ cby_2__4_/left_grid_pin_24_
+ cby_2__4_/left_grid_pin_25_ cby_2__4_/left_grid_pin_26_ cby_2__4_/left_grid_pin_27_
+ cby_2__4_/left_grid_pin_28_ cby_2__4_/left_grid_pin_29_ cby_2__4_/left_grid_pin_30_
+ cby_2__4_/left_grid_pin_31_ sb_2__3_/top_left_grid_pin_42_ sb_2__4_/bottom_left_grid_pin_42_
+ sb_2__3_/top_left_grid_pin_43_ sb_2__4_/bottom_left_grid_pin_43_ sb_2__3_/top_left_grid_pin_44_
+ sb_2__4_/bottom_left_grid_pin_44_ sb_2__3_/top_left_grid_pin_45_ sb_2__4_/bottom_left_grid_pin_45_
+ sb_2__3_/top_left_grid_pin_46_ sb_2__4_/bottom_left_grid_pin_46_ sb_2__3_/top_left_grid_pin_47_
+ sb_2__4_/bottom_left_grid_pin_47_ sb_2__3_/top_left_grid_pin_48_ sb_2__4_/bottom_left_grid_pin_48_
+ sb_2__3_/top_left_grid_pin_49_ sb_2__4_/bottom_left_grid_pin_49_ cbx_2__4_/bottom_grid_pin_0_
+ cbx_2__4_/bottom_grid_pin_10_ cbx_2__4_/bottom_grid_pin_11_ cbx_2__4_/bottom_grid_pin_12_
+ cbx_2__4_/bottom_grid_pin_13_ cbx_2__4_/bottom_grid_pin_14_ cbx_2__4_/bottom_grid_pin_15_
+ cbx_2__4_/bottom_grid_pin_1_ cbx_2__4_/bottom_grid_pin_2_ cbx_2__4_/REGOUT_FEEDTHROUGH
+ grid_clb_2__4_/top_width_0_height_0__pin_33_ sb_2__4_/left_bottom_grid_pin_34_ sb_1__4_/right_bottom_grid_pin_34_
+ sb_2__4_/left_bottom_grid_pin_35_ sb_1__4_/right_bottom_grid_pin_35_ sb_2__4_/left_bottom_grid_pin_36_
+ sb_1__4_/right_bottom_grid_pin_36_ sb_2__4_/left_bottom_grid_pin_37_ sb_1__4_/right_bottom_grid_pin_37_
+ sb_2__4_/left_bottom_grid_pin_38_ sb_1__4_/right_bottom_grid_pin_38_ sb_2__4_/left_bottom_grid_pin_39_
+ sb_1__4_/right_bottom_grid_pin_39_ cbx_2__4_/bottom_grid_pin_3_ sb_2__4_/left_bottom_grid_pin_40_
+ sb_1__4_/right_bottom_grid_pin_40_ sb_2__4_/left_bottom_grid_pin_41_ sb_1__4_/right_bottom_grid_pin_41_
+ cbx_2__4_/bottom_grid_pin_4_ cbx_2__4_/bottom_grid_pin_5_ cbx_2__4_/bottom_grid_pin_6_
+ cbx_2__4_/bottom_grid_pin_7_ cbx_2__4_/bottom_grid_pin_8_ cbx_2__4_/bottom_grid_pin_9_
+ grid_clb
Xsb_7__1_ sb_7__1_/Test_en_N_out sb_7__1_/Test_en_S_in VGND VPWR sb_7__1_/bottom_left_grid_pin_42_
+ sb_7__1_/bottom_left_grid_pin_43_ sb_7__1_/bottom_left_grid_pin_44_ sb_7__1_/bottom_left_grid_pin_45_
+ sb_7__1_/bottom_left_grid_pin_46_ sb_7__1_/bottom_left_grid_pin_47_ sb_7__1_/bottom_left_grid_pin_48_
+ sb_7__1_/bottom_left_grid_pin_49_ sb_7__1_/ccff_head sb_7__1_/ccff_tail sb_7__1_/chanx_left_in[0]
+ sb_7__1_/chanx_left_in[10] sb_7__1_/chanx_left_in[11] sb_7__1_/chanx_left_in[12]
+ sb_7__1_/chanx_left_in[13] sb_7__1_/chanx_left_in[14] sb_7__1_/chanx_left_in[15]
+ sb_7__1_/chanx_left_in[16] sb_7__1_/chanx_left_in[17] sb_7__1_/chanx_left_in[18]
+ sb_7__1_/chanx_left_in[19] sb_7__1_/chanx_left_in[1] sb_7__1_/chanx_left_in[2] sb_7__1_/chanx_left_in[3]
+ sb_7__1_/chanx_left_in[4] sb_7__1_/chanx_left_in[5] sb_7__1_/chanx_left_in[6] sb_7__1_/chanx_left_in[7]
+ sb_7__1_/chanx_left_in[8] sb_7__1_/chanx_left_in[9] sb_7__1_/chanx_left_out[0] sb_7__1_/chanx_left_out[10]
+ sb_7__1_/chanx_left_out[11] sb_7__1_/chanx_left_out[12] sb_7__1_/chanx_left_out[13]
+ sb_7__1_/chanx_left_out[14] sb_7__1_/chanx_left_out[15] sb_7__1_/chanx_left_out[16]
+ sb_7__1_/chanx_left_out[17] sb_7__1_/chanx_left_out[18] sb_7__1_/chanx_left_out[19]
+ sb_7__1_/chanx_left_out[1] sb_7__1_/chanx_left_out[2] sb_7__1_/chanx_left_out[3]
+ sb_7__1_/chanx_left_out[4] sb_7__1_/chanx_left_out[5] sb_7__1_/chanx_left_out[6]
+ sb_7__1_/chanx_left_out[7] sb_7__1_/chanx_left_out[8] sb_7__1_/chanx_left_out[9]
+ sb_7__1_/chanx_right_in[0] sb_7__1_/chanx_right_in[10] sb_7__1_/chanx_right_in[11]
+ sb_7__1_/chanx_right_in[12] sb_7__1_/chanx_right_in[13] sb_7__1_/chanx_right_in[14]
+ sb_7__1_/chanx_right_in[15] sb_7__1_/chanx_right_in[16] sb_7__1_/chanx_right_in[17]
+ sb_7__1_/chanx_right_in[18] sb_7__1_/chanx_right_in[19] sb_7__1_/chanx_right_in[1]
+ sb_7__1_/chanx_right_in[2] sb_7__1_/chanx_right_in[3] sb_7__1_/chanx_right_in[4]
+ sb_7__1_/chanx_right_in[5] sb_7__1_/chanx_right_in[6] sb_7__1_/chanx_right_in[7]
+ sb_7__1_/chanx_right_in[8] sb_7__1_/chanx_right_in[9] cbx_8__1_/chanx_left_in[0]
+ cbx_8__1_/chanx_left_in[10] cbx_8__1_/chanx_left_in[11] cbx_8__1_/chanx_left_in[12]
+ cbx_8__1_/chanx_left_in[13] cbx_8__1_/chanx_left_in[14] cbx_8__1_/chanx_left_in[15]
+ cbx_8__1_/chanx_left_in[16] cbx_8__1_/chanx_left_in[17] cbx_8__1_/chanx_left_in[18]
+ cbx_8__1_/chanx_left_in[19] cbx_8__1_/chanx_left_in[1] cbx_8__1_/chanx_left_in[2]
+ cbx_8__1_/chanx_left_in[3] cbx_8__1_/chanx_left_in[4] cbx_8__1_/chanx_left_in[5]
+ cbx_8__1_/chanx_left_in[6] cbx_8__1_/chanx_left_in[7] cbx_8__1_/chanx_left_in[8]
+ cbx_8__1_/chanx_left_in[9] cby_7__1_/chany_top_out[0] cby_7__1_/chany_top_out[10]
+ cby_7__1_/chany_top_out[11] cby_7__1_/chany_top_out[12] cby_7__1_/chany_top_out[13]
+ cby_7__1_/chany_top_out[14] cby_7__1_/chany_top_out[15] cby_7__1_/chany_top_out[16]
+ cby_7__1_/chany_top_out[17] cby_7__1_/chany_top_out[18] cby_7__1_/chany_top_out[19]
+ cby_7__1_/chany_top_out[1] cby_7__1_/chany_top_out[2] cby_7__1_/chany_top_out[3]
+ cby_7__1_/chany_top_out[4] cby_7__1_/chany_top_out[5] cby_7__1_/chany_top_out[6]
+ cby_7__1_/chany_top_out[7] cby_7__1_/chany_top_out[8] cby_7__1_/chany_top_out[9]
+ cby_7__1_/chany_top_in[0] cby_7__1_/chany_top_in[10] cby_7__1_/chany_top_in[11]
+ cby_7__1_/chany_top_in[12] cby_7__1_/chany_top_in[13] cby_7__1_/chany_top_in[14]
+ cby_7__1_/chany_top_in[15] cby_7__1_/chany_top_in[16] cby_7__1_/chany_top_in[17]
+ cby_7__1_/chany_top_in[18] cby_7__1_/chany_top_in[19] cby_7__1_/chany_top_in[1]
+ cby_7__1_/chany_top_in[2] cby_7__1_/chany_top_in[3] cby_7__1_/chany_top_in[4] cby_7__1_/chany_top_in[5]
+ cby_7__1_/chany_top_in[6] cby_7__1_/chany_top_in[7] cby_7__1_/chany_top_in[8] cby_7__1_/chany_top_in[9]
+ sb_7__1_/chany_top_in[0] sb_7__1_/chany_top_in[10] sb_7__1_/chany_top_in[11] sb_7__1_/chany_top_in[12]
+ sb_7__1_/chany_top_in[13] sb_7__1_/chany_top_in[14] sb_7__1_/chany_top_in[15] sb_7__1_/chany_top_in[16]
+ sb_7__1_/chany_top_in[17] sb_7__1_/chany_top_in[18] sb_7__1_/chany_top_in[19] sb_7__1_/chany_top_in[1]
+ sb_7__1_/chany_top_in[2] sb_7__1_/chany_top_in[3] sb_7__1_/chany_top_in[4] sb_7__1_/chany_top_in[5]
+ sb_7__1_/chany_top_in[6] sb_7__1_/chany_top_in[7] sb_7__1_/chany_top_in[8] sb_7__1_/chany_top_in[9]
+ sb_7__1_/chany_top_out[0] sb_7__1_/chany_top_out[10] sb_7__1_/chany_top_out[11]
+ sb_7__1_/chany_top_out[12] sb_7__1_/chany_top_out[13] sb_7__1_/chany_top_out[14]
+ sb_7__1_/chany_top_out[15] sb_7__1_/chany_top_out[16] sb_7__1_/chany_top_out[17]
+ sb_7__1_/chany_top_out[18] sb_7__1_/chany_top_out[19] sb_7__1_/chany_top_out[1]
+ sb_7__1_/chany_top_out[2] sb_7__1_/chany_top_out[3] sb_7__1_/chany_top_out[4] sb_7__1_/chany_top_out[5]
+ sb_7__1_/chany_top_out[6] sb_7__1_/chany_top_out[7] sb_7__1_/chany_top_out[8] sb_7__1_/chany_top_out[9]
+ sb_7__1_/clk_1_E_out sb_7__1_/clk_1_N_in sb_7__1_/clk_1_W_out sb_7__1_/clk_2_E_out
+ sb_7__1_/clk_2_N_in sb_7__1_/clk_2_N_out sb_7__1_/clk_2_S_out sb_7__1_/clk_2_W_out
+ sb_7__1_/clk_3_E_out sb_7__1_/clk_3_N_in sb_7__1_/clk_3_N_out sb_7__1_/clk_3_S_out
+ sb_7__1_/clk_3_W_out sb_7__1_/left_bottom_grid_pin_34_ sb_7__1_/left_bottom_grid_pin_35_
+ sb_7__1_/left_bottom_grid_pin_36_ sb_7__1_/left_bottom_grid_pin_37_ sb_7__1_/left_bottom_grid_pin_38_
+ sb_7__1_/left_bottom_grid_pin_39_ sb_7__1_/left_bottom_grid_pin_40_ sb_7__1_/left_bottom_grid_pin_41_
+ sb_7__1_/prog_clk_0_N_in sb_7__1_/prog_clk_1_E_out sb_7__1_/prog_clk_1_N_in sb_7__1_/prog_clk_1_W_out
+ sb_7__1_/prog_clk_2_E_out sb_7__1_/prog_clk_2_N_in sb_7__1_/prog_clk_2_N_out sb_7__1_/prog_clk_2_S_out
+ sb_7__1_/prog_clk_2_W_out sb_7__1_/prog_clk_3_E_out sb_7__1_/prog_clk_3_N_in sb_7__1_/prog_clk_3_N_out
+ sb_7__1_/prog_clk_3_S_out sb_7__1_/prog_clk_3_W_out sb_7__1_/right_bottom_grid_pin_34_
+ sb_7__1_/right_bottom_grid_pin_35_ sb_7__1_/right_bottom_grid_pin_36_ sb_7__1_/right_bottom_grid_pin_37_
+ sb_7__1_/right_bottom_grid_pin_38_ sb_7__1_/right_bottom_grid_pin_39_ sb_7__1_/right_bottom_grid_pin_40_
+ sb_7__1_/right_bottom_grid_pin_41_ sb_7__1_/top_left_grid_pin_42_ sb_7__1_/top_left_grid_pin_43_
+ sb_7__1_/top_left_grid_pin_44_ sb_7__1_/top_left_grid_pin_45_ sb_7__1_/top_left_grid_pin_46_
+ sb_7__1_/top_left_grid_pin_47_ sb_7__1_/top_left_grid_pin_48_ sb_7__1_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_0__6_ VGND VPWR sb_0__6_/bottom_left_grid_pin_1_ sb_0__6_/ccff_head sb_0__6_/ccff_tail
+ sb_0__6_/chanx_right_in[0] sb_0__6_/chanx_right_in[10] sb_0__6_/chanx_right_in[11]
+ sb_0__6_/chanx_right_in[12] sb_0__6_/chanx_right_in[13] sb_0__6_/chanx_right_in[14]
+ sb_0__6_/chanx_right_in[15] sb_0__6_/chanx_right_in[16] sb_0__6_/chanx_right_in[17]
+ sb_0__6_/chanx_right_in[18] sb_0__6_/chanx_right_in[19] sb_0__6_/chanx_right_in[1]
+ sb_0__6_/chanx_right_in[2] sb_0__6_/chanx_right_in[3] sb_0__6_/chanx_right_in[4]
+ sb_0__6_/chanx_right_in[5] sb_0__6_/chanx_right_in[6] sb_0__6_/chanx_right_in[7]
+ sb_0__6_/chanx_right_in[8] sb_0__6_/chanx_right_in[9] cbx_1__6_/chanx_left_in[0]
+ cbx_1__6_/chanx_left_in[10] cbx_1__6_/chanx_left_in[11] cbx_1__6_/chanx_left_in[12]
+ cbx_1__6_/chanx_left_in[13] cbx_1__6_/chanx_left_in[14] cbx_1__6_/chanx_left_in[15]
+ cbx_1__6_/chanx_left_in[16] cbx_1__6_/chanx_left_in[17] cbx_1__6_/chanx_left_in[18]
+ cbx_1__6_/chanx_left_in[19] cbx_1__6_/chanx_left_in[1] cbx_1__6_/chanx_left_in[2]
+ cbx_1__6_/chanx_left_in[3] cbx_1__6_/chanx_left_in[4] cbx_1__6_/chanx_left_in[5]
+ cbx_1__6_/chanx_left_in[6] cbx_1__6_/chanx_left_in[7] cbx_1__6_/chanx_left_in[8]
+ cbx_1__6_/chanx_left_in[9] cby_0__6_/chany_top_out[0] cby_0__6_/chany_top_out[10]
+ cby_0__6_/chany_top_out[11] cby_0__6_/chany_top_out[12] cby_0__6_/chany_top_out[13]
+ cby_0__6_/chany_top_out[14] cby_0__6_/chany_top_out[15] cby_0__6_/chany_top_out[16]
+ cby_0__6_/chany_top_out[17] cby_0__6_/chany_top_out[18] cby_0__6_/chany_top_out[19]
+ cby_0__6_/chany_top_out[1] cby_0__6_/chany_top_out[2] cby_0__6_/chany_top_out[3]
+ cby_0__6_/chany_top_out[4] cby_0__6_/chany_top_out[5] cby_0__6_/chany_top_out[6]
+ cby_0__6_/chany_top_out[7] cby_0__6_/chany_top_out[8] cby_0__6_/chany_top_out[9]
+ cby_0__6_/chany_top_in[0] cby_0__6_/chany_top_in[10] cby_0__6_/chany_top_in[11]
+ cby_0__6_/chany_top_in[12] cby_0__6_/chany_top_in[13] cby_0__6_/chany_top_in[14]
+ cby_0__6_/chany_top_in[15] cby_0__6_/chany_top_in[16] cby_0__6_/chany_top_in[17]
+ cby_0__6_/chany_top_in[18] cby_0__6_/chany_top_in[19] cby_0__6_/chany_top_in[1]
+ cby_0__6_/chany_top_in[2] cby_0__6_/chany_top_in[3] cby_0__6_/chany_top_in[4] cby_0__6_/chany_top_in[5]
+ cby_0__6_/chany_top_in[6] cby_0__6_/chany_top_in[7] cby_0__6_/chany_top_in[8] cby_0__6_/chany_top_in[9]
+ sb_0__6_/chany_top_in[0] sb_0__6_/chany_top_in[10] sb_0__6_/chany_top_in[11] sb_0__6_/chany_top_in[12]
+ sb_0__6_/chany_top_in[13] sb_0__6_/chany_top_in[14] sb_0__6_/chany_top_in[15] sb_0__6_/chany_top_in[16]
+ sb_0__6_/chany_top_in[17] sb_0__6_/chany_top_in[18] sb_0__6_/chany_top_in[19] sb_0__6_/chany_top_in[1]
+ sb_0__6_/chany_top_in[2] sb_0__6_/chany_top_in[3] sb_0__6_/chany_top_in[4] sb_0__6_/chany_top_in[5]
+ sb_0__6_/chany_top_in[6] sb_0__6_/chany_top_in[7] sb_0__6_/chany_top_in[8] sb_0__6_/chany_top_in[9]
+ sb_0__6_/chany_top_out[0] sb_0__6_/chany_top_out[10] sb_0__6_/chany_top_out[11]
+ sb_0__6_/chany_top_out[12] sb_0__6_/chany_top_out[13] sb_0__6_/chany_top_out[14]
+ sb_0__6_/chany_top_out[15] sb_0__6_/chany_top_out[16] sb_0__6_/chany_top_out[17]
+ sb_0__6_/chany_top_out[18] sb_0__6_/chany_top_out[19] sb_0__6_/chany_top_out[1]
+ sb_0__6_/chany_top_out[2] sb_0__6_/chany_top_out[3] sb_0__6_/chany_top_out[4] sb_0__6_/chany_top_out[5]
+ sb_0__6_/chany_top_out[6] sb_0__6_/chany_top_out[7] sb_0__6_/chany_top_out[8] sb_0__6_/chany_top_out[9]
+ sb_0__6_/prog_clk_0_E_in sb_0__6_/right_bottom_grid_pin_34_ sb_0__6_/right_bottom_grid_pin_35_
+ sb_0__6_/right_bottom_grid_pin_36_ sb_0__6_/right_bottom_grid_pin_37_ sb_0__6_/right_bottom_grid_pin_38_
+ sb_0__6_/right_bottom_grid_pin_39_ sb_0__6_/right_bottom_grid_pin_40_ sb_0__6_/right_bottom_grid_pin_41_
+ sb_0__6_/top_left_grid_pin_1_ sb_0__1_
Xcby_6__5_ cby_6__5_/Test_en_W_in cby_6__5_/Test_en_E_out cby_6__5_/Test_en_N_out
+ cby_6__5_/Test_en_W_in cby_6__5_/Test_en_W_in cby_6__5_/Test_en_W_out VGND VPWR
+ cby_6__5_/ccff_head cby_6__5_/ccff_tail sb_6__4_/chany_top_out[0] sb_6__4_/chany_top_out[10]
+ sb_6__4_/chany_top_out[11] sb_6__4_/chany_top_out[12] sb_6__4_/chany_top_out[13]
+ sb_6__4_/chany_top_out[14] sb_6__4_/chany_top_out[15] sb_6__4_/chany_top_out[16]
+ sb_6__4_/chany_top_out[17] sb_6__4_/chany_top_out[18] sb_6__4_/chany_top_out[19]
+ sb_6__4_/chany_top_out[1] sb_6__4_/chany_top_out[2] sb_6__4_/chany_top_out[3] sb_6__4_/chany_top_out[4]
+ sb_6__4_/chany_top_out[5] sb_6__4_/chany_top_out[6] sb_6__4_/chany_top_out[7] sb_6__4_/chany_top_out[8]
+ sb_6__4_/chany_top_out[9] sb_6__4_/chany_top_in[0] sb_6__4_/chany_top_in[10] sb_6__4_/chany_top_in[11]
+ sb_6__4_/chany_top_in[12] sb_6__4_/chany_top_in[13] sb_6__4_/chany_top_in[14] sb_6__4_/chany_top_in[15]
+ sb_6__4_/chany_top_in[16] sb_6__4_/chany_top_in[17] sb_6__4_/chany_top_in[18] sb_6__4_/chany_top_in[19]
+ sb_6__4_/chany_top_in[1] sb_6__4_/chany_top_in[2] sb_6__4_/chany_top_in[3] sb_6__4_/chany_top_in[4]
+ sb_6__4_/chany_top_in[5] sb_6__4_/chany_top_in[6] sb_6__4_/chany_top_in[7] sb_6__4_/chany_top_in[8]
+ sb_6__4_/chany_top_in[9] cby_6__5_/chany_top_in[0] cby_6__5_/chany_top_in[10] cby_6__5_/chany_top_in[11]
+ cby_6__5_/chany_top_in[12] cby_6__5_/chany_top_in[13] cby_6__5_/chany_top_in[14]
+ cby_6__5_/chany_top_in[15] cby_6__5_/chany_top_in[16] cby_6__5_/chany_top_in[17]
+ cby_6__5_/chany_top_in[18] cby_6__5_/chany_top_in[19] cby_6__5_/chany_top_in[1]
+ cby_6__5_/chany_top_in[2] cby_6__5_/chany_top_in[3] cby_6__5_/chany_top_in[4] cby_6__5_/chany_top_in[5]
+ cby_6__5_/chany_top_in[6] cby_6__5_/chany_top_in[7] cby_6__5_/chany_top_in[8] cby_6__5_/chany_top_in[9]
+ cby_6__5_/chany_top_out[0] cby_6__5_/chany_top_out[10] cby_6__5_/chany_top_out[11]
+ cby_6__5_/chany_top_out[12] cby_6__5_/chany_top_out[13] cby_6__5_/chany_top_out[14]
+ cby_6__5_/chany_top_out[15] cby_6__5_/chany_top_out[16] cby_6__5_/chany_top_out[17]
+ cby_6__5_/chany_top_out[18] cby_6__5_/chany_top_out[19] cby_6__5_/chany_top_out[1]
+ cby_6__5_/chany_top_out[2] cby_6__5_/chany_top_out[3] cby_6__5_/chany_top_out[4]
+ cby_6__5_/chany_top_out[5] cby_6__5_/chany_top_out[6] cby_6__5_/chany_top_out[7]
+ cby_6__5_/chany_top_out[8] cby_6__5_/chany_top_out[9] cby_6__5_/clk_2_N_out cby_6__5_/clk_2_S_in
+ cby_6__5_/clk_2_S_out sb_6__5_/clk_3_N_in sb_6__4_/clk_3_N_out cby_6__5_/clk_3_S_out
+ cby_6__5_/left_grid_pin_16_ cby_6__5_/left_grid_pin_17_ cby_6__5_/left_grid_pin_18_
+ cby_6__5_/left_grid_pin_19_ cby_6__5_/left_grid_pin_20_ cby_6__5_/left_grid_pin_21_
+ cby_6__5_/left_grid_pin_22_ cby_6__5_/left_grid_pin_23_ cby_6__5_/left_grid_pin_24_
+ cby_6__5_/left_grid_pin_25_ cby_6__5_/left_grid_pin_26_ cby_6__5_/left_grid_pin_27_
+ cby_6__5_/left_grid_pin_28_ cby_6__5_/left_grid_pin_29_ cby_6__5_/left_grid_pin_30_
+ cby_6__5_/left_grid_pin_31_ cby_6__5_/prog_clk_0_N_out sb_6__4_/prog_clk_0_N_in
+ cby_6__5_/prog_clk_0_W_in cby_6__5_/prog_clk_2_N_out cby_6__5_/prog_clk_2_S_in cby_6__5_/prog_clk_2_S_out
+ sb_6__5_/prog_clk_3_N_in sb_6__4_/prog_clk_3_N_out cby_6__5_/prog_clk_3_S_out cby_1__1_
Xcby_3__2_ cby_3__2_/Test_en_W_in cby_3__2_/Test_en_E_out cby_3__2_/Test_en_N_out
+ cby_3__2_/Test_en_W_in cby_3__2_/Test_en_W_in cby_3__2_/Test_en_W_out VGND VPWR
+ cby_3__2_/ccff_head cby_3__2_/ccff_tail sb_3__1_/chany_top_out[0] sb_3__1_/chany_top_out[10]
+ sb_3__1_/chany_top_out[11] sb_3__1_/chany_top_out[12] sb_3__1_/chany_top_out[13]
+ sb_3__1_/chany_top_out[14] sb_3__1_/chany_top_out[15] sb_3__1_/chany_top_out[16]
+ sb_3__1_/chany_top_out[17] sb_3__1_/chany_top_out[18] sb_3__1_/chany_top_out[19]
+ sb_3__1_/chany_top_out[1] sb_3__1_/chany_top_out[2] sb_3__1_/chany_top_out[3] sb_3__1_/chany_top_out[4]
+ sb_3__1_/chany_top_out[5] sb_3__1_/chany_top_out[6] sb_3__1_/chany_top_out[7] sb_3__1_/chany_top_out[8]
+ sb_3__1_/chany_top_out[9] sb_3__1_/chany_top_in[0] sb_3__1_/chany_top_in[10] sb_3__1_/chany_top_in[11]
+ sb_3__1_/chany_top_in[12] sb_3__1_/chany_top_in[13] sb_3__1_/chany_top_in[14] sb_3__1_/chany_top_in[15]
+ sb_3__1_/chany_top_in[16] sb_3__1_/chany_top_in[17] sb_3__1_/chany_top_in[18] sb_3__1_/chany_top_in[19]
+ sb_3__1_/chany_top_in[1] sb_3__1_/chany_top_in[2] sb_3__1_/chany_top_in[3] sb_3__1_/chany_top_in[4]
+ sb_3__1_/chany_top_in[5] sb_3__1_/chany_top_in[6] sb_3__1_/chany_top_in[7] sb_3__1_/chany_top_in[8]
+ sb_3__1_/chany_top_in[9] cby_3__2_/chany_top_in[0] cby_3__2_/chany_top_in[10] cby_3__2_/chany_top_in[11]
+ cby_3__2_/chany_top_in[12] cby_3__2_/chany_top_in[13] cby_3__2_/chany_top_in[14]
+ cby_3__2_/chany_top_in[15] cby_3__2_/chany_top_in[16] cby_3__2_/chany_top_in[17]
+ cby_3__2_/chany_top_in[18] cby_3__2_/chany_top_in[19] cby_3__2_/chany_top_in[1]
+ cby_3__2_/chany_top_in[2] cby_3__2_/chany_top_in[3] cby_3__2_/chany_top_in[4] cby_3__2_/chany_top_in[5]
+ cby_3__2_/chany_top_in[6] cby_3__2_/chany_top_in[7] cby_3__2_/chany_top_in[8] cby_3__2_/chany_top_in[9]
+ cby_3__2_/chany_top_out[0] cby_3__2_/chany_top_out[10] cby_3__2_/chany_top_out[11]
+ cby_3__2_/chany_top_out[12] cby_3__2_/chany_top_out[13] cby_3__2_/chany_top_out[14]
+ cby_3__2_/chany_top_out[15] cby_3__2_/chany_top_out[16] cby_3__2_/chany_top_out[17]
+ cby_3__2_/chany_top_out[18] cby_3__2_/chany_top_out[19] cby_3__2_/chany_top_out[1]
+ cby_3__2_/chany_top_out[2] cby_3__2_/chany_top_out[3] cby_3__2_/chany_top_out[4]
+ cby_3__2_/chany_top_out[5] cby_3__2_/chany_top_out[6] cby_3__2_/chany_top_out[7]
+ cby_3__2_/chany_top_out[8] cby_3__2_/chany_top_out[9] cby_3__2_/clk_2_N_out sb_3__2_/clk_2_S_out
+ sb_3__1_/clk_1_N_in cby_3__2_/clk_3_N_out cby_3__2_/clk_3_S_in cby_3__2_/clk_3_S_out
+ cby_3__2_/left_grid_pin_16_ cby_3__2_/left_grid_pin_17_ cby_3__2_/left_grid_pin_18_
+ cby_3__2_/left_grid_pin_19_ cby_3__2_/left_grid_pin_20_ cby_3__2_/left_grid_pin_21_
+ cby_3__2_/left_grid_pin_22_ cby_3__2_/left_grid_pin_23_ cby_3__2_/left_grid_pin_24_
+ cby_3__2_/left_grid_pin_25_ cby_3__2_/left_grid_pin_26_ cby_3__2_/left_grid_pin_27_
+ cby_3__2_/left_grid_pin_28_ cby_3__2_/left_grid_pin_29_ cby_3__2_/left_grid_pin_30_
+ cby_3__2_/left_grid_pin_31_ cby_3__2_/prog_clk_0_N_out sb_3__1_/prog_clk_0_N_in
+ cby_3__2_/prog_clk_0_W_in cby_3__2_/prog_clk_2_N_out sb_3__2_/prog_clk_2_S_out sb_3__1_/prog_clk_1_N_in
+ cby_3__2_/prog_clk_3_N_out cby_3__2_/prog_clk_3_S_in cby_3__2_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_6__6_ cbx_6__6_/REGIN_FEEDTHROUGH cbx_6__6_/REGOUT_FEEDTHROUGH cbx_6__6_/SC_IN_BOT
+ cbx_6__6_/SC_IN_TOP cbx_6__6_/SC_OUT_BOT cbx_6__6_/SC_OUT_TOP VGND VPWR cbx_6__6_/bottom_grid_pin_0_
+ cbx_6__6_/bottom_grid_pin_10_ cbx_6__6_/bottom_grid_pin_11_ cbx_6__6_/bottom_grid_pin_12_
+ cbx_6__6_/bottom_grid_pin_13_ cbx_6__6_/bottom_grid_pin_14_ cbx_6__6_/bottom_grid_pin_15_
+ cbx_6__6_/bottom_grid_pin_1_ cbx_6__6_/bottom_grid_pin_2_ cbx_6__6_/bottom_grid_pin_3_
+ cbx_6__6_/bottom_grid_pin_4_ cbx_6__6_/bottom_grid_pin_5_ cbx_6__6_/bottom_grid_pin_6_
+ cbx_6__6_/bottom_grid_pin_7_ cbx_6__6_/bottom_grid_pin_8_ cbx_6__6_/bottom_grid_pin_9_
+ sb_6__6_/ccff_tail sb_5__6_/ccff_head cbx_6__6_/chanx_left_in[0] cbx_6__6_/chanx_left_in[10]
+ cbx_6__6_/chanx_left_in[11] cbx_6__6_/chanx_left_in[12] cbx_6__6_/chanx_left_in[13]
+ cbx_6__6_/chanx_left_in[14] cbx_6__6_/chanx_left_in[15] cbx_6__6_/chanx_left_in[16]
+ cbx_6__6_/chanx_left_in[17] cbx_6__6_/chanx_left_in[18] cbx_6__6_/chanx_left_in[19]
+ cbx_6__6_/chanx_left_in[1] cbx_6__6_/chanx_left_in[2] cbx_6__6_/chanx_left_in[3]
+ cbx_6__6_/chanx_left_in[4] cbx_6__6_/chanx_left_in[5] cbx_6__6_/chanx_left_in[6]
+ cbx_6__6_/chanx_left_in[7] cbx_6__6_/chanx_left_in[8] cbx_6__6_/chanx_left_in[9]
+ sb_5__6_/chanx_right_in[0] sb_5__6_/chanx_right_in[10] sb_5__6_/chanx_right_in[11]
+ sb_5__6_/chanx_right_in[12] sb_5__6_/chanx_right_in[13] sb_5__6_/chanx_right_in[14]
+ sb_5__6_/chanx_right_in[15] sb_5__6_/chanx_right_in[16] sb_5__6_/chanx_right_in[17]
+ sb_5__6_/chanx_right_in[18] sb_5__6_/chanx_right_in[19] sb_5__6_/chanx_right_in[1]
+ sb_5__6_/chanx_right_in[2] sb_5__6_/chanx_right_in[3] sb_5__6_/chanx_right_in[4]
+ sb_5__6_/chanx_right_in[5] sb_5__6_/chanx_right_in[6] sb_5__6_/chanx_right_in[7]
+ sb_5__6_/chanx_right_in[8] sb_5__6_/chanx_right_in[9] sb_6__6_/chanx_left_out[0]
+ sb_6__6_/chanx_left_out[10] sb_6__6_/chanx_left_out[11] sb_6__6_/chanx_left_out[12]
+ sb_6__6_/chanx_left_out[13] sb_6__6_/chanx_left_out[14] sb_6__6_/chanx_left_out[15]
+ sb_6__6_/chanx_left_out[16] sb_6__6_/chanx_left_out[17] sb_6__6_/chanx_left_out[18]
+ sb_6__6_/chanx_left_out[19] sb_6__6_/chanx_left_out[1] sb_6__6_/chanx_left_out[2]
+ sb_6__6_/chanx_left_out[3] sb_6__6_/chanx_left_out[4] sb_6__6_/chanx_left_out[5]
+ sb_6__6_/chanx_left_out[6] sb_6__6_/chanx_left_out[7] sb_6__6_/chanx_left_out[8]
+ sb_6__6_/chanx_left_out[9] sb_6__6_/chanx_left_in[0] sb_6__6_/chanx_left_in[10]
+ sb_6__6_/chanx_left_in[11] sb_6__6_/chanx_left_in[12] sb_6__6_/chanx_left_in[13]
+ sb_6__6_/chanx_left_in[14] sb_6__6_/chanx_left_in[15] sb_6__6_/chanx_left_in[16]
+ sb_6__6_/chanx_left_in[17] sb_6__6_/chanx_left_in[18] sb_6__6_/chanx_left_in[19]
+ sb_6__6_/chanx_left_in[1] sb_6__6_/chanx_left_in[2] sb_6__6_/chanx_left_in[3] sb_6__6_/chanx_left_in[4]
+ sb_6__6_/chanx_left_in[5] sb_6__6_/chanx_left_in[6] sb_6__6_/chanx_left_in[7] sb_6__6_/chanx_left_in[8]
+ sb_6__6_/chanx_left_in[9] cbx_6__6_/clk_1_N_out cbx_6__6_/clk_1_S_out cbx_6__6_/clk_1_W_in
+ cbx_6__6_/clk_2_E_out sb_6__6_/clk_2_W_out sb_5__6_/clk_2_N_in cbx_6__6_/clk_3_E_out
+ cbx_6__6_/clk_3_W_in cbx_6__6_/clk_3_W_out cbx_6__6_/prog_clk_0_N_in cbx_6__6_/prog_clk_0_W_out
+ cbx_6__6_/prog_clk_1_N_out cbx_6__6_/prog_clk_1_S_out cbx_6__6_/prog_clk_1_W_in
+ cbx_6__6_/prog_clk_2_E_out sb_6__6_/prog_clk_2_W_out sb_5__6_/prog_clk_2_N_in cbx_6__6_/prog_clk_3_E_out
+ cbx_6__6_/prog_clk_3_W_in cbx_6__6_/prog_clk_3_W_out cbx_1__1_
Xgrid_clb_5__6_ cbx_5__6_/SC_OUT_BOT cbx_5__5_/SC_IN_TOP grid_clb_5__6_/SC_OUT_TOP
+ cby_4__6_/Test_en_E_out cby_5__6_/Test_en_W_in cby_4__6_/Test_en_E_out grid_clb_5__6_/Test_en_W_out
+ VGND VPWR cbx_5__5_/REGIN_FEEDTHROUGH grid_clb_5__6_/bottom_width_0_height_0__pin_51_
+ cby_4__6_/ccff_tail cby_5__6_/ccff_head cbx_5__5_/clk_1_N_out cbx_5__5_/clk_1_N_out
+ cby_5__6_/prog_clk_0_W_in cbx_5__5_/prog_clk_1_N_out grid_clb_5__6_/prog_clk_0_N_out
+ cbx_5__5_/prog_clk_1_N_out cbx_5__5_/prog_clk_0_N_in grid_clb_5__6_/prog_clk_0_W_out
+ cby_5__6_/left_grid_pin_16_ cby_5__6_/left_grid_pin_17_ cby_5__6_/left_grid_pin_18_
+ cby_5__6_/left_grid_pin_19_ cby_5__6_/left_grid_pin_20_ cby_5__6_/left_grid_pin_21_
+ cby_5__6_/left_grid_pin_22_ cby_5__6_/left_grid_pin_23_ cby_5__6_/left_grid_pin_24_
+ cby_5__6_/left_grid_pin_25_ cby_5__6_/left_grid_pin_26_ cby_5__6_/left_grid_pin_27_
+ cby_5__6_/left_grid_pin_28_ cby_5__6_/left_grid_pin_29_ cby_5__6_/left_grid_pin_30_
+ cby_5__6_/left_grid_pin_31_ sb_5__5_/top_left_grid_pin_42_ sb_5__6_/bottom_left_grid_pin_42_
+ sb_5__5_/top_left_grid_pin_43_ sb_5__6_/bottom_left_grid_pin_43_ sb_5__5_/top_left_grid_pin_44_
+ sb_5__6_/bottom_left_grid_pin_44_ sb_5__5_/top_left_grid_pin_45_ sb_5__6_/bottom_left_grid_pin_45_
+ sb_5__5_/top_left_grid_pin_46_ sb_5__6_/bottom_left_grid_pin_46_ sb_5__5_/top_left_grid_pin_47_
+ sb_5__6_/bottom_left_grid_pin_47_ sb_5__5_/top_left_grid_pin_48_ sb_5__6_/bottom_left_grid_pin_48_
+ sb_5__5_/top_left_grid_pin_49_ sb_5__6_/bottom_left_grid_pin_49_ cbx_5__6_/bottom_grid_pin_0_
+ cbx_5__6_/bottom_grid_pin_10_ cbx_5__6_/bottom_grid_pin_11_ cbx_5__6_/bottom_grid_pin_12_
+ cbx_5__6_/bottom_grid_pin_13_ cbx_5__6_/bottom_grid_pin_14_ cbx_5__6_/bottom_grid_pin_15_
+ cbx_5__6_/bottom_grid_pin_1_ cbx_5__6_/bottom_grid_pin_2_ cbx_5__6_/REGOUT_FEEDTHROUGH
+ grid_clb_5__6_/top_width_0_height_0__pin_33_ sb_5__6_/left_bottom_grid_pin_34_ sb_4__6_/right_bottom_grid_pin_34_
+ sb_5__6_/left_bottom_grid_pin_35_ sb_4__6_/right_bottom_grid_pin_35_ sb_5__6_/left_bottom_grid_pin_36_
+ sb_4__6_/right_bottom_grid_pin_36_ sb_5__6_/left_bottom_grid_pin_37_ sb_4__6_/right_bottom_grid_pin_37_
+ sb_5__6_/left_bottom_grid_pin_38_ sb_4__6_/right_bottom_grid_pin_38_ sb_5__6_/left_bottom_grid_pin_39_
+ sb_4__6_/right_bottom_grid_pin_39_ cbx_5__6_/bottom_grid_pin_3_ sb_5__6_/left_bottom_grid_pin_40_
+ sb_4__6_/right_bottom_grid_pin_40_ sb_5__6_/left_bottom_grid_pin_41_ sb_4__6_/right_bottom_grid_pin_41_
+ cbx_5__6_/bottom_grid_pin_4_ cbx_5__6_/bottom_grid_pin_5_ cbx_5__6_/bottom_grid_pin_6_
+ cbx_5__6_/bottom_grid_pin_7_ cbx_5__6_/bottom_grid_pin_8_ cbx_5__6_/bottom_grid_pin_9_
+ grid_clb
Xcbx_3__3_ cbx_3__3_/REGIN_FEEDTHROUGH cbx_3__3_/REGOUT_FEEDTHROUGH cbx_3__3_/SC_IN_BOT
+ cbx_3__3_/SC_IN_TOP cbx_3__3_/SC_OUT_BOT cbx_3__3_/SC_OUT_TOP VGND VPWR cbx_3__3_/bottom_grid_pin_0_
+ cbx_3__3_/bottom_grid_pin_10_ cbx_3__3_/bottom_grid_pin_11_ cbx_3__3_/bottom_grid_pin_12_
+ cbx_3__3_/bottom_grid_pin_13_ cbx_3__3_/bottom_grid_pin_14_ cbx_3__3_/bottom_grid_pin_15_
+ cbx_3__3_/bottom_grid_pin_1_ cbx_3__3_/bottom_grid_pin_2_ cbx_3__3_/bottom_grid_pin_3_
+ cbx_3__3_/bottom_grid_pin_4_ cbx_3__3_/bottom_grid_pin_5_ cbx_3__3_/bottom_grid_pin_6_
+ cbx_3__3_/bottom_grid_pin_7_ cbx_3__3_/bottom_grid_pin_8_ cbx_3__3_/bottom_grid_pin_9_
+ sb_3__3_/ccff_tail sb_2__3_/ccff_head cbx_3__3_/chanx_left_in[0] cbx_3__3_/chanx_left_in[10]
+ cbx_3__3_/chanx_left_in[11] cbx_3__3_/chanx_left_in[12] cbx_3__3_/chanx_left_in[13]
+ cbx_3__3_/chanx_left_in[14] cbx_3__3_/chanx_left_in[15] cbx_3__3_/chanx_left_in[16]
+ cbx_3__3_/chanx_left_in[17] cbx_3__3_/chanx_left_in[18] cbx_3__3_/chanx_left_in[19]
+ cbx_3__3_/chanx_left_in[1] cbx_3__3_/chanx_left_in[2] cbx_3__3_/chanx_left_in[3]
+ cbx_3__3_/chanx_left_in[4] cbx_3__3_/chanx_left_in[5] cbx_3__3_/chanx_left_in[6]
+ cbx_3__3_/chanx_left_in[7] cbx_3__3_/chanx_left_in[8] cbx_3__3_/chanx_left_in[9]
+ sb_2__3_/chanx_right_in[0] sb_2__3_/chanx_right_in[10] sb_2__3_/chanx_right_in[11]
+ sb_2__3_/chanx_right_in[12] sb_2__3_/chanx_right_in[13] sb_2__3_/chanx_right_in[14]
+ sb_2__3_/chanx_right_in[15] sb_2__3_/chanx_right_in[16] sb_2__3_/chanx_right_in[17]
+ sb_2__3_/chanx_right_in[18] sb_2__3_/chanx_right_in[19] sb_2__3_/chanx_right_in[1]
+ sb_2__3_/chanx_right_in[2] sb_2__3_/chanx_right_in[3] sb_2__3_/chanx_right_in[4]
+ sb_2__3_/chanx_right_in[5] sb_2__3_/chanx_right_in[6] sb_2__3_/chanx_right_in[7]
+ sb_2__3_/chanx_right_in[8] sb_2__3_/chanx_right_in[9] sb_3__3_/chanx_left_out[0]
+ sb_3__3_/chanx_left_out[10] sb_3__3_/chanx_left_out[11] sb_3__3_/chanx_left_out[12]
+ sb_3__3_/chanx_left_out[13] sb_3__3_/chanx_left_out[14] sb_3__3_/chanx_left_out[15]
+ sb_3__3_/chanx_left_out[16] sb_3__3_/chanx_left_out[17] sb_3__3_/chanx_left_out[18]
+ sb_3__3_/chanx_left_out[19] sb_3__3_/chanx_left_out[1] sb_3__3_/chanx_left_out[2]
+ sb_3__3_/chanx_left_out[3] sb_3__3_/chanx_left_out[4] sb_3__3_/chanx_left_out[5]
+ sb_3__3_/chanx_left_out[6] sb_3__3_/chanx_left_out[7] sb_3__3_/chanx_left_out[8]
+ sb_3__3_/chanx_left_out[9] sb_3__3_/chanx_left_in[0] sb_3__3_/chanx_left_in[10]
+ sb_3__3_/chanx_left_in[11] sb_3__3_/chanx_left_in[12] sb_3__3_/chanx_left_in[13]
+ sb_3__3_/chanx_left_in[14] sb_3__3_/chanx_left_in[15] sb_3__3_/chanx_left_in[16]
+ sb_3__3_/chanx_left_in[17] sb_3__3_/chanx_left_in[18] sb_3__3_/chanx_left_in[19]
+ sb_3__3_/chanx_left_in[1] sb_3__3_/chanx_left_in[2] sb_3__3_/chanx_left_in[3] sb_3__3_/chanx_left_in[4]
+ sb_3__3_/chanx_left_in[5] sb_3__3_/chanx_left_in[6] sb_3__3_/chanx_left_in[7] sb_3__3_/chanx_left_in[8]
+ sb_3__3_/chanx_left_in[9] cbx_3__3_/clk_1_N_out cbx_3__3_/clk_1_S_out sb_3__3_/clk_1_W_out
+ cbx_3__3_/clk_2_E_out cbx_3__3_/clk_2_W_in cbx_3__3_/clk_2_W_out cbx_3__3_/clk_3_E_out
+ cbx_3__3_/clk_3_W_in cbx_3__3_/clk_3_W_out cbx_3__3_/prog_clk_0_N_in cbx_3__3_/prog_clk_0_W_out
+ cbx_3__3_/prog_clk_1_N_out cbx_3__3_/prog_clk_1_S_out sb_3__3_/prog_clk_1_W_out
+ cbx_3__3_/prog_clk_2_E_out cbx_3__3_/prog_clk_2_W_in cbx_3__3_/prog_clk_2_W_out
+ cbx_3__3_/prog_clk_3_E_out cbx_3__3_/prog_clk_3_W_in cbx_3__3_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_7__0_ sb_7__0_/SC_IN_TOP sb_7__0_/SC_OUT_TOP sb_7__0_/Test_en_N_out sb_7__0_/Test_en_S_in
+ VGND VPWR sb_7__0_/ccff_head sb_7__0_/ccff_tail sb_7__0_/chanx_left_in[0] sb_7__0_/chanx_left_in[10]
+ sb_7__0_/chanx_left_in[11] sb_7__0_/chanx_left_in[12] sb_7__0_/chanx_left_in[13]
+ sb_7__0_/chanx_left_in[14] sb_7__0_/chanx_left_in[15] sb_7__0_/chanx_left_in[16]
+ sb_7__0_/chanx_left_in[17] sb_7__0_/chanx_left_in[18] sb_7__0_/chanx_left_in[19]
+ sb_7__0_/chanx_left_in[1] sb_7__0_/chanx_left_in[2] sb_7__0_/chanx_left_in[3] sb_7__0_/chanx_left_in[4]
+ sb_7__0_/chanx_left_in[5] sb_7__0_/chanx_left_in[6] sb_7__0_/chanx_left_in[7] sb_7__0_/chanx_left_in[8]
+ sb_7__0_/chanx_left_in[9] sb_7__0_/chanx_left_out[0] sb_7__0_/chanx_left_out[10]
+ sb_7__0_/chanx_left_out[11] sb_7__0_/chanx_left_out[12] sb_7__0_/chanx_left_out[13]
+ sb_7__0_/chanx_left_out[14] sb_7__0_/chanx_left_out[15] sb_7__0_/chanx_left_out[16]
+ sb_7__0_/chanx_left_out[17] sb_7__0_/chanx_left_out[18] sb_7__0_/chanx_left_out[19]
+ sb_7__0_/chanx_left_out[1] sb_7__0_/chanx_left_out[2] sb_7__0_/chanx_left_out[3]
+ sb_7__0_/chanx_left_out[4] sb_7__0_/chanx_left_out[5] sb_7__0_/chanx_left_out[6]
+ sb_7__0_/chanx_left_out[7] sb_7__0_/chanx_left_out[8] sb_7__0_/chanx_left_out[9]
+ sb_7__0_/chanx_right_in[0] sb_7__0_/chanx_right_in[10] sb_7__0_/chanx_right_in[11]
+ sb_7__0_/chanx_right_in[12] sb_7__0_/chanx_right_in[13] sb_7__0_/chanx_right_in[14]
+ sb_7__0_/chanx_right_in[15] sb_7__0_/chanx_right_in[16] sb_7__0_/chanx_right_in[17]
+ sb_7__0_/chanx_right_in[18] sb_7__0_/chanx_right_in[19] sb_7__0_/chanx_right_in[1]
+ sb_7__0_/chanx_right_in[2] sb_7__0_/chanx_right_in[3] sb_7__0_/chanx_right_in[4]
+ sb_7__0_/chanx_right_in[5] sb_7__0_/chanx_right_in[6] sb_7__0_/chanx_right_in[7]
+ sb_7__0_/chanx_right_in[8] sb_7__0_/chanx_right_in[9] cbx_8__0_/chanx_left_in[0]
+ cbx_8__0_/chanx_left_in[10] cbx_8__0_/chanx_left_in[11] cbx_8__0_/chanx_left_in[12]
+ cbx_8__0_/chanx_left_in[13] cbx_8__0_/chanx_left_in[14] cbx_8__0_/chanx_left_in[15]
+ cbx_8__0_/chanx_left_in[16] cbx_8__0_/chanx_left_in[17] cbx_8__0_/chanx_left_in[18]
+ cbx_8__0_/chanx_left_in[19] cbx_8__0_/chanx_left_in[1] cbx_8__0_/chanx_left_in[2]
+ cbx_8__0_/chanx_left_in[3] cbx_8__0_/chanx_left_in[4] cbx_8__0_/chanx_left_in[5]
+ cbx_8__0_/chanx_left_in[6] cbx_8__0_/chanx_left_in[7] cbx_8__0_/chanx_left_in[8]
+ cbx_8__0_/chanx_left_in[9] sb_7__0_/chany_top_in[0] sb_7__0_/chany_top_in[10] sb_7__0_/chany_top_in[11]
+ sb_7__0_/chany_top_in[12] sb_7__0_/chany_top_in[13] sb_7__0_/chany_top_in[14] sb_7__0_/chany_top_in[15]
+ sb_7__0_/chany_top_in[16] sb_7__0_/chany_top_in[17] sb_7__0_/chany_top_in[18] sb_7__0_/chany_top_in[19]
+ sb_7__0_/chany_top_in[1] sb_7__0_/chany_top_in[2] sb_7__0_/chany_top_in[3] sb_7__0_/chany_top_in[4]
+ sb_7__0_/chany_top_in[5] sb_7__0_/chany_top_in[6] sb_7__0_/chany_top_in[7] sb_7__0_/chany_top_in[8]
+ sb_7__0_/chany_top_in[9] sb_7__0_/chany_top_out[0] sb_7__0_/chany_top_out[10] sb_7__0_/chany_top_out[11]
+ sb_7__0_/chany_top_out[12] sb_7__0_/chany_top_out[13] sb_7__0_/chany_top_out[14]
+ sb_7__0_/chany_top_out[15] sb_7__0_/chany_top_out[16] sb_7__0_/chany_top_out[17]
+ sb_7__0_/chany_top_out[18] sb_7__0_/chany_top_out[19] sb_7__0_/chany_top_out[1]
+ sb_7__0_/chany_top_out[2] sb_7__0_/chany_top_out[3] sb_7__0_/chany_top_out[4] sb_7__0_/chany_top_out[5]
+ sb_7__0_/chany_top_out[6] sb_7__0_/chany_top_out[7] sb_7__0_/chany_top_out[8] sb_7__0_/chany_top_out[9]
+ sb_7__0_/clk_3_N_out sb_7__0_/clk_3_S_in sb_7__0_/left_bottom_grid_pin_11_ sb_7__0_/left_bottom_grid_pin_13_
+ sb_7__0_/left_bottom_grid_pin_15_ sb_7__0_/left_bottom_grid_pin_17_ sb_7__0_/left_bottom_grid_pin_1_
+ sb_7__0_/left_bottom_grid_pin_3_ sb_7__0_/left_bottom_grid_pin_5_ sb_7__0_/left_bottom_grid_pin_7_
+ sb_7__0_/left_bottom_grid_pin_9_ sb_7__0_/prog_clk_0_N_in sb_7__0_/prog_clk_3_N_out
+ sb_7__0_/prog_clk_3_S_in sb_7__0_/right_bottom_grid_pin_11_ sb_7__0_/right_bottom_grid_pin_13_
+ sb_7__0_/right_bottom_grid_pin_15_ sb_7__0_/right_bottom_grid_pin_17_ sb_7__0_/right_bottom_grid_pin_1_
+ sb_7__0_/right_bottom_grid_pin_3_ sb_7__0_/right_bottom_grid_pin_5_ sb_7__0_/right_bottom_grid_pin_7_
+ sb_7__0_/right_bottom_grid_pin_9_ sb_7__0_/top_left_grid_pin_42_ sb_7__0_/top_left_grid_pin_43_
+ sb_7__0_/top_left_grid_pin_44_ sb_7__0_/top_left_grid_pin_45_ sb_7__0_/top_left_grid_pin_46_
+ sb_7__0_/top_left_grid_pin_47_ sb_7__0_/top_left_grid_pin_48_ sb_7__0_/top_left_grid_pin_49_
+ sb_1__0_
Xsb_3__8_ sb_3__8_/SC_IN_BOT sb_3__8_/SC_OUT_BOT VGND VPWR sb_3__8_/bottom_left_grid_pin_42_
+ sb_3__8_/bottom_left_grid_pin_43_ sb_3__8_/bottom_left_grid_pin_44_ sb_3__8_/bottom_left_grid_pin_45_
+ sb_3__8_/bottom_left_grid_pin_46_ sb_3__8_/bottom_left_grid_pin_47_ sb_3__8_/bottom_left_grid_pin_48_
+ sb_3__8_/bottom_left_grid_pin_49_ sb_3__8_/ccff_head sb_3__8_/ccff_tail sb_3__8_/chanx_left_in[0]
+ sb_3__8_/chanx_left_in[10] sb_3__8_/chanx_left_in[11] sb_3__8_/chanx_left_in[12]
+ sb_3__8_/chanx_left_in[13] sb_3__8_/chanx_left_in[14] sb_3__8_/chanx_left_in[15]
+ sb_3__8_/chanx_left_in[16] sb_3__8_/chanx_left_in[17] sb_3__8_/chanx_left_in[18]
+ sb_3__8_/chanx_left_in[19] sb_3__8_/chanx_left_in[1] sb_3__8_/chanx_left_in[2] sb_3__8_/chanx_left_in[3]
+ sb_3__8_/chanx_left_in[4] sb_3__8_/chanx_left_in[5] sb_3__8_/chanx_left_in[6] sb_3__8_/chanx_left_in[7]
+ sb_3__8_/chanx_left_in[8] sb_3__8_/chanx_left_in[9] sb_3__8_/chanx_left_out[0] sb_3__8_/chanx_left_out[10]
+ sb_3__8_/chanx_left_out[11] sb_3__8_/chanx_left_out[12] sb_3__8_/chanx_left_out[13]
+ sb_3__8_/chanx_left_out[14] sb_3__8_/chanx_left_out[15] sb_3__8_/chanx_left_out[16]
+ sb_3__8_/chanx_left_out[17] sb_3__8_/chanx_left_out[18] sb_3__8_/chanx_left_out[19]
+ sb_3__8_/chanx_left_out[1] sb_3__8_/chanx_left_out[2] sb_3__8_/chanx_left_out[3]
+ sb_3__8_/chanx_left_out[4] sb_3__8_/chanx_left_out[5] sb_3__8_/chanx_left_out[6]
+ sb_3__8_/chanx_left_out[7] sb_3__8_/chanx_left_out[8] sb_3__8_/chanx_left_out[9]
+ sb_3__8_/chanx_right_in[0] sb_3__8_/chanx_right_in[10] sb_3__8_/chanx_right_in[11]
+ sb_3__8_/chanx_right_in[12] sb_3__8_/chanx_right_in[13] sb_3__8_/chanx_right_in[14]
+ sb_3__8_/chanx_right_in[15] sb_3__8_/chanx_right_in[16] sb_3__8_/chanx_right_in[17]
+ sb_3__8_/chanx_right_in[18] sb_3__8_/chanx_right_in[19] sb_3__8_/chanx_right_in[1]
+ sb_3__8_/chanx_right_in[2] sb_3__8_/chanx_right_in[3] sb_3__8_/chanx_right_in[4]
+ sb_3__8_/chanx_right_in[5] sb_3__8_/chanx_right_in[6] sb_3__8_/chanx_right_in[7]
+ sb_3__8_/chanx_right_in[8] sb_3__8_/chanx_right_in[9] cbx_4__8_/chanx_left_in[0]
+ cbx_4__8_/chanx_left_in[10] cbx_4__8_/chanx_left_in[11] cbx_4__8_/chanx_left_in[12]
+ cbx_4__8_/chanx_left_in[13] cbx_4__8_/chanx_left_in[14] cbx_4__8_/chanx_left_in[15]
+ cbx_4__8_/chanx_left_in[16] cbx_4__8_/chanx_left_in[17] cbx_4__8_/chanx_left_in[18]
+ cbx_4__8_/chanx_left_in[19] cbx_4__8_/chanx_left_in[1] cbx_4__8_/chanx_left_in[2]
+ cbx_4__8_/chanx_left_in[3] cbx_4__8_/chanx_left_in[4] cbx_4__8_/chanx_left_in[5]
+ cbx_4__8_/chanx_left_in[6] cbx_4__8_/chanx_left_in[7] cbx_4__8_/chanx_left_in[8]
+ cbx_4__8_/chanx_left_in[9] cby_3__8_/chany_top_out[0] cby_3__8_/chany_top_out[10]
+ cby_3__8_/chany_top_out[11] cby_3__8_/chany_top_out[12] cby_3__8_/chany_top_out[13]
+ cby_3__8_/chany_top_out[14] cby_3__8_/chany_top_out[15] cby_3__8_/chany_top_out[16]
+ cby_3__8_/chany_top_out[17] cby_3__8_/chany_top_out[18] cby_3__8_/chany_top_out[19]
+ cby_3__8_/chany_top_out[1] cby_3__8_/chany_top_out[2] cby_3__8_/chany_top_out[3]
+ cby_3__8_/chany_top_out[4] cby_3__8_/chany_top_out[5] cby_3__8_/chany_top_out[6]
+ cby_3__8_/chany_top_out[7] cby_3__8_/chany_top_out[8] cby_3__8_/chany_top_out[9]
+ cby_3__8_/chany_top_in[0] cby_3__8_/chany_top_in[10] cby_3__8_/chany_top_in[11]
+ cby_3__8_/chany_top_in[12] cby_3__8_/chany_top_in[13] cby_3__8_/chany_top_in[14]
+ cby_3__8_/chany_top_in[15] cby_3__8_/chany_top_in[16] cby_3__8_/chany_top_in[17]
+ cby_3__8_/chany_top_in[18] cby_3__8_/chany_top_in[19] cby_3__8_/chany_top_in[1]
+ cby_3__8_/chany_top_in[2] cby_3__8_/chany_top_in[3] cby_3__8_/chany_top_in[4] cby_3__8_/chany_top_in[5]
+ cby_3__8_/chany_top_in[6] cby_3__8_/chany_top_in[7] cby_3__8_/chany_top_in[8] cby_3__8_/chany_top_in[9]
+ sb_3__8_/left_bottom_grid_pin_34_ sb_3__8_/left_bottom_grid_pin_35_ sb_3__8_/left_bottom_grid_pin_36_
+ sb_3__8_/left_bottom_grid_pin_37_ sb_3__8_/left_bottom_grid_pin_38_ sb_3__8_/left_bottom_grid_pin_39_
+ sb_3__8_/left_bottom_grid_pin_40_ sb_3__8_/left_bottom_grid_pin_41_ sb_3__8_/left_top_grid_pin_1_
+ sb_3__8_/prog_clk_0_S_in sb_3__8_/right_bottom_grid_pin_34_ sb_3__8_/right_bottom_grid_pin_35_
+ sb_3__8_/right_bottom_grid_pin_36_ sb_3__8_/right_bottom_grid_pin_37_ sb_3__8_/right_bottom_grid_pin_38_
+ sb_3__8_/right_bottom_grid_pin_39_ sb_3__8_/right_bottom_grid_pin_40_ sb_3__8_/right_bottom_grid_pin_41_
+ sb_3__8_/right_top_grid_pin_1_ sb_1__2_
Xgrid_clb_2__3_ cbx_2__2_/SC_OUT_TOP grid_clb_2__3_/SC_OUT_BOT cbx_2__3_/SC_IN_BOT
+ cby_2__3_/Test_en_W_out grid_clb_2__3_/Test_en_E_out cby_2__3_/Test_en_W_out cby_1__3_/Test_en_W_in
+ VGND VPWR cbx_2__2_/REGIN_FEEDTHROUGH grid_clb_2__3_/bottom_width_0_height_0__pin_51_
+ cby_1__3_/ccff_tail cby_2__3_/ccff_head cbx_2__3_/clk_1_S_out cbx_2__3_/clk_1_S_out
+ cby_2__3_/prog_clk_0_W_in cbx_2__3_/prog_clk_1_S_out grid_clb_2__3_/prog_clk_0_N_out
+ cbx_2__3_/prog_clk_1_S_out cbx_2__2_/prog_clk_0_N_in grid_clb_2__3_/prog_clk_0_W_out
+ cby_2__3_/left_grid_pin_16_ cby_2__3_/left_grid_pin_17_ cby_2__3_/left_grid_pin_18_
+ cby_2__3_/left_grid_pin_19_ cby_2__3_/left_grid_pin_20_ cby_2__3_/left_grid_pin_21_
+ cby_2__3_/left_grid_pin_22_ cby_2__3_/left_grid_pin_23_ cby_2__3_/left_grid_pin_24_
+ cby_2__3_/left_grid_pin_25_ cby_2__3_/left_grid_pin_26_ cby_2__3_/left_grid_pin_27_
+ cby_2__3_/left_grid_pin_28_ cby_2__3_/left_grid_pin_29_ cby_2__3_/left_grid_pin_30_
+ cby_2__3_/left_grid_pin_31_ sb_2__2_/top_left_grid_pin_42_ sb_2__3_/bottom_left_grid_pin_42_
+ sb_2__2_/top_left_grid_pin_43_ sb_2__3_/bottom_left_grid_pin_43_ sb_2__2_/top_left_grid_pin_44_
+ sb_2__3_/bottom_left_grid_pin_44_ sb_2__2_/top_left_grid_pin_45_ sb_2__3_/bottom_left_grid_pin_45_
+ sb_2__2_/top_left_grid_pin_46_ sb_2__3_/bottom_left_grid_pin_46_ sb_2__2_/top_left_grid_pin_47_
+ sb_2__3_/bottom_left_grid_pin_47_ sb_2__2_/top_left_grid_pin_48_ sb_2__3_/bottom_left_grid_pin_48_
+ sb_2__2_/top_left_grid_pin_49_ sb_2__3_/bottom_left_grid_pin_49_ cbx_2__3_/bottom_grid_pin_0_
+ cbx_2__3_/bottom_grid_pin_10_ cbx_2__3_/bottom_grid_pin_11_ cbx_2__3_/bottom_grid_pin_12_
+ cbx_2__3_/bottom_grid_pin_13_ cbx_2__3_/bottom_grid_pin_14_ cbx_2__3_/bottom_grid_pin_15_
+ cbx_2__3_/bottom_grid_pin_1_ cbx_2__3_/bottom_grid_pin_2_ cbx_2__3_/REGOUT_FEEDTHROUGH
+ grid_clb_2__3_/top_width_0_height_0__pin_33_ sb_2__3_/left_bottom_grid_pin_34_ sb_1__3_/right_bottom_grid_pin_34_
+ sb_2__3_/left_bottom_grid_pin_35_ sb_1__3_/right_bottom_grid_pin_35_ sb_2__3_/left_bottom_grid_pin_36_
+ sb_1__3_/right_bottom_grid_pin_36_ sb_2__3_/left_bottom_grid_pin_37_ sb_1__3_/right_bottom_grid_pin_37_
+ sb_2__3_/left_bottom_grid_pin_38_ sb_1__3_/right_bottom_grid_pin_38_ sb_2__3_/left_bottom_grid_pin_39_
+ sb_1__3_/right_bottom_grid_pin_39_ cbx_2__3_/bottom_grid_pin_3_ sb_2__3_/left_bottom_grid_pin_40_
+ sb_1__3_/right_bottom_grid_pin_40_ sb_2__3_/left_bottom_grid_pin_41_ sb_1__3_/right_bottom_grid_pin_41_
+ cbx_2__3_/bottom_grid_pin_4_ cbx_2__3_/bottom_grid_pin_5_ cbx_2__3_/bottom_grid_pin_6_
+ cbx_2__3_/bottom_grid_pin_7_ cbx_2__3_/bottom_grid_pin_8_ cbx_2__3_/bottom_grid_pin_9_
+ grid_clb
Xsb_0__5_ VGND VPWR sb_0__5_/bottom_left_grid_pin_1_ sb_0__5_/ccff_head sb_0__5_/ccff_tail
+ sb_0__5_/chanx_right_in[0] sb_0__5_/chanx_right_in[10] sb_0__5_/chanx_right_in[11]
+ sb_0__5_/chanx_right_in[12] sb_0__5_/chanx_right_in[13] sb_0__5_/chanx_right_in[14]
+ sb_0__5_/chanx_right_in[15] sb_0__5_/chanx_right_in[16] sb_0__5_/chanx_right_in[17]
+ sb_0__5_/chanx_right_in[18] sb_0__5_/chanx_right_in[19] sb_0__5_/chanx_right_in[1]
+ sb_0__5_/chanx_right_in[2] sb_0__5_/chanx_right_in[3] sb_0__5_/chanx_right_in[4]
+ sb_0__5_/chanx_right_in[5] sb_0__5_/chanx_right_in[6] sb_0__5_/chanx_right_in[7]
+ sb_0__5_/chanx_right_in[8] sb_0__5_/chanx_right_in[9] cbx_1__5_/chanx_left_in[0]
+ cbx_1__5_/chanx_left_in[10] cbx_1__5_/chanx_left_in[11] cbx_1__5_/chanx_left_in[12]
+ cbx_1__5_/chanx_left_in[13] cbx_1__5_/chanx_left_in[14] cbx_1__5_/chanx_left_in[15]
+ cbx_1__5_/chanx_left_in[16] cbx_1__5_/chanx_left_in[17] cbx_1__5_/chanx_left_in[18]
+ cbx_1__5_/chanx_left_in[19] cbx_1__5_/chanx_left_in[1] cbx_1__5_/chanx_left_in[2]
+ cbx_1__5_/chanx_left_in[3] cbx_1__5_/chanx_left_in[4] cbx_1__5_/chanx_left_in[5]
+ cbx_1__5_/chanx_left_in[6] cbx_1__5_/chanx_left_in[7] cbx_1__5_/chanx_left_in[8]
+ cbx_1__5_/chanx_left_in[9] cby_0__5_/chany_top_out[0] cby_0__5_/chany_top_out[10]
+ cby_0__5_/chany_top_out[11] cby_0__5_/chany_top_out[12] cby_0__5_/chany_top_out[13]
+ cby_0__5_/chany_top_out[14] cby_0__5_/chany_top_out[15] cby_0__5_/chany_top_out[16]
+ cby_0__5_/chany_top_out[17] cby_0__5_/chany_top_out[18] cby_0__5_/chany_top_out[19]
+ cby_0__5_/chany_top_out[1] cby_0__5_/chany_top_out[2] cby_0__5_/chany_top_out[3]
+ cby_0__5_/chany_top_out[4] cby_0__5_/chany_top_out[5] cby_0__5_/chany_top_out[6]
+ cby_0__5_/chany_top_out[7] cby_0__5_/chany_top_out[8] cby_0__5_/chany_top_out[9]
+ cby_0__5_/chany_top_in[0] cby_0__5_/chany_top_in[10] cby_0__5_/chany_top_in[11]
+ cby_0__5_/chany_top_in[12] cby_0__5_/chany_top_in[13] cby_0__5_/chany_top_in[14]
+ cby_0__5_/chany_top_in[15] cby_0__5_/chany_top_in[16] cby_0__5_/chany_top_in[17]
+ cby_0__5_/chany_top_in[18] cby_0__5_/chany_top_in[19] cby_0__5_/chany_top_in[1]
+ cby_0__5_/chany_top_in[2] cby_0__5_/chany_top_in[3] cby_0__5_/chany_top_in[4] cby_0__5_/chany_top_in[5]
+ cby_0__5_/chany_top_in[6] cby_0__5_/chany_top_in[7] cby_0__5_/chany_top_in[8] cby_0__5_/chany_top_in[9]
+ sb_0__5_/chany_top_in[0] sb_0__5_/chany_top_in[10] sb_0__5_/chany_top_in[11] sb_0__5_/chany_top_in[12]
+ sb_0__5_/chany_top_in[13] sb_0__5_/chany_top_in[14] sb_0__5_/chany_top_in[15] sb_0__5_/chany_top_in[16]
+ sb_0__5_/chany_top_in[17] sb_0__5_/chany_top_in[18] sb_0__5_/chany_top_in[19] sb_0__5_/chany_top_in[1]
+ sb_0__5_/chany_top_in[2] sb_0__5_/chany_top_in[3] sb_0__5_/chany_top_in[4] sb_0__5_/chany_top_in[5]
+ sb_0__5_/chany_top_in[6] sb_0__5_/chany_top_in[7] sb_0__5_/chany_top_in[8] sb_0__5_/chany_top_in[9]
+ sb_0__5_/chany_top_out[0] sb_0__5_/chany_top_out[10] sb_0__5_/chany_top_out[11]
+ sb_0__5_/chany_top_out[12] sb_0__5_/chany_top_out[13] sb_0__5_/chany_top_out[14]
+ sb_0__5_/chany_top_out[15] sb_0__5_/chany_top_out[16] sb_0__5_/chany_top_out[17]
+ sb_0__5_/chany_top_out[18] sb_0__5_/chany_top_out[19] sb_0__5_/chany_top_out[1]
+ sb_0__5_/chany_top_out[2] sb_0__5_/chany_top_out[3] sb_0__5_/chany_top_out[4] sb_0__5_/chany_top_out[5]
+ sb_0__5_/chany_top_out[6] sb_0__5_/chany_top_out[7] sb_0__5_/chany_top_out[8] sb_0__5_/chany_top_out[9]
+ sb_0__5_/prog_clk_0_E_in sb_0__5_/right_bottom_grid_pin_34_ sb_0__5_/right_bottom_grid_pin_35_
+ sb_0__5_/right_bottom_grid_pin_36_ sb_0__5_/right_bottom_grid_pin_37_ sb_0__5_/right_bottom_grid_pin_38_
+ sb_0__5_/right_bottom_grid_pin_39_ sb_0__5_/right_bottom_grid_pin_40_ sb_0__5_/right_bottom_grid_pin_41_
+ sb_0__5_/top_left_grid_pin_1_ sb_0__1_
Xcby_6__4_ cby_6__4_/Test_en_W_in cby_6__4_/Test_en_E_out cby_6__4_/Test_en_N_out
+ cby_6__4_/Test_en_W_in cby_6__4_/Test_en_W_in cby_6__4_/Test_en_W_out VGND VPWR
+ cby_6__4_/ccff_head cby_6__4_/ccff_tail sb_6__3_/chany_top_out[0] sb_6__3_/chany_top_out[10]
+ sb_6__3_/chany_top_out[11] sb_6__3_/chany_top_out[12] sb_6__3_/chany_top_out[13]
+ sb_6__3_/chany_top_out[14] sb_6__3_/chany_top_out[15] sb_6__3_/chany_top_out[16]
+ sb_6__3_/chany_top_out[17] sb_6__3_/chany_top_out[18] sb_6__3_/chany_top_out[19]
+ sb_6__3_/chany_top_out[1] sb_6__3_/chany_top_out[2] sb_6__3_/chany_top_out[3] sb_6__3_/chany_top_out[4]
+ sb_6__3_/chany_top_out[5] sb_6__3_/chany_top_out[6] sb_6__3_/chany_top_out[7] sb_6__3_/chany_top_out[8]
+ sb_6__3_/chany_top_out[9] sb_6__3_/chany_top_in[0] sb_6__3_/chany_top_in[10] sb_6__3_/chany_top_in[11]
+ sb_6__3_/chany_top_in[12] sb_6__3_/chany_top_in[13] sb_6__3_/chany_top_in[14] sb_6__3_/chany_top_in[15]
+ sb_6__3_/chany_top_in[16] sb_6__3_/chany_top_in[17] sb_6__3_/chany_top_in[18] sb_6__3_/chany_top_in[19]
+ sb_6__3_/chany_top_in[1] sb_6__3_/chany_top_in[2] sb_6__3_/chany_top_in[3] sb_6__3_/chany_top_in[4]
+ sb_6__3_/chany_top_in[5] sb_6__3_/chany_top_in[6] sb_6__3_/chany_top_in[7] sb_6__3_/chany_top_in[8]
+ sb_6__3_/chany_top_in[9] cby_6__4_/chany_top_in[0] cby_6__4_/chany_top_in[10] cby_6__4_/chany_top_in[11]
+ cby_6__4_/chany_top_in[12] cby_6__4_/chany_top_in[13] cby_6__4_/chany_top_in[14]
+ cby_6__4_/chany_top_in[15] cby_6__4_/chany_top_in[16] cby_6__4_/chany_top_in[17]
+ cby_6__4_/chany_top_in[18] cby_6__4_/chany_top_in[19] cby_6__4_/chany_top_in[1]
+ cby_6__4_/chany_top_in[2] cby_6__4_/chany_top_in[3] cby_6__4_/chany_top_in[4] cby_6__4_/chany_top_in[5]
+ cby_6__4_/chany_top_in[6] cby_6__4_/chany_top_in[7] cby_6__4_/chany_top_in[8] cby_6__4_/chany_top_in[9]
+ cby_6__4_/chany_top_out[0] cby_6__4_/chany_top_out[10] cby_6__4_/chany_top_out[11]
+ cby_6__4_/chany_top_out[12] cby_6__4_/chany_top_out[13] cby_6__4_/chany_top_out[14]
+ cby_6__4_/chany_top_out[15] cby_6__4_/chany_top_out[16] cby_6__4_/chany_top_out[17]
+ cby_6__4_/chany_top_out[18] cby_6__4_/chany_top_out[19] cby_6__4_/chany_top_out[1]
+ cby_6__4_/chany_top_out[2] cby_6__4_/chany_top_out[3] cby_6__4_/chany_top_out[4]
+ cby_6__4_/chany_top_out[5] cby_6__4_/chany_top_out[6] cby_6__4_/chany_top_out[7]
+ cby_6__4_/chany_top_out[8] cby_6__4_/chany_top_out[9] cby_6__4_/clk_2_N_out cby_6__4_/clk_2_S_in
+ cby_6__4_/clk_2_S_out cby_6__4_/clk_3_N_out sb_6__4_/clk_3_S_out sb_6__3_/clk_3_N_in
+ cby_6__4_/left_grid_pin_16_ cby_6__4_/left_grid_pin_17_ cby_6__4_/left_grid_pin_18_
+ cby_6__4_/left_grid_pin_19_ cby_6__4_/left_grid_pin_20_ cby_6__4_/left_grid_pin_21_
+ cby_6__4_/left_grid_pin_22_ cby_6__4_/left_grid_pin_23_ cby_6__4_/left_grid_pin_24_
+ cby_6__4_/left_grid_pin_25_ cby_6__4_/left_grid_pin_26_ cby_6__4_/left_grid_pin_27_
+ cby_6__4_/left_grid_pin_28_ cby_6__4_/left_grid_pin_29_ cby_6__4_/left_grid_pin_30_
+ cby_6__4_/left_grid_pin_31_ cby_6__4_/prog_clk_0_N_out sb_6__3_/prog_clk_0_N_in
+ cby_6__4_/prog_clk_0_W_in cby_6__4_/prog_clk_2_N_out cby_6__4_/prog_clk_2_S_in cby_6__4_/prog_clk_2_S_out
+ cby_6__4_/prog_clk_3_N_out sb_6__4_/prog_clk_3_S_out sb_6__3_/prog_clk_3_N_in cby_1__1_
Xtie_array VGND VPWR tie_array/x[0] tie_array/x[1] tie_array/x[2] tie_array/x[3] tie_array/x[4]
+ tie_array/x[5] tie_array/x[6] tie_array/x[7] tie_array
Xgrid_clb_8__8_ cbx_8__7_/SC_OUT_TOP grid_clb_8__8_/SC_OUT_BOT cbx_8__8_/SC_IN_BOT
+ cby_7__8_/Test_en_E_out grid_clb_8__8_/Test_en_E_out cby_7__8_/Test_en_E_out grid_clb_8__8_/Test_en_W_out
+ VGND VPWR cbx_8__7_/REGIN_FEEDTHROUGH grid_clb_8__8_/bottom_width_0_height_0__pin_51_
+ cby_7__8_/ccff_tail cby_8__8_/ccff_head cbx_8__7_/clk_1_N_out cbx_8__7_/clk_1_N_out
+ cby_8__8_/prog_clk_0_W_in cbx_8__7_/prog_clk_1_N_out cbx_8__8_/prog_clk_0_S_in cbx_8__7_/prog_clk_1_N_out
+ cbx_8__7_/prog_clk_0_N_in grid_clb_8__8_/prog_clk_0_W_out cby_8__8_/left_grid_pin_16_
+ cby_8__8_/left_grid_pin_17_ cby_8__8_/left_grid_pin_18_ cby_8__8_/left_grid_pin_19_
+ cby_8__8_/left_grid_pin_20_ cby_8__8_/left_grid_pin_21_ cby_8__8_/left_grid_pin_22_
+ cby_8__8_/left_grid_pin_23_ cby_8__8_/left_grid_pin_24_ cby_8__8_/left_grid_pin_25_
+ cby_8__8_/left_grid_pin_26_ cby_8__8_/left_grid_pin_27_ cby_8__8_/left_grid_pin_28_
+ cby_8__8_/left_grid_pin_29_ cby_8__8_/left_grid_pin_30_ cby_8__8_/left_grid_pin_31_
+ sb_8__7_/top_left_grid_pin_42_ sb_8__8_/bottom_left_grid_pin_42_ sb_8__7_/top_left_grid_pin_43_
+ sb_8__8_/bottom_left_grid_pin_43_ sb_8__7_/top_left_grid_pin_44_ sb_8__8_/bottom_left_grid_pin_44_
+ sb_8__7_/top_left_grid_pin_45_ sb_8__8_/bottom_left_grid_pin_45_ sb_8__7_/top_left_grid_pin_46_
+ sb_8__8_/bottom_left_grid_pin_46_ sb_8__7_/top_left_grid_pin_47_ sb_8__8_/bottom_left_grid_pin_47_
+ sb_8__7_/top_left_grid_pin_48_ sb_8__8_/bottom_left_grid_pin_48_ sb_8__7_/top_left_grid_pin_49_
+ sb_8__8_/bottom_left_grid_pin_49_ cbx_8__8_/bottom_grid_pin_0_ cbx_8__8_/bottom_grid_pin_10_
+ cbx_8__8_/bottom_grid_pin_11_ cbx_8__8_/bottom_grid_pin_12_ cbx_8__8_/bottom_grid_pin_13_
+ cbx_8__8_/bottom_grid_pin_14_ cbx_8__8_/bottom_grid_pin_15_ cbx_8__8_/bottom_grid_pin_1_
+ cbx_8__8_/bottom_grid_pin_2_ tie_array/x[7] grid_clb_8__8_/top_width_0_height_0__pin_33_
+ sb_8__8_/left_bottom_grid_pin_34_ sb_7__8_/right_bottom_grid_pin_34_ sb_8__8_/left_bottom_grid_pin_35_
+ sb_7__8_/right_bottom_grid_pin_35_ sb_8__8_/left_bottom_grid_pin_36_ sb_7__8_/right_bottom_grid_pin_36_
+ sb_8__8_/left_bottom_grid_pin_37_ sb_7__8_/right_bottom_grid_pin_37_ sb_8__8_/left_bottom_grid_pin_38_
+ sb_7__8_/right_bottom_grid_pin_38_ sb_8__8_/left_bottom_grid_pin_39_ sb_7__8_/right_bottom_grid_pin_39_
+ cbx_8__8_/bottom_grid_pin_3_ sb_8__8_/left_bottom_grid_pin_40_ sb_7__8_/right_bottom_grid_pin_40_
+ sb_8__8_/left_bottom_grid_pin_41_ sb_7__8_/right_bottom_grid_pin_41_ cbx_8__8_/bottom_grid_pin_4_
+ cbx_8__8_/bottom_grid_pin_5_ cbx_8__8_/bottom_grid_pin_6_ cbx_8__8_/bottom_grid_pin_7_
+ cbx_8__8_/bottom_grid_pin_8_ cbx_8__8_/bottom_grid_pin_9_ grid_clb
Xcbx_6__5_ cbx_6__5_/REGIN_FEEDTHROUGH cbx_6__5_/REGOUT_FEEDTHROUGH cbx_6__5_/SC_IN_BOT
+ cbx_6__5_/SC_IN_TOP cbx_6__5_/SC_OUT_BOT cbx_6__5_/SC_OUT_TOP VGND VPWR cbx_6__5_/bottom_grid_pin_0_
+ cbx_6__5_/bottom_grid_pin_10_ cbx_6__5_/bottom_grid_pin_11_ cbx_6__5_/bottom_grid_pin_12_
+ cbx_6__5_/bottom_grid_pin_13_ cbx_6__5_/bottom_grid_pin_14_ cbx_6__5_/bottom_grid_pin_15_
+ cbx_6__5_/bottom_grid_pin_1_ cbx_6__5_/bottom_grid_pin_2_ cbx_6__5_/bottom_grid_pin_3_
+ cbx_6__5_/bottom_grid_pin_4_ cbx_6__5_/bottom_grid_pin_5_ cbx_6__5_/bottom_grid_pin_6_
+ cbx_6__5_/bottom_grid_pin_7_ cbx_6__5_/bottom_grid_pin_8_ cbx_6__5_/bottom_grid_pin_9_
+ sb_6__5_/ccff_tail sb_5__5_/ccff_head cbx_6__5_/chanx_left_in[0] cbx_6__5_/chanx_left_in[10]
+ cbx_6__5_/chanx_left_in[11] cbx_6__5_/chanx_left_in[12] cbx_6__5_/chanx_left_in[13]
+ cbx_6__5_/chanx_left_in[14] cbx_6__5_/chanx_left_in[15] cbx_6__5_/chanx_left_in[16]
+ cbx_6__5_/chanx_left_in[17] cbx_6__5_/chanx_left_in[18] cbx_6__5_/chanx_left_in[19]
+ cbx_6__5_/chanx_left_in[1] cbx_6__5_/chanx_left_in[2] cbx_6__5_/chanx_left_in[3]
+ cbx_6__5_/chanx_left_in[4] cbx_6__5_/chanx_left_in[5] cbx_6__5_/chanx_left_in[6]
+ cbx_6__5_/chanx_left_in[7] cbx_6__5_/chanx_left_in[8] cbx_6__5_/chanx_left_in[9]
+ sb_5__5_/chanx_right_in[0] sb_5__5_/chanx_right_in[10] sb_5__5_/chanx_right_in[11]
+ sb_5__5_/chanx_right_in[12] sb_5__5_/chanx_right_in[13] sb_5__5_/chanx_right_in[14]
+ sb_5__5_/chanx_right_in[15] sb_5__5_/chanx_right_in[16] sb_5__5_/chanx_right_in[17]
+ sb_5__5_/chanx_right_in[18] sb_5__5_/chanx_right_in[19] sb_5__5_/chanx_right_in[1]
+ sb_5__5_/chanx_right_in[2] sb_5__5_/chanx_right_in[3] sb_5__5_/chanx_right_in[4]
+ sb_5__5_/chanx_right_in[5] sb_5__5_/chanx_right_in[6] sb_5__5_/chanx_right_in[7]
+ sb_5__5_/chanx_right_in[8] sb_5__5_/chanx_right_in[9] sb_6__5_/chanx_left_out[0]
+ sb_6__5_/chanx_left_out[10] sb_6__5_/chanx_left_out[11] sb_6__5_/chanx_left_out[12]
+ sb_6__5_/chanx_left_out[13] sb_6__5_/chanx_left_out[14] sb_6__5_/chanx_left_out[15]
+ sb_6__5_/chanx_left_out[16] sb_6__5_/chanx_left_out[17] sb_6__5_/chanx_left_out[18]
+ sb_6__5_/chanx_left_out[19] sb_6__5_/chanx_left_out[1] sb_6__5_/chanx_left_out[2]
+ sb_6__5_/chanx_left_out[3] sb_6__5_/chanx_left_out[4] sb_6__5_/chanx_left_out[5]
+ sb_6__5_/chanx_left_out[6] sb_6__5_/chanx_left_out[7] sb_6__5_/chanx_left_out[8]
+ sb_6__5_/chanx_left_out[9] sb_6__5_/chanx_left_in[0] sb_6__5_/chanx_left_in[10]
+ sb_6__5_/chanx_left_in[11] sb_6__5_/chanx_left_in[12] sb_6__5_/chanx_left_in[13]
+ sb_6__5_/chanx_left_in[14] sb_6__5_/chanx_left_in[15] sb_6__5_/chanx_left_in[16]
+ sb_6__5_/chanx_left_in[17] sb_6__5_/chanx_left_in[18] sb_6__5_/chanx_left_in[19]
+ sb_6__5_/chanx_left_in[1] sb_6__5_/chanx_left_in[2] sb_6__5_/chanx_left_in[3] sb_6__5_/chanx_left_in[4]
+ sb_6__5_/chanx_left_in[5] sb_6__5_/chanx_left_in[6] sb_6__5_/chanx_left_in[7] sb_6__5_/chanx_left_in[8]
+ sb_6__5_/chanx_left_in[9] cbx_6__5_/clk_1_N_out cbx_6__5_/clk_1_S_out sb_5__5_/clk_1_E_out
+ cbx_6__5_/clk_2_E_out cbx_6__5_/clk_2_W_in cbx_6__5_/clk_2_W_out cbx_6__5_/clk_3_E_out
+ cbx_6__5_/clk_3_W_in cbx_6__5_/clk_3_W_out cbx_6__5_/prog_clk_0_N_in cbx_6__5_/prog_clk_0_W_out
+ cbx_6__5_/prog_clk_1_N_out cbx_6__5_/prog_clk_1_S_out sb_5__5_/prog_clk_1_E_out
+ cbx_6__5_/prog_clk_2_E_out cbx_6__5_/prog_clk_2_W_in cbx_6__5_/prog_clk_2_W_out
+ cbx_6__5_/prog_clk_3_E_out cbx_6__5_/prog_clk_3_W_in cbx_6__5_/prog_clk_3_W_out
+ cbx_1__1_
Xcby_3__1_ cby_3__1_/Test_en_W_in cby_3__1_/Test_en_E_out cby_3__1_/Test_en_N_out
+ cby_3__1_/Test_en_W_in cby_3__1_/Test_en_W_in cby_3__1_/Test_en_W_out VGND VPWR
+ cby_3__1_/ccff_head cby_3__1_/ccff_tail sb_3__0_/chany_top_out[0] sb_3__0_/chany_top_out[10]
+ sb_3__0_/chany_top_out[11] sb_3__0_/chany_top_out[12] sb_3__0_/chany_top_out[13]
+ sb_3__0_/chany_top_out[14] sb_3__0_/chany_top_out[15] sb_3__0_/chany_top_out[16]
+ sb_3__0_/chany_top_out[17] sb_3__0_/chany_top_out[18] sb_3__0_/chany_top_out[19]
+ sb_3__0_/chany_top_out[1] sb_3__0_/chany_top_out[2] sb_3__0_/chany_top_out[3] sb_3__0_/chany_top_out[4]
+ sb_3__0_/chany_top_out[5] sb_3__0_/chany_top_out[6] sb_3__0_/chany_top_out[7] sb_3__0_/chany_top_out[8]
+ sb_3__0_/chany_top_out[9] sb_3__0_/chany_top_in[0] sb_3__0_/chany_top_in[10] sb_3__0_/chany_top_in[11]
+ sb_3__0_/chany_top_in[12] sb_3__0_/chany_top_in[13] sb_3__0_/chany_top_in[14] sb_3__0_/chany_top_in[15]
+ sb_3__0_/chany_top_in[16] sb_3__0_/chany_top_in[17] sb_3__0_/chany_top_in[18] sb_3__0_/chany_top_in[19]
+ sb_3__0_/chany_top_in[1] sb_3__0_/chany_top_in[2] sb_3__0_/chany_top_in[3] sb_3__0_/chany_top_in[4]
+ sb_3__0_/chany_top_in[5] sb_3__0_/chany_top_in[6] sb_3__0_/chany_top_in[7] sb_3__0_/chany_top_in[8]
+ sb_3__0_/chany_top_in[9] cby_3__1_/chany_top_in[0] cby_3__1_/chany_top_in[10] cby_3__1_/chany_top_in[11]
+ cby_3__1_/chany_top_in[12] cby_3__1_/chany_top_in[13] cby_3__1_/chany_top_in[14]
+ cby_3__1_/chany_top_in[15] cby_3__1_/chany_top_in[16] cby_3__1_/chany_top_in[17]
+ cby_3__1_/chany_top_in[18] cby_3__1_/chany_top_in[19] cby_3__1_/chany_top_in[1]
+ cby_3__1_/chany_top_in[2] cby_3__1_/chany_top_in[3] cby_3__1_/chany_top_in[4] cby_3__1_/chany_top_in[5]
+ cby_3__1_/chany_top_in[6] cby_3__1_/chany_top_in[7] cby_3__1_/chany_top_in[8] cby_3__1_/chany_top_in[9]
+ cby_3__1_/chany_top_out[0] cby_3__1_/chany_top_out[10] cby_3__1_/chany_top_out[11]
+ cby_3__1_/chany_top_out[12] cby_3__1_/chany_top_out[13] cby_3__1_/chany_top_out[14]
+ cby_3__1_/chany_top_out[15] cby_3__1_/chany_top_out[16] cby_3__1_/chany_top_out[17]
+ cby_3__1_/chany_top_out[18] cby_3__1_/chany_top_out[19] cby_3__1_/chany_top_out[1]
+ cby_3__1_/chany_top_out[2] cby_3__1_/chany_top_out[3] cby_3__1_/chany_top_out[4]
+ cby_3__1_/chany_top_out[5] cby_3__1_/chany_top_out[6] cby_3__1_/chany_top_out[7]
+ cby_3__1_/chany_top_out[8] cby_3__1_/chany_top_out[9] cby_3__1_/clk_2_N_out cby_3__1_/clk_2_S_in
+ cby_3__1_/clk_2_S_out cby_3__1_/clk_3_N_out cby_3__1_/clk_3_S_in cby_3__1_/clk_3_S_out
+ cby_3__1_/left_grid_pin_16_ cby_3__1_/left_grid_pin_17_ cby_3__1_/left_grid_pin_18_
+ cby_3__1_/left_grid_pin_19_ cby_3__1_/left_grid_pin_20_ cby_3__1_/left_grid_pin_21_
+ cby_3__1_/left_grid_pin_22_ cby_3__1_/left_grid_pin_23_ cby_3__1_/left_grid_pin_24_
+ cby_3__1_/left_grid_pin_25_ cby_3__1_/left_grid_pin_26_ cby_3__1_/left_grid_pin_27_
+ cby_3__1_/left_grid_pin_28_ cby_3__1_/left_grid_pin_29_ cby_3__1_/left_grid_pin_30_
+ cby_3__1_/left_grid_pin_31_ cby_3__1_/prog_clk_0_N_out sb_3__0_/prog_clk_0_N_in
+ cby_3__1_/prog_clk_0_W_in cby_3__1_/prog_clk_2_N_out cby_3__1_/prog_clk_2_S_in cby_3__1_/prog_clk_2_S_out
+ cby_3__1_/prog_clk_3_N_out cby_3__1_/prog_clk_3_S_in cby_3__1_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_5__5_ cbx_5__5_/SC_OUT_BOT cbx_5__4_/SC_IN_TOP grid_clb_5__5_/SC_OUT_TOP
+ cby_4__5_/Test_en_E_out cby_5__5_/Test_en_W_in cby_4__5_/Test_en_E_out grid_clb_5__5_/Test_en_W_out
+ VGND VPWR cbx_5__4_/REGIN_FEEDTHROUGH grid_clb_5__5_/bottom_width_0_height_0__pin_51_
+ cby_4__5_/ccff_tail cby_5__5_/ccff_head cbx_5__5_/clk_1_S_out cbx_5__5_/clk_1_S_out
+ cby_5__5_/prog_clk_0_W_in cbx_5__5_/prog_clk_1_S_out grid_clb_5__5_/prog_clk_0_N_out
+ cbx_5__5_/prog_clk_1_S_out cbx_5__4_/prog_clk_0_N_in grid_clb_5__5_/prog_clk_0_W_out
+ cby_5__5_/left_grid_pin_16_ cby_5__5_/left_grid_pin_17_ cby_5__5_/left_grid_pin_18_
+ cby_5__5_/left_grid_pin_19_ cby_5__5_/left_grid_pin_20_ cby_5__5_/left_grid_pin_21_
+ cby_5__5_/left_grid_pin_22_ cby_5__5_/left_grid_pin_23_ cby_5__5_/left_grid_pin_24_
+ cby_5__5_/left_grid_pin_25_ cby_5__5_/left_grid_pin_26_ cby_5__5_/left_grid_pin_27_
+ cby_5__5_/left_grid_pin_28_ cby_5__5_/left_grid_pin_29_ cby_5__5_/left_grid_pin_30_
+ cby_5__5_/left_grid_pin_31_ sb_5__4_/top_left_grid_pin_42_ sb_5__5_/bottom_left_grid_pin_42_
+ sb_5__4_/top_left_grid_pin_43_ sb_5__5_/bottom_left_grid_pin_43_ sb_5__4_/top_left_grid_pin_44_
+ sb_5__5_/bottom_left_grid_pin_44_ sb_5__4_/top_left_grid_pin_45_ sb_5__5_/bottom_left_grid_pin_45_
+ sb_5__4_/top_left_grid_pin_46_ sb_5__5_/bottom_left_grid_pin_46_ sb_5__4_/top_left_grid_pin_47_
+ sb_5__5_/bottom_left_grid_pin_47_ sb_5__4_/top_left_grid_pin_48_ sb_5__5_/bottom_left_grid_pin_48_
+ sb_5__4_/top_left_grid_pin_49_ sb_5__5_/bottom_left_grid_pin_49_ cbx_5__5_/bottom_grid_pin_0_
+ cbx_5__5_/bottom_grid_pin_10_ cbx_5__5_/bottom_grid_pin_11_ cbx_5__5_/bottom_grid_pin_12_
+ cbx_5__5_/bottom_grid_pin_13_ cbx_5__5_/bottom_grid_pin_14_ cbx_5__5_/bottom_grid_pin_15_
+ cbx_5__5_/bottom_grid_pin_1_ cbx_5__5_/bottom_grid_pin_2_ cbx_5__5_/REGOUT_FEEDTHROUGH
+ grid_clb_5__5_/top_width_0_height_0__pin_33_ sb_5__5_/left_bottom_grid_pin_34_ sb_4__5_/right_bottom_grid_pin_34_
+ sb_5__5_/left_bottom_grid_pin_35_ sb_4__5_/right_bottom_grid_pin_35_ sb_5__5_/left_bottom_grid_pin_36_
+ sb_4__5_/right_bottom_grid_pin_36_ sb_5__5_/left_bottom_grid_pin_37_ sb_4__5_/right_bottom_grid_pin_37_
+ sb_5__5_/left_bottom_grid_pin_38_ sb_4__5_/right_bottom_grid_pin_38_ sb_5__5_/left_bottom_grid_pin_39_
+ sb_4__5_/right_bottom_grid_pin_39_ cbx_5__5_/bottom_grid_pin_3_ sb_5__5_/left_bottom_grid_pin_40_
+ sb_4__5_/right_bottom_grid_pin_40_ sb_5__5_/left_bottom_grid_pin_41_ sb_4__5_/right_bottom_grid_pin_41_
+ cbx_5__5_/bottom_grid_pin_4_ cbx_5__5_/bottom_grid_pin_5_ cbx_5__5_/bottom_grid_pin_6_
+ cbx_5__5_/bottom_grid_pin_7_ cbx_5__5_/bottom_grid_pin_8_ cbx_5__5_/bottom_grid_pin_9_
+ grid_clb
Xgrid_clb_2__2_ cbx_2__1_/SC_OUT_TOP grid_clb_2__2_/SC_OUT_BOT cbx_2__2_/SC_IN_BOT
+ cby_2__2_/Test_en_W_out grid_clb_2__2_/Test_en_E_out cby_2__2_/Test_en_W_out cby_1__2_/Test_en_W_in
+ VGND VPWR cbx_2__1_/REGIN_FEEDTHROUGH grid_clb_2__2_/bottom_width_0_height_0__pin_51_
+ cby_1__2_/ccff_tail cby_2__2_/ccff_head cbx_2__1_/clk_1_N_out cbx_2__1_/clk_1_N_out
+ cby_2__2_/prog_clk_0_W_in cbx_2__1_/prog_clk_1_N_out grid_clb_2__2_/prog_clk_0_N_out
+ cbx_2__1_/prog_clk_1_N_out cbx_2__1_/prog_clk_0_N_in grid_clb_2__2_/prog_clk_0_W_out
+ cby_2__2_/left_grid_pin_16_ cby_2__2_/left_grid_pin_17_ cby_2__2_/left_grid_pin_18_
+ cby_2__2_/left_grid_pin_19_ cby_2__2_/left_grid_pin_20_ cby_2__2_/left_grid_pin_21_
+ cby_2__2_/left_grid_pin_22_ cby_2__2_/left_grid_pin_23_ cby_2__2_/left_grid_pin_24_
+ cby_2__2_/left_grid_pin_25_ cby_2__2_/left_grid_pin_26_ cby_2__2_/left_grid_pin_27_
+ cby_2__2_/left_grid_pin_28_ cby_2__2_/left_grid_pin_29_ cby_2__2_/left_grid_pin_30_
+ cby_2__2_/left_grid_pin_31_ sb_2__1_/top_left_grid_pin_42_ sb_2__2_/bottom_left_grid_pin_42_
+ sb_2__1_/top_left_grid_pin_43_ sb_2__2_/bottom_left_grid_pin_43_ sb_2__1_/top_left_grid_pin_44_
+ sb_2__2_/bottom_left_grid_pin_44_ sb_2__1_/top_left_grid_pin_45_ sb_2__2_/bottom_left_grid_pin_45_
+ sb_2__1_/top_left_grid_pin_46_ sb_2__2_/bottom_left_grid_pin_46_ sb_2__1_/top_left_grid_pin_47_
+ sb_2__2_/bottom_left_grid_pin_47_ sb_2__1_/top_left_grid_pin_48_ sb_2__2_/bottom_left_grid_pin_48_
+ sb_2__1_/top_left_grid_pin_49_ sb_2__2_/bottom_left_grid_pin_49_ cbx_2__2_/bottom_grid_pin_0_
+ cbx_2__2_/bottom_grid_pin_10_ cbx_2__2_/bottom_grid_pin_11_ cbx_2__2_/bottom_grid_pin_12_
+ cbx_2__2_/bottom_grid_pin_13_ cbx_2__2_/bottom_grid_pin_14_ cbx_2__2_/bottom_grid_pin_15_
+ cbx_2__2_/bottom_grid_pin_1_ cbx_2__2_/bottom_grid_pin_2_ cbx_2__2_/REGOUT_FEEDTHROUGH
+ grid_clb_2__2_/top_width_0_height_0__pin_33_ sb_2__2_/left_bottom_grid_pin_34_ sb_1__2_/right_bottom_grid_pin_34_
+ sb_2__2_/left_bottom_grid_pin_35_ sb_1__2_/right_bottom_grid_pin_35_ sb_2__2_/left_bottom_grid_pin_36_
+ sb_1__2_/right_bottom_grid_pin_36_ sb_2__2_/left_bottom_grid_pin_37_ sb_1__2_/right_bottom_grid_pin_37_
+ sb_2__2_/left_bottom_grid_pin_38_ sb_1__2_/right_bottom_grid_pin_38_ sb_2__2_/left_bottom_grid_pin_39_
+ sb_1__2_/right_bottom_grid_pin_39_ cbx_2__2_/bottom_grid_pin_3_ sb_2__2_/left_bottom_grid_pin_40_
+ sb_1__2_/right_bottom_grid_pin_40_ sb_2__2_/left_bottom_grid_pin_41_ sb_1__2_/right_bottom_grid_pin_41_
+ cbx_2__2_/bottom_grid_pin_4_ cbx_2__2_/bottom_grid_pin_5_ cbx_2__2_/bottom_grid_pin_6_
+ cbx_2__2_/bottom_grid_pin_7_ cbx_2__2_/bottom_grid_pin_8_ cbx_2__2_/bottom_grid_pin_9_
+ grid_clb
Xcbx_3__2_ cbx_3__2_/REGIN_FEEDTHROUGH cbx_3__2_/REGOUT_FEEDTHROUGH cbx_3__2_/SC_IN_BOT
+ cbx_3__2_/SC_IN_TOP cbx_3__2_/SC_OUT_BOT cbx_3__2_/SC_OUT_TOP VGND VPWR cbx_3__2_/bottom_grid_pin_0_
+ cbx_3__2_/bottom_grid_pin_10_ cbx_3__2_/bottom_grid_pin_11_ cbx_3__2_/bottom_grid_pin_12_
+ cbx_3__2_/bottom_grid_pin_13_ cbx_3__2_/bottom_grid_pin_14_ cbx_3__2_/bottom_grid_pin_15_
+ cbx_3__2_/bottom_grid_pin_1_ cbx_3__2_/bottom_grid_pin_2_ cbx_3__2_/bottom_grid_pin_3_
+ cbx_3__2_/bottom_grid_pin_4_ cbx_3__2_/bottom_grid_pin_5_ cbx_3__2_/bottom_grid_pin_6_
+ cbx_3__2_/bottom_grid_pin_7_ cbx_3__2_/bottom_grid_pin_8_ cbx_3__2_/bottom_grid_pin_9_
+ sb_3__2_/ccff_tail sb_2__2_/ccff_head cbx_3__2_/chanx_left_in[0] cbx_3__2_/chanx_left_in[10]
+ cbx_3__2_/chanx_left_in[11] cbx_3__2_/chanx_left_in[12] cbx_3__2_/chanx_left_in[13]
+ cbx_3__2_/chanx_left_in[14] cbx_3__2_/chanx_left_in[15] cbx_3__2_/chanx_left_in[16]
+ cbx_3__2_/chanx_left_in[17] cbx_3__2_/chanx_left_in[18] cbx_3__2_/chanx_left_in[19]
+ cbx_3__2_/chanx_left_in[1] cbx_3__2_/chanx_left_in[2] cbx_3__2_/chanx_left_in[3]
+ cbx_3__2_/chanx_left_in[4] cbx_3__2_/chanx_left_in[5] cbx_3__2_/chanx_left_in[6]
+ cbx_3__2_/chanx_left_in[7] cbx_3__2_/chanx_left_in[8] cbx_3__2_/chanx_left_in[9]
+ sb_2__2_/chanx_right_in[0] sb_2__2_/chanx_right_in[10] sb_2__2_/chanx_right_in[11]
+ sb_2__2_/chanx_right_in[12] sb_2__2_/chanx_right_in[13] sb_2__2_/chanx_right_in[14]
+ sb_2__2_/chanx_right_in[15] sb_2__2_/chanx_right_in[16] sb_2__2_/chanx_right_in[17]
+ sb_2__2_/chanx_right_in[18] sb_2__2_/chanx_right_in[19] sb_2__2_/chanx_right_in[1]
+ sb_2__2_/chanx_right_in[2] sb_2__2_/chanx_right_in[3] sb_2__2_/chanx_right_in[4]
+ sb_2__2_/chanx_right_in[5] sb_2__2_/chanx_right_in[6] sb_2__2_/chanx_right_in[7]
+ sb_2__2_/chanx_right_in[8] sb_2__2_/chanx_right_in[9] sb_3__2_/chanx_left_out[0]
+ sb_3__2_/chanx_left_out[10] sb_3__2_/chanx_left_out[11] sb_3__2_/chanx_left_out[12]
+ sb_3__2_/chanx_left_out[13] sb_3__2_/chanx_left_out[14] sb_3__2_/chanx_left_out[15]
+ sb_3__2_/chanx_left_out[16] sb_3__2_/chanx_left_out[17] sb_3__2_/chanx_left_out[18]
+ sb_3__2_/chanx_left_out[19] sb_3__2_/chanx_left_out[1] sb_3__2_/chanx_left_out[2]
+ sb_3__2_/chanx_left_out[3] sb_3__2_/chanx_left_out[4] sb_3__2_/chanx_left_out[5]
+ sb_3__2_/chanx_left_out[6] sb_3__2_/chanx_left_out[7] sb_3__2_/chanx_left_out[8]
+ sb_3__2_/chanx_left_out[9] sb_3__2_/chanx_left_in[0] sb_3__2_/chanx_left_in[10]
+ sb_3__2_/chanx_left_in[11] sb_3__2_/chanx_left_in[12] sb_3__2_/chanx_left_in[13]
+ sb_3__2_/chanx_left_in[14] sb_3__2_/chanx_left_in[15] sb_3__2_/chanx_left_in[16]
+ sb_3__2_/chanx_left_in[17] sb_3__2_/chanx_left_in[18] sb_3__2_/chanx_left_in[19]
+ sb_3__2_/chanx_left_in[1] sb_3__2_/chanx_left_in[2] sb_3__2_/chanx_left_in[3] sb_3__2_/chanx_left_in[4]
+ sb_3__2_/chanx_left_in[5] sb_3__2_/chanx_left_in[6] sb_3__2_/chanx_left_in[7] sb_3__2_/chanx_left_in[8]
+ sb_3__2_/chanx_left_in[9] cbx_3__2_/clk_1_N_out cbx_3__2_/clk_1_S_out cbx_3__2_/clk_1_W_in
+ sb_3__2_/clk_2_N_in sb_2__2_/clk_2_E_out cbx_3__2_/clk_2_W_out cbx_3__2_/clk_3_E_out
+ cbx_3__2_/clk_3_W_in cbx_3__2_/clk_3_W_out cbx_3__2_/prog_clk_0_N_in cbx_3__2_/prog_clk_0_W_out
+ cbx_3__2_/prog_clk_1_N_out cbx_3__2_/prog_clk_1_S_out cbx_3__2_/prog_clk_1_W_in
+ sb_3__2_/prog_clk_2_N_in sb_2__2_/prog_clk_2_E_out cbx_3__2_/prog_clk_2_W_out cbx_3__2_/prog_clk_3_E_out
+ cbx_3__2_/prog_clk_3_W_in cbx_3__2_/prog_clk_3_W_out cbx_1__1_
Xsb_3__7_ sb_3__7_/Test_en_N_out sb_3__7_/Test_en_S_in VGND VPWR sb_3__7_/bottom_left_grid_pin_42_
+ sb_3__7_/bottom_left_grid_pin_43_ sb_3__7_/bottom_left_grid_pin_44_ sb_3__7_/bottom_left_grid_pin_45_
+ sb_3__7_/bottom_left_grid_pin_46_ sb_3__7_/bottom_left_grid_pin_47_ sb_3__7_/bottom_left_grid_pin_48_
+ sb_3__7_/bottom_left_grid_pin_49_ sb_3__7_/ccff_head sb_3__7_/ccff_tail sb_3__7_/chanx_left_in[0]
+ sb_3__7_/chanx_left_in[10] sb_3__7_/chanx_left_in[11] sb_3__7_/chanx_left_in[12]
+ sb_3__7_/chanx_left_in[13] sb_3__7_/chanx_left_in[14] sb_3__7_/chanx_left_in[15]
+ sb_3__7_/chanx_left_in[16] sb_3__7_/chanx_left_in[17] sb_3__7_/chanx_left_in[18]
+ sb_3__7_/chanx_left_in[19] sb_3__7_/chanx_left_in[1] sb_3__7_/chanx_left_in[2] sb_3__7_/chanx_left_in[3]
+ sb_3__7_/chanx_left_in[4] sb_3__7_/chanx_left_in[5] sb_3__7_/chanx_left_in[6] sb_3__7_/chanx_left_in[7]
+ sb_3__7_/chanx_left_in[8] sb_3__7_/chanx_left_in[9] sb_3__7_/chanx_left_out[0] sb_3__7_/chanx_left_out[10]
+ sb_3__7_/chanx_left_out[11] sb_3__7_/chanx_left_out[12] sb_3__7_/chanx_left_out[13]
+ sb_3__7_/chanx_left_out[14] sb_3__7_/chanx_left_out[15] sb_3__7_/chanx_left_out[16]
+ sb_3__7_/chanx_left_out[17] sb_3__7_/chanx_left_out[18] sb_3__7_/chanx_left_out[19]
+ sb_3__7_/chanx_left_out[1] sb_3__7_/chanx_left_out[2] sb_3__7_/chanx_left_out[3]
+ sb_3__7_/chanx_left_out[4] sb_3__7_/chanx_left_out[5] sb_3__7_/chanx_left_out[6]
+ sb_3__7_/chanx_left_out[7] sb_3__7_/chanx_left_out[8] sb_3__7_/chanx_left_out[9]
+ sb_3__7_/chanx_right_in[0] sb_3__7_/chanx_right_in[10] sb_3__7_/chanx_right_in[11]
+ sb_3__7_/chanx_right_in[12] sb_3__7_/chanx_right_in[13] sb_3__7_/chanx_right_in[14]
+ sb_3__7_/chanx_right_in[15] sb_3__7_/chanx_right_in[16] sb_3__7_/chanx_right_in[17]
+ sb_3__7_/chanx_right_in[18] sb_3__7_/chanx_right_in[19] sb_3__7_/chanx_right_in[1]
+ sb_3__7_/chanx_right_in[2] sb_3__7_/chanx_right_in[3] sb_3__7_/chanx_right_in[4]
+ sb_3__7_/chanx_right_in[5] sb_3__7_/chanx_right_in[6] sb_3__7_/chanx_right_in[7]
+ sb_3__7_/chanx_right_in[8] sb_3__7_/chanx_right_in[9] cbx_4__7_/chanx_left_in[0]
+ cbx_4__7_/chanx_left_in[10] cbx_4__7_/chanx_left_in[11] cbx_4__7_/chanx_left_in[12]
+ cbx_4__7_/chanx_left_in[13] cbx_4__7_/chanx_left_in[14] cbx_4__7_/chanx_left_in[15]
+ cbx_4__7_/chanx_left_in[16] cbx_4__7_/chanx_left_in[17] cbx_4__7_/chanx_left_in[18]
+ cbx_4__7_/chanx_left_in[19] cbx_4__7_/chanx_left_in[1] cbx_4__7_/chanx_left_in[2]
+ cbx_4__7_/chanx_left_in[3] cbx_4__7_/chanx_left_in[4] cbx_4__7_/chanx_left_in[5]
+ cbx_4__7_/chanx_left_in[6] cbx_4__7_/chanx_left_in[7] cbx_4__7_/chanx_left_in[8]
+ cbx_4__7_/chanx_left_in[9] cby_3__7_/chany_top_out[0] cby_3__7_/chany_top_out[10]
+ cby_3__7_/chany_top_out[11] cby_3__7_/chany_top_out[12] cby_3__7_/chany_top_out[13]
+ cby_3__7_/chany_top_out[14] cby_3__7_/chany_top_out[15] cby_3__7_/chany_top_out[16]
+ cby_3__7_/chany_top_out[17] cby_3__7_/chany_top_out[18] cby_3__7_/chany_top_out[19]
+ cby_3__7_/chany_top_out[1] cby_3__7_/chany_top_out[2] cby_3__7_/chany_top_out[3]
+ cby_3__7_/chany_top_out[4] cby_3__7_/chany_top_out[5] cby_3__7_/chany_top_out[6]
+ cby_3__7_/chany_top_out[7] cby_3__7_/chany_top_out[8] cby_3__7_/chany_top_out[9]
+ cby_3__7_/chany_top_in[0] cby_3__7_/chany_top_in[10] cby_3__7_/chany_top_in[11]
+ cby_3__7_/chany_top_in[12] cby_3__7_/chany_top_in[13] cby_3__7_/chany_top_in[14]
+ cby_3__7_/chany_top_in[15] cby_3__7_/chany_top_in[16] cby_3__7_/chany_top_in[17]
+ cby_3__7_/chany_top_in[18] cby_3__7_/chany_top_in[19] cby_3__7_/chany_top_in[1]
+ cby_3__7_/chany_top_in[2] cby_3__7_/chany_top_in[3] cby_3__7_/chany_top_in[4] cby_3__7_/chany_top_in[5]
+ cby_3__7_/chany_top_in[6] cby_3__7_/chany_top_in[7] cby_3__7_/chany_top_in[8] cby_3__7_/chany_top_in[9]
+ sb_3__7_/chany_top_in[0] sb_3__7_/chany_top_in[10] sb_3__7_/chany_top_in[11] sb_3__7_/chany_top_in[12]
+ sb_3__7_/chany_top_in[13] sb_3__7_/chany_top_in[14] sb_3__7_/chany_top_in[15] sb_3__7_/chany_top_in[16]
+ sb_3__7_/chany_top_in[17] sb_3__7_/chany_top_in[18] sb_3__7_/chany_top_in[19] sb_3__7_/chany_top_in[1]
+ sb_3__7_/chany_top_in[2] sb_3__7_/chany_top_in[3] sb_3__7_/chany_top_in[4] sb_3__7_/chany_top_in[5]
+ sb_3__7_/chany_top_in[6] sb_3__7_/chany_top_in[7] sb_3__7_/chany_top_in[8] sb_3__7_/chany_top_in[9]
+ sb_3__7_/chany_top_out[0] sb_3__7_/chany_top_out[10] sb_3__7_/chany_top_out[11]
+ sb_3__7_/chany_top_out[12] sb_3__7_/chany_top_out[13] sb_3__7_/chany_top_out[14]
+ sb_3__7_/chany_top_out[15] sb_3__7_/chany_top_out[16] sb_3__7_/chany_top_out[17]
+ sb_3__7_/chany_top_out[18] sb_3__7_/chany_top_out[19] sb_3__7_/chany_top_out[1]
+ sb_3__7_/chany_top_out[2] sb_3__7_/chany_top_out[3] sb_3__7_/chany_top_out[4] sb_3__7_/chany_top_out[5]
+ sb_3__7_/chany_top_out[6] sb_3__7_/chany_top_out[7] sb_3__7_/chany_top_out[8] sb_3__7_/chany_top_out[9]
+ sb_3__7_/clk_1_E_out sb_3__7_/clk_1_N_in sb_3__7_/clk_1_W_out sb_3__7_/clk_2_E_out
+ sb_3__7_/clk_2_N_in sb_3__7_/clk_2_N_out sb_3__7_/clk_2_S_out sb_3__7_/clk_2_W_out
+ sb_3__7_/clk_3_E_out sb_3__7_/clk_3_N_in sb_3__7_/clk_3_N_out sb_3__7_/clk_3_S_out
+ sb_3__7_/clk_3_W_out sb_3__7_/left_bottom_grid_pin_34_ sb_3__7_/left_bottom_grid_pin_35_
+ sb_3__7_/left_bottom_grid_pin_36_ sb_3__7_/left_bottom_grid_pin_37_ sb_3__7_/left_bottom_grid_pin_38_
+ sb_3__7_/left_bottom_grid_pin_39_ sb_3__7_/left_bottom_grid_pin_40_ sb_3__7_/left_bottom_grid_pin_41_
+ sb_3__7_/prog_clk_0_N_in sb_3__7_/prog_clk_1_E_out sb_3__7_/prog_clk_1_N_in sb_3__7_/prog_clk_1_W_out
+ sb_3__7_/prog_clk_2_E_out sb_3__7_/prog_clk_2_N_in sb_3__7_/prog_clk_2_N_out sb_3__7_/prog_clk_2_S_out
+ sb_3__7_/prog_clk_2_W_out sb_3__7_/prog_clk_3_E_out sb_3__7_/prog_clk_3_N_in sb_3__7_/prog_clk_3_N_out
+ sb_3__7_/prog_clk_3_S_out sb_3__7_/prog_clk_3_W_out sb_3__7_/right_bottom_grid_pin_34_
+ sb_3__7_/right_bottom_grid_pin_35_ sb_3__7_/right_bottom_grid_pin_36_ sb_3__7_/right_bottom_grid_pin_37_
+ sb_3__7_/right_bottom_grid_pin_38_ sb_3__7_/right_bottom_grid_pin_39_ sb_3__7_/right_bottom_grid_pin_40_
+ sb_3__7_/right_bottom_grid_pin_41_ sb_3__7_/top_left_grid_pin_42_ sb_3__7_/top_left_grid_pin_43_
+ sb_3__7_/top_left_grid_pin_44_ sb_3__7_/top_left_grid_pin_45_ sb_3__7_/top_left_grid_pin_46_
+ sb_3__7_/top_left_grid_pin_47_ sb_3__7_/top_left_grid_pin_48_ sb_3__7_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_0__4_ VGND VPWR sb_0__4_/bottom_left_grid_pin_1_ sb_0__4_/ccff_head sb_0__4_/ccff_tail
+ sb_0__4_/chanx_right_in[0] sb_0__4_/chanx_right_in[10] sb_0__4_/chanx_right_in[11]
+ sb_0__4_/chanx_right_in[12] sb_0__4_/chanx_right_in[13] sb_0__4_/chanx_right_in[14]
+ sb_0__4_/chanx_right_in[15] sb_0__4_/chanx_right_in[16] sb_0__4_/chanx_right_in[17]
+ sb_0__4_/chanx_right_in[18] sb_0__4_/chanx_right_in[19] sb_0__4_/chanx_right_in[1]
+ sb_0__4_/chanx_right_in[2] sb_0__4_/chanx_right_in[3] sb_0__4_/chanx_right_in[4]
+ sb_0__4_/chanx_right_in[5] sb_0__4_/chanx_right_in[6] sb_0__4_/chanx_right_in[7]
+ sb_0__4_/chanx_right_in[8] sb_0__4_/chanx_right_in[9] cbx_1__4_/chanx_left_in[0]
+ cbx_1__4_/chanx_left_in[10] cbx_1__4_/chanx_left_in[11] cbx_1__4_/chanx_left_in[12]
+ cbx_1__4_/chanx_left_in[13] cbx_1__4_/chanx_left_in[14] cbx_1__4_/chanx_left_in[15]
+ cbx_1__4_/chanx_left_in[16] cbx_1__4_/chanx_left_in[17] cbx_1__4_/chanx_left_in[18]
+ cbx_1__4_/chanx_left_in[19] cbx_1__4_/chanx_left_in[1] cbx_1__4_/chanx_left_in[2]
+ cbx_1__4_/chanx_left_in[3] cbx_1__4_/chanx_left_in[4] cbx_1__4_/chanx_left_in[5]
+ cbx_1__4_/chanx_left_in[6] cbx_1__4_/chanx_left_in[7] cbx_1__4_/chanx_left_in[8]
+ cbx_1__4_/chanx_left_in[9] cby_0__4_/chany_top_out[0] cby_0__4_/chany_top_out[10]
+ cby_0__4_/chany_top_out[11] cby_0__4_/chany_top_out[12] cby_0__4_/chany_top_out[13]
+ cby_0__4_/chany_top_out[14] cby_0__4_/chany_top_out[15] cby_0__4_/chany_top_out[16]
+ cby_0__4_/chany_top_out[17] cby_0__4_/chany_top_out[18] cby_0__4_/chany_top_out[19]
+ cby_0__4_/chany_top_out[1] cby_0__4_/chany_top_out[2] cby_0__4_/chany_top_out[3]
+ cby_0__4_/chany_top_out[4] cby_0__4_/chany_top_out[5] cby_0__4_/chany_top_out[6]
+ cby_0__4_/chany_top_out[7] cby_0__4_/chany_top_out[8] cby_0__4_/chany_top_out[9]
+ cby_0__4_/chany_top_in[0] cby_0__4_/chany_top_in[10] cby_0__4_/chany_top_in[11]
+ cby_0__4_/chany_top_in[12] cby_0__4_/chany_top_in[13] cby_0__4_/chany_top_in[14]
+ cby_0__4_/chany_top_in[15] cby_0__4_/chany_top_in[16] cby_0__4_/chany_top_in[17]
+ cby_0__4_/chany_top_in[18] cby_0__4_/chany_top_in[19] cby_0__4_/chany_top_in[1]
+ cby_0__4_/chany_top_in[2] cby_0__4_/chany_top_in[3] cby_0__4_/chany_top_in[4] cby_0__4_/chany_top_in[5]
+ cby_0__4_/chany_top_in[6] cby_0__4_/chany_top_in[7] cby_0__4_/chany_top_in[8] cby_0__4_/chany_top_in[9]
+ sb_0__4_/chany_top_in[0] sb_0__4_/chany_top_in[10] sb_0__4_/chany_top_in[11] sb_0__4_/chany_top_in[12]
+ sb_0__4_/chany_top_in[13] sb_0__4_/chany_top_in[14] sb_0__4_/chany_top_in[15] sb_0__4_/chany_top_in[16]
+ sb_0__4_/chany_top_in[17] sb_0__4_/chany_top_in[18] sb_0__4_/chany_top_in[19] sb_0__4_/chany_top_in[1]
+ sb_0__4_/chany_top_in[2] sb_0__4_/chany_top_in[3] sb_0__4_/chany_top_in[4] sb_0__4_/chany_top_in[5]
+ sb_0__4_/chany_top_in[6] sb_0__4_/chany_top_in[7] sb_0__4_/chany_top_in[8] sb_0__4_/chany_top_in[9]
+ sb_0__4_/chany_top_out[0] sb_0__4_/chany_top_out[10] sb_0__4_/chany_top_out[11]
+ sb_0__4_/chany_top_out[12] sb_0__4_/chany_top_out[13] sb_0__4_/chany_top_out[14]
+ sb_0__4_/chany_top_out[15] sb_0__4_/chany_top_out[16] sb_0__4_/chany_top_out[17]
+ sb_0__4_/chany_top_out[18] sb_0__4_/chany_top_out[19] sb_0__4_/chany_top_out[1]
+ sb_0__4_/chany_top_out[2] sb_0__4_/chany_top_out[3] sb_0__4_/chany_top_out[4] sb_0__4_/chany_top_out[5]
+ sb_0__4_/chany_top_out[6] sb_0__4_/chany_top_out[7] sb_0__4_/chany_top_out[8] sb_0__4_/chany_top_out[9]
+ sb_0__4_/prog_clk_0_E_in sb_0__4_/right_bottom_grid_pin_34_ sb_0__4_/right_bottom_grid_pin_35_
+ sb_0__4_/right_bottom_grid_pin_36_ sb_0__4_/right_bottom_grid_pin_37_ sb_0__4_/right_bottom_grid_pin_38_
+ sb_0__4_/right_bottom_grid_pin_39_ sb_0__4_/right_bottom_grid_pin_40_ sb_0__4_/right_bottom_grid_pin_41_
+ sb_0__4_/top_left_grid_pin_1_ sb_0__1_
Xcby_6__3_ cby_6__3_/Test_en_W_in cby_6__3_/Test_en_E_out cby_6__3_/Test_en_N_out
+ cby_6__3_/Test_en_W_in cby_6__3_/Test_en_W_in cby_6__3_/Test_en_W_out VGND VPWR
+ cby_6__3_/ccff_head cby_6__3_/ccff_tail sb_6__2_/chany_top_out[0] sb_6__2_/chany_top_out[10]
+ sb_6__2_/chany_top_out[11] sb_6__2_/chany_top_out[12] sb_6__2_/chany_top_out[13]
+ sb_6__2_/chany_top_out[14] sb_6__2_/chany_top_out[15] sb_6__2_/chany_top_out[16]
+ sb_6__2_/chany_top_out[17] sb_6__2_/chany_top_out[18] sb_6__2_/chany_top_out[19]
+ sb_6__2_/chany_top_out[1] sb_6__2_/chany_top_out[2] sb_6__2_/chany_top_out[3] sb_6__2_/chany_top_out[4]
+ sb_6__2_/chany_top_out[5] sb_6__2_/chany_top_out[6] sb_6__2_/chany_top_out[7] sb_6__2_/chany_top_out[8]
+ sb_6__2_/chany_top_out[9] sb_6__2_/chany_top_in[0] sb_6__2_/chany_top_in[10] sb_6__2_/chany_top_in[11]
+ sb_6__2_/chany_top_in[12] sb_6__2_/chany_top_in[13] sb_6__2_/chany_top_in[14] sb_6__2_/chany_top_in[15]
+ sb_6__2_/chany_top_in[16] sb_6__2_/chany_top_in[17] sb_6__2_/chany_top_in[18] sb_6__2_/chany_top_in[19]
+ sb_6__2_/chany_top_in[1] sb_6__2_/chany_top_in[2] sb_6__2_/chany_top_in[3] sb_6__2_/chany_top_in[4]
+ sb_6__2_/chany_top_in[5] sb_6__2_/chany_top_in[6] sb_6__2_/chany_top_in[7] sb_6__2_/chany_top_in[8]
+ sb_6__2_/chany_top_in[9] cby_6__3_/chany_top_in[0] cby_6__3_/chany_top_in[10] cby_6__3_/chany_top_in[11]
+ cby_6__3_/chany_top_in[12] cby_6__3_/chany_top_in[13] cby_6__3_/chany_top_in[14]
+ cby_6__3_/chany_top_in[15] cby_6__3_/chany_top_in[16] cby_6__3_/chany_top_in[17]
+ cby_6__3_/chany_top_in[18] cby_6__3_/chany_top_in[19] cby_6__3_/chany_top_in[1]
+ cby_6__3_/chany_top_in[2] cby_6__3_/chany_top_in[3] cby_6__3_/chany_top_in[4] cby_6__3_/chany_top_in[5]
+ cby_6__3_/chany_top_in[6] cby_6__3_/chany_top_in[7] cby_6__3_/chany_top_in[8] cby_6__3_/chany_top_in[9]
+ cby_6__3_/chany_top_out[0] cby_6__3_/chany_top_out[10] cby_6__3_/chany_top_out[11]
+ cby_6__3_/chany_top_out[12] cby_6__3_/chany_top_out[13] cby_6__3_/chany_top_out[14]
+ cby_6__3_/chany_top_out[15] cby_6__3_/chany_top_out[16] cby_6__3_/chany_top_out[17]
+ cby_6__3_/chany_top_out[18] cby_6__3_/chany_top_out[19] cby_6__3_/chany_top_out[1]
+ cby_6__3_/chany_top_out[2] cby_6__3_/chany_top_out[3] cby_6__3_/chany_top_out[4]
+ cby_6__3_/chany_top_out[5] cby_6__3_/chany_top_out[6] cby_6__3_/chany_top_out[7]
+ cby_6__3_/chany_top_out[8] cby_6__3_/chany_top_out[9] cby_6__3_/clk_2_N_out cby_6__3_/clk_2_S_in
+ cby_6__3_/clk_2_S_out cby_6__3_/clk_3_N_out sb_6__3_/clk_3_S_out sb_6__2_/clk_2_N_in
+ cby_6__3_/left_grid_pin_16_ cby_6__3_/left_grid_pin_17_ cby_6__3_/left_grid_pin_18_
+ cby_6__3_/left_grid_pin_19_ cby_6__3_/left_grid_pin_20_ cby_6__3_/left_grid_pin_21_
+ cby_6__3_/left_grid_pin_22_ cby_6__3_/left_grid_pin_23_ cby_6__3_/left_grid_pin_24_
+ cby_6__3_/left_grid_pin_25_ cby_6__3_/left_grid_pin_26_ cby_6__3_/left_grid_pin_27_
+ cby_6__3_/left_grid_pin_28_ cby_6__3_/left_grid_pin_29_ cby_6__3_/left_grid_pin_30_
+ cby_6__3_/left_grid_pin_31_ cby_6__3_/prog_clk_0_N_out sb_6__2_/prog_clk_0_N_in
+ cby_6__3_/prog_clk_0_W_in cby_6__3_/prog_clk_2_N_out cby_6__3_/prog_clk_2_S_in cby_6__3_/prog_clk_2_S_out
+ cby_6__3_/prog_clk_3_N_out sb_6__3_/prog_clk_3_S_out sb_6__2_/prog_clk_2_N_in cby_1__1_
Xgrid_clb_8__7_ cbx_8__6_/SC_OUT_TOP grid_clb_8__7_/SC_OUT_BOT cbx_8__7_/SC_IN_BOT
+ cby_7__7_/Test_en_E_out grid_clb_8__7_/Test_en_E_out cby_7__7_/Test_en_E_out grid_clb_8__7_/Test_en_W_out
+ VGND VPWR cbx_8__6_/REGIN_FEEDTHROUGH grid_clb_8__7_/bottom_width_0_height_0__pin_51_
+ cby_7__7_/ccff_tail cby_8__7_/ccff_head cbx_8__7_/clk_1_S_out cbx_8__7_/clk_1_S_out
+ cby_8__7_/prog_clk_0_W_in cbx_8__7_/prog_clk_1_S_out grid_clb_8__7_/prog_clk_0_N_out
+ cbx_8__7_/prog_clk_1_S_out cbx_8__6_/prog_clk_0_N_in grid_clb_8__7_/prog_clk_0_W_out
+ cby_8__7_/left_grid_pin_16_ cby_8__7_/left_grid_pin_17_ cby_8__7_/left_grid_pin_18_
+ cby_8__7_/left_grid_pin_19_ cby_8__7_/left_grid_pin_20_ cby_8__7_/left_grid_pin_21_
+ cby_8__7_/left_grid_pin_22_ cby_8__7_/left_grid_pin_23_ cby_8__7_/left_grid_pin_24_
+ cby_8__7_/left_grid_pin_25_ cby_8__7_/left_grid_pin_26_ cby_8__7_/left_grid_pin_27_
+ cby_8__7_/left_grid_pin_28_ cby_8__7_/left_grid_pin_29_ cby_8__7_/left_grid_pin_30_
+ cby_8__7_/left_grid_pin_31_ sb_8__6_/top_left_grid_pin_42_ sb_8__7_/bottom_left_grid_pin_42_
+ sb_8__6_/top_left_grid_pin_43_ sb_8__7_/bottom_left_grid_pin_43_ sb_8__6_/top_left_grid_pin_44_
+ sb_8__7_/bottom_left_grid_pin_44_ sb_8__6_/top_left_grid_pin_45_ sb_8__7_/bottom_left_grid_pin_45_
+ sb_8__6_/top_left_grid_pin_46_ sb_8__7_/bottom_left_grid_pin_46_ sb_8__6_/top_left_grid_pin_47_
+ sb_8__7_/bottom_left_grid_pin_47_ sb_8__6_/top_left_grid_pin_48_ sb_8__7_/bottom_left_grid_pin_48_
+ sb_8__6_/top_left_grid_pin_49_ sb_8__7_/bottom_left_grid_pin_49_ cbx_8__7_/bottom_grid_pin_0_
+ cbx_8__7_/bottom_grid_pin_10_ cbx_8__7_/bottom_grid_pin_11_ cbx_8__7_/bottom_grid_pin_12_
+ cbx_8__7_/bottom_grid_pin_13_ cbx_8__7_/bottom_grid_pin_14_ cbx_8__7_/bottom_grid_pin_15_
+ cbx_8__7_/bottom_grid_pin_1_ cbx_8__7_/bottom_grid_pin_2_ cbx_8__7_/REGOUT_FEEDTHROUGH
+ grid_clb_8__7_/top_width_0_height_0__pin_33_ sb_8__7_/left_bottom_grid_pin_34_ sb_7__7_/right_bottom_grid_pin_34_
+ sb_8__7_/left_bottom_grid_pin_35_ sb_7__7_/right_bottom_grid_pin_35_ sb_8__7_/left_bottom_grid_pin_36_
+ sb_7__7_/right_bottom_grid_pin_36_ sb_8__7_/left_bottom_grid_pin_37_ sb_7__7_/right_bottom_grid_pin_37_
+ sb_8__7_/left_bottom_grid_pin_38_ sb_7__7_/right_bottom_grid_pin_38_ sb_8__7_/left_bottom_grid_pin_39_
+ sb_7__7_/right_bottom_grid_pin_39_ cbx_8__7_/bottom_grid_pin_3_ sb_8__7_/left_bottom_grid_pin_40_
+ sb_7__7_/right_bottom_grid_pin_40_ sb_8__7_/left_bottom_grid_pin_41_ sb_7__7_/right_bottom_grid_pin_41_
+ cbx_8__7_/bottom_grid_pin_4_ cbx_8__7_/bottom_grid_pin_5_ cbx_8__7_/bottom_grid_pin_6_
+ cbx_8__7_/bottom_grid_pin_7_ cbx_8__7_/bottom_grid_pin_8_ cbx_8__7_/bottom_grid_pin_9_
+ grid_clb
Xcbx_6__4_ cbx_6__4_/REGIN_FEEDTHROUGH cbx_6__4_/REGOUT_FEEDTHROUGH cbx_6__4_/SC_IN_BOT
+ cbx_6__4_/SC_IN_TOP cbx_6__4_/SC_OUT_BOT cbx_6__4_/SC_OUT_TOP VGND VPWR cbx_6__4_/bottom_grid_pin_0_
+ cbx_6__4_/bottom_grid_pin_10_ cbx_6__4_/bottom_grid_pin_11_ cbx_6__4_/bottom_grid_pin_12_
+ cbx_6__4_/bottom_grid_pin_13_ cbx_6__4_/bottom_grid_pin_14_ cbx_6__4_/bottom_grid_pin_15_
+ cbx_6__4_/bottom_grid_pin_1_ cbx_6__4_/bottom_grid_pin_2_ cbx_6__4_/bottom_grid_pin_3_
+ cbx_6__4_/bottom_grid_pin_4_ cbx_6__4_/bottom_grid_pin_5_ cbx_6__4_/bottom_grid_pin_6_
+ cbx_6__4_/bottom_grid_pin_7_ cbx_6__4_/bottom_grid_pin_8_ cbx_6__4_/bottom_grid_pin_9_
+ sb_6__4_/ccff_tail sb_5__4_/ccff_head cbx_6__4_/chanx_left_in[0] cbx_6__4_/chanx_left_in[10]
+ cbx_6__4_/chanx_left_in[11] cbx_6__4_/chanx_left_in[12] cbx_6__4_/chanx_left_in[13]
+ cbx_6__4_/chanx_left_in[14] cbx_6__4_/chanx_left_in[15] cbx_6__4_/chanx_left_in[16]
+ cbx_6__4_/chanx_left_in[17] cbx_6__4_/chanx_left_in[18] cbx_6__4_/chanx_left_in[19]
+ cbx_6__4_/chanx_left_in[1] cbx_6__4_/chanx_left_in[2] cbx_6__4_/chanx_left_in[3]
+ cbx_6__4_/chanx_left_in[4] cbx_6__4_/chanx_left_in[5] cbx_6__4_/chanx_left_in[6]
+ cbx_6__4_/chanx_left_in[7] cbx_6__4_/chanx_left_in[8] cbx_6__4_/chanx_left_in[9]
+ sb_5__4_/chanx_right_in[0] sb_5__4_/chanx_right_in[10] sb_5__4_/chanx_right_in[11]
+ sb_5__4_/chanx_right_in[12] sb_5__4_/chanx_right_in[13] sb_5__4_/chanx_right_in[14]
+ sb_5__4_/chanx_right_in[15] sb_5__4_/chanx_right_in[16] sb_5__4_/chanx_right_in[17]
+ sb_5__4_/chanx_right_in[18] sb_5__4_/chanx_right_in[19] sb_5__4_/chanx_right_in[1]
+ sb_5__4_/chanx_right_in[2] sb_5__4_/chanx_right_in[3] sb_5__4_/chanx_right_in[4]
+ sb_5__4_/chanx_right_in[5] sb_5__4_/chanx_right_in[6] sb_5__4_/chanx_right_in[7]
+ sb_5__4_/chanx_right_in[8] sb_5__4_/chanx_right_in[9] sb_6__4_/chanx_left_out[0]
+ sb_6__4_/chanx_left_out[10] sb_6__4_/chanx_left_out[11] sb_6__4_/chanx_left_out[12]
+ sb_6__4_/chanx_left_out[13] sb_6__4_/chanx_left_out[14] sb_6__4_/chanx_left_out[15]
+ sb_6__4_/chanx_left_out[16] sb_6__4_/chanx_left_out[17] sb_6__4_/chanx_left_out[18]
+ sb_6__4_/chanx_left_out[19] sb_6__4_/chanx_left_out[1] sb_6__4_/chanx_left_out[2]
+ sb_6__4_/chanx_left_out[3] sb_6__4_/chanx_left_out[4] sb_6__4_/chanx_left_out[5]
+ sb_6__4_/chanx_left_out[6] sb_6__4_/chanx_left_out[7] sb_6__4_/chanx_left_out[8]
+ sb_6__4_/chanx_left_out[9] sb_6__4_/chanx_left_in[0] sb_6__4_/chanx_left_in[10]
+ sb_6__4_/chanx_left_in[11] sb_6__4_/chanx_left_in[12] sb_6__4_/chanx_left_in[13]
+ sb_6__4_/chanx_left_in[14] sb_6__4_/chanx_left_in[15] sb_6__4_/chanx_left_in[16]
+ sb_6__4_/chanx_left_in[17] sb_6__4_/chanx_left_in[18] sb_6__4_/chanx_left_in[19]
+ sb_6__4_/chanx_left_in[1] sb_6__4_/chanx_left_in[2] sb_6__4_/chanx_left_in[3] sb_6__4_/chanx_left_in[4]
+ sb_6__4_/chanx_left_in[5] sb_6__4_/chanx_left_in[6] sb_6__4_/chanx_left_in[7] sb_6__4_/chanx_left_in[8]
+ sb_6__4_/chanx_left_in[9] cbx_6__4_/clk_1_N_out cbx_6__4_/clk_1_S_out cbx_6__4_/clk_1_W_in
+ cbx_6__4_/clk_2_E_out cbx_6__4_/clk_2_W_in cbx_6__4_/clk_2_W_out sb_6__4_/clk_3_N_in
+ sb_5__4_/clk_3_E_out cbx_6__4_/clk_3_W_out cbx_6__4_/prog_clk_0_N_in cbx_6__4_/prog_clk_0_W_out
+ cbx_6__4_/prog_clk_1_N_out cbx_6__4_/prog_clk_1_S_out cbx_6__4_/prog_clk_1_W_in
+ cbx_6__4_/prog_clk_2_E_out cbx_6__4_/prog_clk_2_W_in cbx_6__4_/prog_clk_2_W_out
+ sb_6__4_/prog_clk_3_N_in sb_5__4_/prog_clk_3_E_out cbx_6__4_/prog_clk_3_W_out cbx_1__1_
Xgrid_clb_5__4_ cbx_5__4_/SC_OUT_BOT cbx_5__3_/SC_IN_TOP grid_clb_5__4_/SC_OUT_TOP
+ cby_4__4_/Test_en_E_out cby_5__4_/Test_en_W_in cby_4__4_/Test_en_E_out grid_clb_5__4_/Test_en_W_out
+ VGND VPWR cbx_5__3_/REGIN_FEEDTHROUGH grid_clb_5__4_/bottom_width_0_height_0__pin_51_
+ cby_4__4_/ccff_tail cby_5__4_/ccff_head cbx_5__3_/clk_1_N_out cbx_5__3_/clk_1_N_out
+ cby_5__4_/prog_clk_0_W_in cbx_5__3_/prog_clk_1_N_out grid_clb_5__4_/prog_clk_0_N_out
+ cbx_5__3_/prog_clk_1_N_out cbx_5__3_/prog_clk_0_N_in grid_clb_5__4_/prog_clk_0_W_out
+ cby_5__4_/left_grid_pin_16_ cby_5__4_/left_grid_pin_17_ cby_5__4_/left_grid_pin_18_
+ cby_5__4_/left_grid_pin_19_ cby_5__4_/left_grid_pin_20_ cby_5__4_/left_grid_pin_21_
+ cby_5__4_/left_grid_pin_22_ cby_5__4_/left_grid_pin_23_ cby_5__4_/left_grid_pin_24_
+ cby_5__4_/left_grid_pin_25_ cby_5__4_/left_grid_pin_26_ cby_5__4_/left_grid_pin_27_
+ cby_5__4_/left_grid_pin_28_ cby_5__4_/left_grid_pin_29_ cby_5__4_/left_grid_pin_30_
+ cby_5__4_/left_grid_pin_31_ sb_5__3_/top_left_grid_pin_42_ sb_5__4_/bottom_left_grid_pin_42_
+ sb_5__3_/top_left_grid_pin_43_ sb_5__4_/bottom_left_grid_pin_43_ sb_5__3_/top_left_grid_pin_44_
+ sb_5__4_/bottom_left_grid_pin_44_ sb_5__3_/top_left_grid_pin_45_ sb_5__4_/bottom_left_grid_pin_45_
+ sb_5__3_/top_left_grid_pin_46_ sb_5__4_/bottom_left_grid_pin_46_ sb_5__3_/top_left_grid_pin_47_
+ sb_5__4_/bottom_left_grid_pin_47_ sb_5__3_/top_left_grid_pin_48_ sb_5__4_/bottom_left_grid_pin_48_
+ sb_5__3_/top_left_grid_pin_49_ sb_5__4_/bottom_left_grid_pin_49_ cbx_5__4_/bottom_grid_pin_0_
+ cbx_5__4_/bottom_grid_pin_10_ cbx_5__4_/bottom_grid_pin_11_ cbx_5__4_/bottom_grid_pin_12_
+ cbx_5__4_/bottom_grid_pin_13_ cbx_5__4_/bottom_grid_pin_14_ cbx_5__4_/bottom_grid_pin_15_
+ cbx_5__4_/bottom_grid_pin_1_ cbx_5__4_/bottom_grid_pin_2_ cbx_5__4_/REGOUT_FEEDTHROUGH
+ grid_clb_5__4_/top_width_0_height_0__pin_33_ sb_5__4_/left_bottom_grid_pin_34_ sb_4__4_/right_bottom_grid_pin_34_
+ sb_5__4_/left_bottom_grid_pin_35_ sb_4__4_/right_bottom_grid_pin_35_ sb_5__4_/left_bottom_grid_pin_36_
+ sb_4__4_/right_bottom_grid_pin_36_ sb_5__4_/left_bottom_grid_pin_37_ sb_4__4_/right_bottom_grid_pin_37_
+ sb_5__4_/left_bottom_grid_pin_38_ sb_4__4_/right_bottom_grid_pin_38_ sb_5__4_/left_bottom_grid_pin_39_
+ sb_4__4_/right_bottom_grid_pin_39_ cbx_5__4_/bottom_grid_pin_3_ sb_5__4_/left_bottom_grid_pin_40_
+ sb_4__4_/right_bottom_grid_pin_40_ sb_5__4_/left_bottom_grid_pin_41_ sb_4__4_/right_bottom_grid_pin_41_
+ cbx_5__4_/bottom_grid_pin_4_ cbx_5__4_/bottom_grid_pin_5_ cbx_5__4_/bottom_grid_pin_6_
+ cbx_5__4_/bottom_grid_pin_7_ cbx_5__4_/bottom_grid_pin_8_ cbx_5__4_/bottom_grid_pin_9_
+ grid_clb
Xcbx_3__1_ cbx_3__1_/REGIN_FEEDTHROUGH cbx_3__1_/REGOUT_FEEDTHROUGH cbx_3__1_/SC_IN_BOT
+ cbx_3__1_/SC_IN_TOP cbx_3__1_/SC_OUT_BOT cbx_3__1_/SC_OUT_TOP VGND VPWR cbx_3__1_/bottom_grid_pin_0_
+ cbx_3__1_/bottom_grid_pin_10_ cbx_3__1_/bottom_grid_pin_11_ cbx_3__1_/bottom_grid_pin_12_
+ cbx_3__1_/bottom_grid_pin_13_ cbx_3__1_/bottom_grid_pin_14_ cbx_3__1_/bottom_grid_pin_15_
+ cbx_3__1_/bottom_grid_pin_1_ cbx_3__1_/bottom_grid_pin_2_ cbx_3__1_/bottom_grid_pin_3_
+ cbx_3__1_/bottom_grid_pin_4_ cbx_3__1_/bottom_grid_pin_5_ cbx_3__1_/bottom_grid_pin_6_
+ cbx_3__1_/bottom_grid_pin_7_ cbx_3__1_/bottom_grid_pin_8_ cbx_3__1_/bottom_grid_pin_9_
+ sb_3__1_/ccff_tail sb_2__1_/ccff_head cbx_3__1_/chanx_left_in[0] cbx_3__1_/chanx_left_in[10]
+ cbx_3__1_/chanx_left_in[11] cbx_3__1_/chanx_left_in[12] cbx_3__1_/chanx_left_in[13]
+ cbx_3__1_/chanx_left_in[14] cbx_3__1_/chanx_left_in[15] cbx_3__1_/chanx_left_in[16]
+ cbx_3__1_/chanx_left_in[17] cbx_3__1_/chanx_left_in[18] cbx_3__1_/chanx_left_in[19]
+ cbx_3__1_/chanx_left_in[1] cbx_3__1_/chanx_left_in[2] cbx_3__1_/chanx_left_in[3]
+ cbx_3__1_/chanx_left_in[4] cbx_3__1_/chanx_left_in[5] cbx_3__1_/chanx_left_in[6]
+ cbx_3__1_/chanx_left_in[7] cbx_3__1_/chanx_left_in[8] cbx_3__1_/chanx_left_in[9]
+ sb_2__1_/chanx_right_in[0] sb_2__1_/chanx_right_in[10] sb_2__1_/chanx_right_in[11]
+ sb_2__1_/chanx_right_in[12] sb_2__1_/chanx_right_in[13] sb_2__1_/chanx_right_in[14]
+ sb_2__1_/chanx_right_in[15] sb_2__1_/chanx_right_in[16] sb_2__1_/chanx_right_in[17]
+ sb_2__1_/chanx_right_in[18] sb_2__1_/chanx_right_in[19] sb_2__1_/chanx_right_in[1]
+ sb_2__1_/chanx_right_in[2] sb_2__1_/chanx_right_in[3] sb_2__1_/chanx_right_in[4]
+ sb_2__1_/chanx_right_in[5] sb_2__1_/chanx_right_in[6] sb_2__1_/chanx_right_in[7]
+ sb_2__1_/chanx_right_in[8] sb_2__1_/chanx_right_in[9] sb_3__1_/chanx_left_out[0]
+ sb_3__1_/chanx_left_out[10] sb_3__1_/chanx_left_out[11] sb_3__1_/chanx_left_out[12]
+ sb_3__1_/chanx_left_out[13] sb_3__1_/chanx_left_out[14] sb_3__1_/chanx_left_out[15]
+ sb_3__1_/chanx_left_out[16] sb_3__1_/chanx_left_out[17] sb_3__1_/chanx_left_out[18]
+ sb_3__1_/chanx_left_out[19] sb_3__1_/chanx_left_out[1] sb_3__1_/chanx_left_out[2]
+ sb_3__1_/chanx_left_out[3] sb_3__1_/chanx_left_out[4] sb_3__1_/chanx_left_out[5]
+ sb_3__1_/chanx_left_out[6] sb_3__1_/chanx_left_out[7] sb_3__1_/chanx_left_out[8]
+ sb_3__1_/chanx_left_out[9] sb_3__1_/chanx_left_in[0] sb_3__1_/chanx_left_in[10]
+ sb_3__1_/chanx_left_in[11] sb_3__1_/chanx_left_in[12] sb_3__1_/chanx_left_in[13]
+ sb_3__1_/chanx_left_in[14] sb_3__1_/chanx_left_in[15] sb_3__1_/chanx_left_in[16]
+ sb_3__1_/chanx_left_in[17] sb_3__1_/chanx_left_in[18] sb_3__1_/chanx_left_in[19]
+ sb_3__1_/chanx_left_in[1] sb_3__1_/chanx_left_in[2] sb_3__1_/chanx_left_in[3] sb_3__1_/chanx_left_in[4]
+ sb_3__1_/chanx_left_in[5] sb_3__1_/chanx_left_in[6] sb_3__1_/chanx_left_in[7] sb_3__1_/chanx_left_in[8]
+ sb_3__1_/chanx_left_in[9] cbx_3__1_/clk_1_N_out cbx_3__1_/clk_1_S_out sb_3__1_/clk_1_W_out
+ cbx_3__1_/clk_2_E_out cbx_3__1_/clk_2_W_in cbx_3__1_/clk_2_W_out cbx_3__1_/clk_3_E_out
+ cbx_3__1_/clk_3_W_in cbx_3__1_/clk_3_W_out cbx_3__1_/prog_clk_0_N_in cbx_3__1_/prog_clk_0_W_out
+ cbx_3__1_/prog_clk_1_N_out cbx_3__1_/prog_clk_1_S_out sb_3__1_/prog_clk_1_W_out
+ cbx_3__1_/prog_clk_2_E_out cbx_3__1_/prog_clk_2_W_in cbx_3__1_/prog_clk_2_W_out
+ cbx_3__1_/prog_clk_3_E_out cbx_3__1_/prog_clk_3_W_in cbx_3__1_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_3__6_ sb_3__6_/Test_en_N_out sb_3__6_/Test_en_S_in VGND VPWR sb_3__6_/bottom_left_grid_pin_42_
+ sb_3__6_/bottom_left_grid_pin_43_ sb_3__6_/bottom_left_grid_pin_44_ sb_3__6_/bottom_left_grid_pin_45_
+ sb_3__6_/bottom_left_grid_pin_46_ sb_3__6_/bottom_left_grid_pin_47_ sb_3__6_/bottom_left_grid_pin_48_
+ sb_3__6_/bottom_left_grid_pin_49_ sb_3__6_/ccff_head sb_3__6_/ccff_tail sb_3__6_/chanx_left_in[0]
+ sb_3__6_/chanx_left_in[10] sb_3__6_/chanx_left_in[11] sb_3__6_/chanx_left_in[12]
+ sb_3__6_/chanx_left_in[13] sb_3__6_/chanx_left_in[14] sb_3__6_/chanx_left_in[15]
+ sb_3__6_/chanx_left_in[16] sb_3__6_/chanx_left_in[17] sb_3__6_/chanx_left_in[18]
+ sb_3__6_/chanx_left_in[19] sb_3__6_/chanx_left_in[1] sb_3__6_/chanx_left_in[2] sb_3__6_/chanx_left_in[3]
+ sb_3__6_/chanx_left_in[4] sb_3__6_/chanx_left_in[5] sb_3__6_/chanx_left_in[6] sb_3__6_/chanx_left_in[7]
+ sb_3__6_/chanx_left_in[8] sb_3__6_/chanx_left_in[9] sb_3__6_/chanx_left_out[0] sb_3__6_/chanx_left_out[10]
+ sb_3__6_/chanx_left_out[11] sb_3__6_/chanx_left_out[12] sb_3__6_/chanx_left_out[13]
+ sb_3__6_/chanx_left_out[14] sb_3__6_/chanx_left_out[15] sb_3__6_/chanx_left_out[16]
+ sb_3__6_/chanx_left_out[17] sb_3__6_/chanx_left_out[18] sb_3__6_/chanx_left_out[19]
+ sb_3__6_/chanx_left_out[1] sb_3__6_/chanx_left_out[2] sb_3__6_/chanx_left_out[3]
+ sb_3__6_/chanx_left_out[4] sb_3__6_/chanx_left_out[5] sb_3__6_/chanx_left_out[6]
+ sb_3__6_/chanx_left_out[7] sb_3__6_/chanx_left_out[8] sb_3__6_/chanx_left_out[9]
+ sb_3__6_/chanx_right_in[0] sb_3__6_/chanx_right_in[10] sb_3__6_/chanx_right_in[11]
+ sb_3__6_/chanx_right_in[12] sb_3__6_/chanx_right_in[13] sb_3__6_/chanx_right_in[14]
+ sb_3__6_/chanx_right_in[15] sb_3__6_/chanx_right_in[16] sb_3__6_/chanx_right_in[17]
+ sb_3__6_/chanx_right_in[18] sb_3__6_/chanx_right_in[19] sb_3__6_/chanx_right_in[1]
+ sb_3__6_/chanx_right_in[2] sb_3__6_/chanx_right_in[3] sb_3__6_/chanx_right_in[4]
+ sb_3__6_/chanx_right_in[5] sb_3__6_/chanx_right_in[6] sb_3__6_/chanx_right_in[7]
+ sb_3__6_/chanx_right_in[8] sb_3__6_/chanx_right_in[9] cbx_4__6_/chanx_left_in[0]
+ cbx_4__6_/chanx_left_in[10] cbx_4__6_/chanx_left_in[11] cbx_4__6_/chanx_left_in[12]
+ cbx_4__6_/chanx_left_in[13] cbx_4__6_/chanx_left_in[14] cbx_4__6_/chanx_left_in[15]
+ cbx_4__6_/chanx_left_in[16] cbx_4__6_/chanx_left_in[17] cbx_4__6_/chanx_left_in[18]
+ cbx_4__6_/chanx_left_in[19] cbx_4__6_/chanx_left_in[1] cbx_4__6_/chanx_left_in[2]
+ cbx_4__6_/chanx_left_in[3] cbx_4__6_/chanx_left_in[4] cbx_4__6_/chanx_left_in[5]
+ cbx_4__6_/chanx_left_in[6] cbx_4__6_/chanx_left_in[7] cbx_4__6_/chanx_left_in[8]
+ cbx_4__6_/chanx_left_in[9] cby_3__6_/chany_top_out[0] cby_3__6_/chany_top_out[10]
+ cby_3__6_/chany_top_out[11] cby_3__6_/chany_top_out[12] cby_3__6_/chany_top_out[13]
+ cby_3__6_/chany_top_out[14] cby_3__6_/chany_top_out[15] cby_3__6_/chany_top_out[16]
+ cby_3__6_/chany_top_out[17] cby_3__6_/chany_top_out[18] cby_3__6_/chany_top_out[19]
+ cby_3__6_/chany_top_out[1] cby_3__6_/chany_top_out[2] cby_3__6_/chany_top_out[3]
+ cby_3__6_/chany_top_out[4] cby_3__6_/chany_top_out[5] cby_3__6_/chany_top_out[6]
+ cby_3__6_/chany_top_out[7] cby_3__6_/chany_top_out[8] cby_3__6_/chany_top_out[9]
+ cby_3__6_/chany_top_in[0] cby_3__6_/chany_top_in[10] cby_3__6_/chany_top_in[11]
+ cby_3__6_/chany_top_in[12] cby_3__6_/chany_top_in[13] cby_3__6_/chany_top_in[14]
+ cby_3__6_/chany_top_in[15] cby_3__6_/chany_top_in[16] cby_3__6_/chany_top_in[17]
+ cby_3__6_/chany_top_in[18] cby_3__6_/chany_top_in[19] cby_3__6_/chany_top_in[1]
+ cby_3__6_/chany_top_in[2] cby_3__6_/chany_top_in[3] cby_3__6_/chany_top_in[4] cby_3__6_/chany_top_in[5]
+ cby_3__6_/chany_top_in[6] cby_3__6_/chany_top_in[7] cby_3__6_/chany_top_in[8] cby_3__6_/chany_top_in[9]
+ sb_3__6_/chany_top_in[0] sb_3__6_/chany_top_in[10] sb_3__6_/chany_top_in[11] sb_3__6_/chany_top_in[12]
+ sb_3__6_/chany_top_in[13] sb_3__6_/chany_top_in[14] sb_3__6_/chany_top_in[15] sb_3__6_/chany_top_in[16]
+ sb_3__6_/chany_top_in[17] sb_3__6_/chany_top_in[18] sb_3__6_/chany_top_in[19] sb_3__6_/chany_top_in[1]
+ sb_3__6_/chany_top_in[2] sb_3__6_/chany_top_in[3] sb_3__6_/chany_top_in[4] sb_3__6_/chany_top_in[5]
+ sb_3__6_/chany_top_in[6] sb_3__6_/chany_top_in[7] sb_3__6_/chany_top_in[8] sb_3__6_/chany_top_in[9]
+ sb_3__6_/chany_top_out[0] sb_3__6_/chany_top_out[10] sb_3__6_/chany_top_out[11]
+ sb_3__6_/chany_top_out[12] sb_3__6_/chany_top_out[13] sb_3__6_/chany_top_out[14]
+ sb_3__6_/chany_top_out[15] sb_3__6_/chany_top_out[16] sb_3__6_/chany_top_out[17]
+ sb_3__6_/chany_top_out[18] sb_3__6_/chany_top_out[19] sb_3__6_/chany_top_out[1]
+ sb_3__6_/chany_top_out[2] sb_3__6_/chany_top_out[3] sb_3__6_/chany_top_out[4] sb_3__6_/chany_top_out[5]
+ sb_3__6_/chany_top_out[6] sb_3__6_/chany_top_out[7] sb_3__6_/chany_top_out[8] sb_3__6_/chany_top_out[9]
+ sb_3__6_/clk_1_E_out sb_3__6_/clk_1_N_in sb_3__6_/clk_1_W_out sb_3__6_/clk_2_E_out
+ sb_3__6_/clk_2_N_in sb_3__6_/clk_2_N_out sb_3__6_/clk_2_S_out sb_3__6_/clk_2_W_out
+ sb_3__6_/clk_3_E_out sb_3__6_/clk_3_N_in sb_3__6_/clk_3_N_out sb_3__6_/clk_3_S_out
+ sb_3__6_/clk_3_W_out sb_3__6_/left_bottom_grid_pin_34_ sb_3__6_/left_bottom_grid_pin_35_
+ sb_3__6_/left_bottom_grid_pin_36_ sb_3__6_/left_bottom_grid_pin_37_ sb_3__6_/left_bottom_grid_pin_38_
+ sb_3__6_/left_bottom_grid_pin_39_ sb_3__6_/left_bottom_grid_pin_40_ sb_3__6_/left_bottom_grid_pin_41_
+ sb_3__6_/prog_clk_0_N_in sb_3__6_/prog_clk_1_E_out sb_3__6_/prog_clk_1_N_in sb_3__6_/prog_clk_1_W_out
+ sb_3__6_/prog_clk_2_E_out sb_3__6_/prog_clk_2_N_in sb_3__6_/prog_clk_2_N_out sb_3__6_/prog_clk_2_S_out
+ sb_3__6_/prog_clk_2_W_out sb_3__6_/prog_clk_3_E_out sb_3__6_/prog_clk_3_N_in sb_3__6_/prog_clk_3_N_out
+ sb_3__6_/prog_clk_3_S_out sb_3__6_/prog_clk_3_W_out sb_3__6_/right_bottom_grid_pin_34_
+ sb_3__6_/right_bottom_grid_pin_35_ sb_3__6_/right_bottom_grid_pin_36_ sb_3__6_/right_bottom_grid_pin_37_
+ sb_3__6_/right_bottom_grid_pin_38_ sb_3__6_/right_bottom_grid_pin_39_ sb_3__6_/right_bottom_grid_pin_40_
+ sb_3__6_/right_bottom_grid_pin_41_ sb_3__6_/top_left_grid_pin_42_ sb_3__6_/top_left_grid_pin_43_
+ sb_3__6_/top_left_grid_pin_44_ sb_3__6_/top_left_grid_pin_45_ sb_3__6_/top_left_grid_pin_46_
+ sb_3__6_/top_left_grid_pin_47_ sb_3__6_/top_left_grid_pin_48_ sb_3__6_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_2__1_ cbx_2__0_/SC_OUT_TOP grid_clb_2__1_/SC_OUT_BOT cbx_2__1_/SC_IN_BOT
+ cby_2__1_/Test_en_W_out grid_clb_2__1_/Test_en_E_out cby_2__1_/Test_en_W_out cby_1__1_/Test_en_W_in
+ VGND VPWR grid_clb_2__1_/bottom_width_0_height_0__pin_50_ grid_clb_2__1_/bottom_width_0_height_0__pin_51_
+ cby_1__1_/ccff_tail cby_2__1_/ccff_head cbx_2__1_/clk_1_S_out cbx_2__1_/clk_1_S_out
+ cby_2__1_/prog_clk_0_W_in cbx_2__1_/prog_clk_1_S_out grid_clb_2__1_/prog_clk_0_N_out
+ cbx_2__1_/prog_clk_1_S_out cbx_2__0_/prog_clk_0_N_in grid_clb_2__1_/prog_clk_0_W_out
+ cby_2__1_/left_grid_pin_16_ cby_2__1_/left_grid_pin_17_ cby_2__1_/left_grid_pin_18_
+ cby_2__1_/left_grid_pin_19_ cby_2__1_/left_grid_pin_20_ cby_2__1_/left_grid_pin_21_
+ cby_2__1_/left_grid_pin_22_ cby_2__1_/left_grid_pin_23_ cby_2__1_/left_grid_pin_24_
+ cby_2__1_/left_grid_pin_25_ cby_2__1_/left_grid_pin_26_ cby_2__1_/left_grid_pin_27_
+ cby_2__1_/left_grid_pin_28_ cby_2__1_/left_grid_pin_29_ cby_2__1_/left_grid_pin_30_
+ cby_2__1_/left_grid_pin_31_ sb_2__0_/top_left_grid_pin_42_ sb_2__1_/bottom_left_grid_pin_42_
+ sb_2__0_/top_left_grid_pin_43_ sb_2__1_/bottom_left_grid_pin_43_ sb_2__0_/top_left_grid_pin_44_
+ sb_2__1_/bottom_left_grid_pin_44_ sb_2__0_/top_left_grid_pin_45_ sb_2__1_/bottom_left_grid_pin_45_
+ sb_2__0_/top_left_grid_pin_46_ sb_2__1_/bottom_left_grid_pin_46_ sb_2__0_/top_left_grid_pin_47_
+ sb_2__1_/bottom_left_grid_pin_47_ sb_2__0_/top_left_grid_pin_48_ sb_2__1_/bottom_left_grid_pin_48_
+ sb_2__0_/top_left_grid_pin_49_ sb_2__1_/bottom_left_grid_pin_49_ cbx_2__1_/bottom_grid_pin_0_
+ cbx_2__1_/bottom_grid_pin_10_ cbx_2__1_/bottom_grid_pin_11_ cbx_2__1_/bottom_grid_pin_12_
+ cbx_2__1_/bottom_grid_pin_13_ cbx_2__1_/bottom_grid_pin_14_ cbx_2__1_/bottom_grid_pin_15_
+ cbx_2__1_/bottom_grid_pin_1_ cbx_2__1_/bottom_grid_pin_2_ cbx_2__1_/REGOUT_FEEDTHROUGH
+ grid_clb_2__1_/top_width_0_height_0__pin_33_ sb_2__1_/left_bottom_grid_pin_34_ sb_1__1_/right_bottom_grid_pin_34_
+ sb_2__1_/left_bottom_grid_pin_35_ sb_1__1_/right_bottom_grid_pin_35_ sb_2__1_/left_bottom_grid_pin_36_
+ sb_1__1_/right_bottom_grid_pin_36_ sb_2__1_/left_bottom_grid_pin_37_ sb_1__1_/right_bottom_grid_pin_37_
+ sb_2__1_/left_bottom_grid_pin_38_ sb_1__1_/right_bottom_grid_pin_38_ sb_2__1_/left_bottom_grid_pin_39_
+ sb_1__1_/right_bottom_grid_pin_39_ cbx_2__1_/bottom_grid_pin_3_ sb_2__1_/left_bottom_grid_pin_40_
+ sb_1__1_/right_bottom_grid_pin_40_ sb_2__1_/left_bottom_grid_pin_41_ sb_1__1_/right_bottom_grid_pin_41_
+ cbx_2__1_/bottom_grid_pin_4_ cbx_2__1_/bottom_grid_pin_5_ cbx_2__1_/bottom_grid_pin_6_
+ cbx_2__1_/bottom_grid_pin_7_ cbx_2__1_/bottom_grid_pin_8_ cbx_2__1_/bottom_grid_pin_9_
+ grid_clb
Xsb_0__3_ VGND VPWR sb_0__3_/bottom_left_grid_pin_1_ sb_0__3_/ccff_head sb_0__3_/ccff_tail
+ sb_0__3_/chanx_right_in[0] sb_0__3_/chanx_right_in[10] sb_0__3_/chanx_right_in[11]
+ sb_0__3_/chanx_right_in[12] sb_0__3_/chanx_right_in[13] sb_0__3_/chanx_right_in[14]
+ sb_0__3_/chanx_right_in[15] sb_0__3_/chanx_right_in[16] sb_0__3_/chanx_right_in[17]
+ sb_0__3_/chanx_right_in[18] sb_0__3_/chanx_right_in[19] sb_0__3_/chanx_right_in[1]
+ sb_0__3_/chanx_right_in[2] sb_0__3_/chanx_right_in[3] sb_0__3_/chanx_right_in[4]
+ sb_0__3_/chanx_right_in[5] sb_0__3_/chanx_right_in[6] sb_0__3_/chanx_right_in[7]
+ sb_0__3_/chanx_right_in[8] sb_0__3_/chanx_right_in[9] cbx_1__3_/chanx_left_in[0]
+ cbx_1__3_/chanx_left_in[10] cbx_1__3_/chanx_left_in[11] cbx_1__3_/chanx_left_in[12]
+ cbx_1__3_/chanx_left_in[13] cbx_1__3_/chanx_left_in[14] cbx_1__3_/chanx_left_in[15]
+ cbx_1__3_/chanx_left_in[16] cbx_1__3_/chanx_left_in[17] cbx_1__3_/chanx_left_in[18]
+ cbx_1__3_/chanx_left_in[19] cbx_1__3_/chanx_left_in[1] cbx_1__3_/chanx_left_in[2]
+ cbx_1__3_/chanx_left_in[3] cbx_1__3_/chanx_left_in[4] cbx_1__3_/chanx_left_in[5]
+ cbx_1__3_/chanx_left_in[6] cbx_1__3_/chanx_left_in[7] cbx_1__3_/chanx_left_in[8]
+ cbx_1__3_/chanx_left_in[9] cby_0__3_/chany_top_out[0] cby_0__3_/chany_top_out[10]
+ cby_0__3_/chany_top_out[11] cby_0__3_/chany_top_out[12] cby_0__3_/chany_top_out[13]
+ cby_0__3_/chany_top_out[14] cby_0__3_/chany_top_out[15] cby_0__3_/chany_top_out[16]
+ cby_0__3_/chany_top_out[17] cby_0__3_/chany_top_out[18] cby_0__3_/chany_top_out[19]
+ cby_0__3_/chany_top_out[1] cby_0__3_/chany_top_out[2] cby_0__3_/chany_top_out[3]
+ cby_0__3_/chany_top_out[4] cby_0__3_/chany_top_out[5] cby_0__3_/chany_top_out[6]
+ cby_0__3_/chany_top_out[7] cby_0__3_/chany_top_out[8] cby_0__3_/chany_top_out[9]
+ cby_0__3_/chany_top_in[0] cby_0__3_/chany_top_in[10] cby_0__3_/chany_top_in[11]
+ cby_0__3_/chany_top_in[12] cby_0__3_/chany_top_in[13] cby_0__3_/chany_top_in[14]
+ cby_0__3_/chany_top_in[15] cby_0__3_/chany_top_in[16] cby_0__3_/chany_top_in[17]
+ cby_0__3_/chany_top_in[18] cby_0__3_/chany_top_in[19] cby_0__3_/chany_top_in[1]
+ cby_0__3_/chany_top_in[2] cby_0__3_/chany_top_in[3] cby_0__3_/chany_top_in[4] cby_0__3_/chany_top_in[5]
+ cby_0__3_/chany_top_in[6] cby_0__3_/chany_top_in[7] cby_0__3_/chany_top_in[8] cby_0__3_/chany_top_in[9]
+ sb_0__3_/chany_top_in[0] sb_0__3_/chany_top_in[10] sb_0__3_/chany_top_in[11] sb_0__3_/chany_top_in[12]
+ sb_0__3_/chany_top_in[13] sb_0__3_/chany_top_in[14] sb_0__3_/chany_top_in[15] sb_0__3_/chany_top_in[16]
+ sb_0__3_/chany_top_in[17] sb_0__3_/chany_top_in[18] sb_0__3_/chany_top_in[19] sb_0__3_/chany_top_in[1]
+ sb_0__3_/chany_top_in[2] sb_0__3_/chany_top_in[3] sb_0__3_/chany_top_in[4] sb_0__3_/chany_top_in[5]
+ sb_0__3_/chany_top_in[6] sb_0__3_/chany_top_in[7] sb_0__3_/chany_top_in[8] sb_0__3_/chany_top_in[9]
+ sb_0__3_/chany_top_out[0] sb_0__3_/chany_top_out[10] sb_0__3_/chany_top_out[11]
+ sb_0__3_/chany_top_out[12] sb_0__3_/chany_top_out[13] sb_0__3_/chany_top_out[14]
+ sb_0__3_/chany_top_out[15] sb_0__3_/chany_top_out[16] sb_0__3_/chany_top_out[17]
+ sb_0__3_/chany_top_out[18] sb_0__3_/chany_top_out[19] sb_0__3_/chany_top_out[1]
+ sb_0__3_/chany_top_out[2] sb_0__3_/chany_top_out[3] sb_0__3_/chany_top_out[4] sb_0__3_/chany_top_out[5]
+ sb_0__3_/chany_top_out[6] sb_0__3_/chany_top_out[7] sb_0__3_/chany_top_out[8] sb_0__3_/chany_top_out[9]
+ sb_0__3_/prog_clk_0_E_in sb_0__3_/right_bottom_grid_pin_34_ sb_0__3_/right_bottom_grid_pin_35_
+ sb_0__3_/right_bottom_grid_pin_36_ sb_0__3_/right_bottom_grid_pin_37_ sb_0__3_/right_bottom_grid_pin_38_
+ sb_0__3_/right_bottom_grid_pin_39_ sb_0__3_/right_bottom_grid_pin_40_ sb_0__3_/right_bottom_grid_pin_41_
+ sb_0__3_/top_left_grid_pin_1_ sb_0__1_
Xcby_6__2_ cby_6__2_/Test_en_W_in cby_6__2_/Test_en_E_out cby_6__2_/Test_en_N_out
+ cby_6__2_/Test_en_W_in cby_6__2_/Test_en_W_in cby_6__2_/Test_en_W_out VGND VPWR
+ cby_6__2_/ccff_head cby_6__2_/ccff_tail sb_6__1_/chany_top_out[0] sb_6__1_/chany_top_out[10]
+ sb_6__1_/chany_top_out[11] sb_6__1_/chany_top_out[12] sb_6__1_/chany_top_out[13]
+ sb_6__1_/chany_top_out[14] sb_6__1_/chany_top_out[15] sb_6__1_/chany_top_out[16]
+ sb_6__1_/chany_top_out[17] sb_6__1_/chany_top_out[18] sb_6__1_/chany_top_out[19]
+ sb_6__1_/chany_top_out[1] sb_6__1_/chany_top_out[2] sb_6__1_/chany_top_out[3] sb_6__1_/chany_top_out[4]
+ sb_6__1_/chany_top_out[5] sb_6__1_/chany_top_out[6] sb_6__1_/chany_top_out[7] sb_6__1_/chany_top_out[8]
+ sb_6__1_/chany_top_out[9] sb_6__1_/chany_top_in[0] sb_6__1_/chany_top_in[10] sb_6__1_/chany_top_in[11]
+ sb_6__1_/chany_top_in[12] sb_6__1_/chany_top_in[13] sb_6__1_/chany_top_in[14] sb_6__1_/chany_top_in[15]
+ sb_6__1_/chany_top_in[16] sb_6__1_/chany_top_in[17] sb_6__1_/chany_top_in[18] sb_6__1_/chany_top_in[19]
+ sb_6__1_/chany_top_in[1] sb_6__1_/chany_top_in[2] sb_6__1_/chany_top_in[3] sb_6__1_/chany_top_in[4]
+ sb_6__1_/chany_top_in[5] sb_6__1_/chany_top_in[6] sb_6__1_/chany_top_in[7] sb_6__1_/chany_top_in[8]
+ sb_6__1_/chany_top_in[9] cby_6__2_/chany_top_in[0] cby_6__2_/chany_top_in[10] cby_6__2_/chany_top_in[11]
+ cby_6__2_/chany_top_in[12] cby_6__2_/chany_top_in[13] cby_6__2_/chany_top_in[14]
+ cby_6__2_/chany_top_in[15] cby_6__2_/chany_top_in[16] cby_6__2_/chany_top_in[17]
+ cby_6__2_/chany_top_in[18] cby_6__2_/chany_top_in[19] cby_6__2_/chany_top_in[1]
+ cby_6__2_/chany_top_in[2] cby_6__2_/chany_top_in[3] cby_6__2_/chany_top_in[4] cby_6__2_/chany_top_in[5]
+ cby_6__2_/chany_top_in[6] cby_6__2_/chany_top_in[7] cby_6__2_/chany_top_in[8] cby_6__2_/chany_top_in[9]
+ cby_6__2_/chany_top_out[0] cby_6__2_/chany_top_out[10] cby_6__2_/chany_top_out[11]
+ cby_6__2_/chany_top_out[12] cby_6__2_/chany_top_out[13] cby_6__2_/chany_top_out[14]
+ cby_6__2_/chany_top_out[15] cby_6__2_/chany_top_out[16] cby_6__2_/chany_top_out[17]
+ cby_6__2_/chany_top_out[18] cby_6__2_/chany_top_out[19] cby_6__2_/chany_top_out[1]
+ cby_6__2_/chany_top_out[2] cby_6__2_/chany_top_out[3] cby_6__2_/chany_top_out[4]
+ cby_6__2_/chany_top_out[5] cby_6__2_/chany_top_out[6] cby_6__2_/chany_top_out[7]
+ cby_6__2_/chany_top_out[8] cby_6__2_/chany_top_out[9] cby_6__2_/clk_2_N_out cby_6__2_/clk_2_S_in
+ cby_6__2_/clk_2_S_out cby_6__2_/clk_3_N_out cby_6__2_/clk_3_S_in cby_6__2_/clk_3_S_out
+ cby_6__2_/left_grid_pin_16_ cby_6__2_/left_grid_pin_17_ cby_6__2_/left_grid_pin_18_
+ cby_6__2_/left_grid_pin_19_ cby_6__2_/left_grid_pin_20_ cby_6__2_/left_grid_pin_21_
+ cby_6__2_/left_grid_pin_22_ cby_6__2_/left_grid_pin_23_ cby_6__2_/left_grid_pin_24_
+ cby_6__2_/left_grid_pin_25_ cby_6__2_/left_grid_pin_26_ cby_6__2_/left_grid_pin_27_
+ cby_6__2_/left_grid_pin_28_ cby_6__2_/left_grid_pin_29_ cby_6__2_/left_grid_pin_30_
+ cby_6__2_/left_grid_pin_31_ cby_6__2_/prog_clk_0_N_out sb_6__1_/prog_clk_0_N_in
+ cby_6__2_/prog_clk_0_W_in cby_6__2_/prog_clk_2_N_out cby_6__2_/prog_clk_2_S_in cby_6__2_/prog_clk_2_S_out
+ cby_6__2_/prog_clk_3_N_out cby_6__2_/prog_clk_3_S_in cby_6__2_/prog_clk_3_S_out
+ cby_1__1_
Xcbx_6__3_ cbx_6__3_/REGIN_FEEDTHROUGH cbx_6__3_/REGOUT_FEEDTHROUGH cbx_6__3_/SC_IN_BOT
+ cbx_6__3_/SC_IN_TOP cbx_6__3_/SC_OUT_BOT cbx_6__3_/SC_OUT_TOP VGND VPWR cbx_6__3_/bottom_grid_pin_0_
+ cbx_6__3_/bottom_grid_pin_10_ cbx_6__3_/bottom_grid_pin_11_ cbx_6__3_/bottom_grid_pin_12_
+ cbx_6__3_/bottom_grid_pin_13_ cbx_6__3_/bottom_grid_pin_14_ cbx_6__3_/bottom_grid_pin_15_
+ cbx_6__3_/bottom_grid_pin_1_ cbx_6__3_/bottom_grid_pin_2_ cbx_6__3_/bottom_grid_pin_3_
+ cbx_6__3_/bottom_grid_pin_4_ cbx_6__3_/bottom_grid_pin_5_ cbx_6__3_/bottom_grid_pin_6_
+ cbx_6__3_/bottom_grid_pin_7_ cbx_6__3_/bottom_grid_pin_8_ cbx_6__3_/bottom_grid_pin_9_
+ sb_6__3_/ccff_tail sb_5__3_/ccff_head cbx_6__3_/chanx_left_in[0] cbx_6__3_/chanx_left_in[10]
+ cbx_6__3_/chanx_left_in[11] cbx_6__3_/chanx_left_in[12] cbx_6__3_/chanx_left_in[13]
+ cbx_6__3_/chanx_left_in[14] cbx_6__3_/chanx_left_in[15] cbx_6__3_/chanx_left_in[16]
+ cbx_6__3_/chanx_left_in[17] cbx_6__3_/chanx_left_in[18] cbx_6__3_/chanx_left_in[19]
+ cbx_6__3_/chanx_left_in[1] cbx_6__3_/chanx_left_in[2] cbx_6__3_/chanx_left_in[3]
+ cbx_6__3_/chanx_left_in[4] cbx_6__3_/chanx_left_in[5] cbx_6__3_/chanx_left_in[6]
+ cbx_6__3_/chanx_left_in[7] cbx_6__3_/chanx_left_in[8] cbx_6__3_/chanx_left_in[9]
+ sb_5__3_/chanx_right_in[0] sb_5__3_/chanx_right_in[10] sb_5__3_/chanx_right_in[11]
+ sb_5__3_/chanx_right_in[12] sb_5__3_/chanx_right_in[13] sb_5__3_/chanx_right_in[14]
+ sb_5__3_/chanx_right_in[15] sb_5__3_/chanx_right_in[16] sb_5__3_/chanx_right_in[17]
+ sb_5__3_/chanx_right_in[18] sb_5__3_/chanx_right_in[19] sb_5__3_/chanx_right_in[1]
+ sb_5__3_/chanx_right_in[2] sb_5__3_/chanx_right_in[3] sb_5__3_/chanx_right_in[4]
+ sb_5__3_/chanx_right_in[5] sb_5__3_/chanx_right_in[6] sb_5__3_/chanx_right_in[7]
+ sb_5__3_/chanx_right_in[8] sb_5__3_/chanx_right_in[9] sb_6__3_/chanx_left_out[0]
+ sb_6__3_/chanx_left_out[10] sb_6__3_/chanx_left_out[11] sb_6__3_/chanx_left_out[12]
+ sb_6__3_/chanx_left_out[13] sb_6__3_/chanx_left_out[14] sb_6__3_/chanx_left_out[15]
+ sb_6__3_/chanx_left_out[16] sb_6__3_/chanx_left_out[17] sb_6__3_/chanx_left_out[18]
+ sb_6__3_/chanx_left_out[19] sb_6__3_/chanx_left_out[1] sb_6__3_/chanx_left_out[2]
+ sb_6__3_/chanx_left_out[3] sb_6__3_/chanx_left_out[4] sb_6__3_/chanx_left_out[5]
+ sb_6__3_/chanx_left_out[6] sb_6__3_/chanx_left_out[7] sb_6__3_/chanx_left_out[8]
+ sb_6__3_/chanx_left_out[9] sb_6__3_/chanx_left_in[0] sb_6__3_/chanx_left_in[10]
+ sb_6__3_/chanx_left_in[11] sb_6__3_/chanx_left_in[12] sb_6__3_/chanx_left_in[13]
+ sb_6__3_/chanx_left_in[14] sb_6__3_/chanx_left_in[15] sb_6__3_/chanx_left_in[16]
+ sb_6__3_/chanx_left_in[17] sb_6__3_/chanx_left_in[18] sb_6__3_/chanx_left_in[19]
+ sb_6__3_/chanx_left_in[1] sb_6__3_/chanx_left_in[2] sb_6__3_/chanx_left_in[3] sb_6__3_/chanx_left_in[4]
+ sb_6__3_/chanx_left_in[5] sb_6__3_/chanx_left_in[6] sb_6__3_/chanx_left_in[7] sb_6__3_/chanx_left_in[8]
+ sb_6__3_/chanx_left_in[9] cbx_6__3_/clk_1_N_out cbx_6__3_/clk_1_S_out sb_5__3_/clk_1_E_out
+ cbx_6__3_/clk_2_E_out cbx_6__3_/clk_2_W_in cbx_6__3_/clk_2_W_out cbx_6__3_/clk_3_E_out
+ cbx_6__3_/clk_3_W_in cbx_6__3_/clk_3_W_out cbx_6__3_/prog_clk_0_N_in cbx_6__3_/prog_clk_0_W_out
+ cbx_6__3_/prog_clk_1_N_out cbx_6__3_/prog_clk_1_S_out sb_5__3_/prog_clk_1_E_out
+ cbx_6__3_/prog_clk_2_E_out cbx_6__3_/prog_clk_2_W_in cbx_6__3_/prog_clk_2_W_out
+ cbx_6__3_/prog_clk_3_E_out cbx_6__3_/prog_clk_3_W_in cbx_6__3_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_6__8_ sb_6__8_/SC_IN_BOT sb_6__8_/SC_OUT_BOT VGND VPWR sb_6__8_/bottom_left_grid_pin_42_
+ sb_6__8_/bottom_left_grid_pin_43_ sb_6__8_/bottom_left_grid_pin_44_ sb_6__8_/bottom_left_grid_pin_45_
+ sb_6__8_/bottom_left_grid_pin_46_ sb_6__8_/bottom_left_grid_pin_47_ sb_6__8_/bottom_left_grid_pin_48_
+ sb_6__8_/bottom_left_grid_pin_49_ sb_6__8_/ccff_head sb_6__8_/ccff_tail sb_6__8_/chanx_left_in[0]
+ sb_6__8_/chanx_left_in[10] sb_6__8_/chanx_left_in[11] sb_6__8_/chanx_left_in[12]
+ sb_6__8_/chanx_left_in[13] sb_6__8_/chanx_left_in[14] sb_6__8_/chanx_left_in[15]
+ sb_6__8_/chanx_left_in[16] sb_6__8_/chanx_left_in[17] sb_6__8_/chanx_left_in[18]
+ sb_6__8_/chanx_left_in[19] sb_6__8_/chanx_left_in[1] sb_6__8_/chanx_left_in[2] sb_6__8_/chanx_left_in[3]
+ sb_6__8_/chanx_left_in[4] sb_6__8_/chanx_left_in[5] sb_6__8_/chanx_left_in[6] sb_6__8_/chanx_left_in[7]
+ sb_6__8_/chanx_left_in[8] sb_6__8_/chanx_left_in[9] sb_6__8_/chanx_left_out[0] sb_6__8_/chanx_left_out[10]
+ sb_6__8_/chanx_left_out[11] sb_6__8_/chanx_left_out[12] sb_6__8_/chanx_left_out[13]
+ sb_6__8_/chanx_left_out[14] sb_6__8_/chanx_left_out[15] sb_6__8_/chanx_left_out[16]
+ sb_6__8_/chanx_left_out[17] sb_6__8_/chanx_left_out[18] sb_6__8_/chanx_left_out[19]
+ sb_6__8_/chanx_left_out[1] sb_6__8_/chanx_left_out[2] sb_6__8_/chanx_left_out[3]
+ sb_6__8_/chanx_left_out[4] sb_6__8_/chanx_left_out[5] sb_6__8_/chanx_left_out[6]
+ sb_6__8_/chanx_left_out[7] sb_6__8_/chanx_left_out[8] sb_6__8_/chanx_left_out[9]
+ sb_6__8_/chanx_right_in[0] sb_6__8_/chanx_right_in[10] sb_6__8_/chanx_right_in[11]
+ sb_6__8_/chanx_right_in[12] sb_6__8_/chanx_right_in[13] sb_6__8_/chanx_right_in[14]
+ sb_6__8_/chanx_right_in[15] sb_6__8_/chanx_right_in[16] sb_6__8_/chanx_right_in[17]
+ sb_6__8_/chanx_right_in[18] sb_6__8_/chanx_right_in[19] sb_6__8_/chanx_right_in[1]
+ sb_6__8_/chanx_right_in[2] sb_6__8_/chanx_right_in[3] sb_6__8_/chanx_right_in[4]
+ sb_6__8_/chanx_right_in[5] sb_6__8_/chanx_right_in[6] sb_6__8_/chanx_right_in[7]
+ sb_6__8_/chanx_right_in[8] sb_6__8_/chanx_right_in[9] cbx_7__8_/chanx_left_in[0]
+ cbx_7__8_/chanx_left_in[10] cbx_7__8_/chanx_left_in[11] cbx_7__8_/chanx_left_in[12]
+ cbx_7__8_/chanx_left_in[13] cbx_7__8_/chanx_left_in[14] cbx_7__8_/chanx_left_in[15]
+ cbx_7__8_/chanx_left_in[16] cbx_7__8_/chanx_left_in[17] cbx_7__8_/chanx_left_in[18]
+ cbx_7__8_/chanx_left_in[19] cbx_7__8_/chanx_left_in[1] cbx_7__8_/chanx_left_in[2]
+ cbx_7__8_/chanx_left_in[3] cbx_7__8_/chanx_left_in[4] cbx_7__8_/chanx_left_in[5]
+ cbx_7__8_/chanx_left_in[6] cbx_7__8_/chanx_left_in[7] cbx_7__8_/chanx_left_in[8]
+ cbx_7__8_/chanx_left_in[9] cby_6__8_/chany_top_out[0] cby_6__8_/chany_top_out[10]
+ cby_6__8_/chany_top_out[11] cby_6__8_/chany_top_out[12] cby_6__8_/chany_top_out[13]
+ cby_6__8_/chany_top_out[14] cby_6__8_/chany_top_out[15] cby_6__8_/chany_top_out[16]
+ cby_6__8_/chany_top_out[17] cby_6__8_/chany_top_out[18] cby_6__8_/chany_top_out[19]
+ cby_6__8_/chany_top_out[1] cby_6__8_/chany_top_out[2] cby_6__8_/chany_top_out[3]
+ cby_6__8_/chany_top_out[4] cby_6__8_/chany_top_out[5] cby_6__8_/chany_top_out[6]
+ cby_6__8_/chany_top_out[7] cby_6__8_/chany_top_out[8] cby_6__8_/chany_top_out[9]
+ cby_6__8_/chany_top_in[0] cby_6__8_/chany_top_in[10] cby_6__8_/chany_top_in[11]
+ cby_6__8_/chany_top_in[12] cby_6__8_/chany_top_in[13] cby_6__8_/chany_top_in[14]
+ cby_6__8_/chany_top_in[15] cby_6__8_/chany_top_in[16] cby_6__8_/chany_top_in[17]
+ cby_6__8_/chany_top_in[18] cby_6__8_/chany_top_in[19] cby_6__8_/chany_top_in[1]
+ cby_6__8_/chany_top_in[2] cby_6__8_/chany_top_in[3] cby_6__8_/chany_top_in[4] cby_6__8_/chany_top_in[5]
+ cby_6__8_/chany_top_in[6] cby_6__8_/chany_top_in[7] cby_6__8_/chany_top_in[8] cby_6__8_/chany_top_in[9]
+ sb_6__8_/left_bottom_grid_pin_34_ sb_6__8_/left_bottom_grid_pin_35_ sb_6__8_/left_bottom_grid_pin_36_
+ sb_6__8_/left_bottom_grid_pin_37_ sb_6__8_/left_bottom_grid_pin_38_ sb_6__8_/left_bottom_grid_pin_39_
+ sb_6__8_/left_bottom_grid_pin_40_ sb_6__8_/left_bottom_grid_pin_41_ sb_6__8_/left_top_grid_pin_1_
+ sb_6__8_/prog_clk_0_S_in sb_6__8_/right_bottom_grid_pin_34_ sb_6__8_/right_bottom_grid_pin_35_
+ sb_6__8_/right_bottom_grid_pin_36_ sb_6__8_/right_bottom_grid_pin_37_ sb_6__8_/right_bottom_grid_pin_38_
+ sb_6__8_/right_bottom_grid_pin_39_ sb_6__8_/right_bottom_grid_pin_40_ sb_6__8_/right_bottom_grid_pin_41_
+ sb_6__8_/right_top_grid_pin_1_ sb_1__2_
Xgrid_clb_8__6_ cbx_8__5_/SC_OUT_TOP grid_clb_8__6_/SC_OUT_BOT cbx_8__6_/SC_IN_BOT
+ cby_7__6_/Test_en_E_out grid_clb_8__6_/Test_en_E_out cby_7__6_/Test_en_E_out grid_clb_8__6_/Test_en_W_out
+ VGND VPWR cbx_8__5_/REGIN_FEEDTHROUGH grid_clb_8__6_/bottom_width_0_height_0__pin_51_
+ cby_7__6_/ccff_tail cby_8__6_/ccff_head cbx_8__5_/clk_1_N_out cbx_8__5_/clk_1_N_out
+ cby_8__6_/prog_clk_0_W_in cbx_8__5_/prog_clk_1_N_out grid_clb_8__6_/prog_clk_0_N_out
+ cbx_8__5_/prog_clk_1_N_out cbx_8__5_/prog_clk_0_N_in grid_clb_8__6_/prog_clk_0_W_out
+ cby_8__6_/left_grid_pin_16_ cby_8__6_/left_grid_pin_17_ cby_8__6_/left_grid_pin_18_
+ cby_8__6_/left_grid_pin_19_ cby_8__6_/left_grid_pin_20_ cby_8__6_/left_grid_pin_21_
+ cby_8__6_/left_grid_pin_22_ cby_8__6_/left_grid_pin_23_ cby_8__6_/left_grid_pin_24_
+ cby_8__6_/left_grid_pin_25_ cby_8__6_/left_grid_pin_26_ cby_8__6_/left_grid_pin_27_
+ cby_8__6_/left_grid_pin_28_ cby_8__6_/left_grid_pin_29_ cby_8__6_/left_grid_pin_30_
+ cby_8__6_/left_grid_pin_31_ sb_8__5_/top_left_grid_pin_42_ sb_8__6_/bottom_left_grid_pin_42_
+ sb_8__5_/top_left_grid_pin_43_ sb_8__6_/bottom_left_grid_pin_43_ sb_8__5_/top_left_grid_pin_44_
+ sb_8__6_/bottom_left_grid_pin_44_ sb_8__5_/top_left_grid_pin_45_ sb_8__6_/bottom_left_grid_pin_45_
+ sb_8__5_/top_left_grid_pin_46_ sb_8__6_/bottom_left_grid_pin_46_ sb_8__5_/top_left_grid_pin_47_
+ sb_8__6_/bottom_left_grid_pin_47_ sb_8__5_/top_left_grid_pin_48_ sb_8__6_/bottom_left_grid_pin_48_
+ sb_8__5_/top_left_grid_pin_49_ sb_8__6_/bottom_left_grid_pin_49_ cbx_8__6_/bottom_grid_pin_0_
+ cbx_8__6_/bottom_grid_pin_10_ cbx_8__6_/bottom_grid_pin_11_ cbx_8__6_/bottom_grid_pin_12_
+ cbx_8__6_/bottom_grid_pin_13_ cbx_8__6_/bottom_grid_pin_14_ cbx_8__6_/bottom_grid_pin_15_
+ cbx_8__6_/bottom_grid_pin_1_ cbx_8__6_/bottom_grid_pin_2_ cbx_8__6_/REGOUT_FEEDTHROUGH
+ grid_clb_8__6_/top_width_0_height_0__pin_33_ sb_8__6_/left_bottom_grid_pin_34_ sb_7__6_/right_bottom_grid_pin_34_
+ sb_8__6_/left_bottom_grid_pin_35_ sb_7__6_/right_bottom_grid_pin_35_ sb_8__6_/left_bottom_grid_pin_36_
+ sb_7__6_/right_bottom_grid_pin_36_ sb_8__6_/left_bottom_grid_pin_37_ sb_7__6_/right_bottom_grid_pin_37_
+ sb_8__6_/left_bottom_grid_pin_38_ sb_7__6_/right_bottom_grid_pin_38_ sb_8__6_/left_bottom_grid_pin_39_
+ sb_7__6_/right_bottom_grid_pin_39_ cbx_8__6_/bottom_grid_pin_3_ sb_8__6_/left_bottom_grid_pin_40_
+ sb_7__6_/right_bottom_grid_pin_40_ sb_8__6_/left_bottom_grid_pin_41_ sb_7__6_/right_bottom_grid_pin_41_
+ cbx_8__6_/bottom_grid_pin_4_ cbx_8__6_/bottom_grid_pin_5_ cbx_8__6_/bottom_grid_pin_6_
+ cbx_8__6_/bottom_grid_pin_7_ cbx_8__6_/bottom_grid_pin_8_ cbx_8__6_/bottom_grid_pin_9_
+ grid_clb
Xcbx_3__0_ IO_ISOL_N cbx_3__0_/SC_IN_BOT cbx_3__0_/SC_IN_TOP sb_3__0_/SC_IN_TOP cbx_3__0_/SC_OUT_TOP
+ VGND VPWR cbx_3__0_/bottom_grid_pin_0_ cbx_3__0_/bottom_grid_pin_10_ cbx_3__0_/bottom_grid_pin_12_
+ cbx_3__0_/bottom_grid_pin_14_ cbx_3__0_/bottom_grid_pin_16_ cbx_3__0_/bottom_grid_pin_2_
+ cbx_3__0_/bottom_grid_pin_4_ cbx_3__0_/bottom_grid_pin_6_ cbx_3__0_/bottom_grid_pin_8_
+ sb_3__0_/ccff_tail sb_2__0_/ccff_head cbx_3__0_/chanx_left_in[0] cbx_3__0_/chanx_left_in[10]
+ cbx_3__0_/chanx_left_in[11] cbx_3__0_/chanx_left_in[12] cbx_3__0_/chanx_left_in[13]
+ cbx_3__0_/chanx_left_in[14] cbx_3__0_/chanx_left_in[15] cbx_3__0_/chanx_left_in[16]
+ cbx_3__0_/chanx_left_in[17] cbx_3__0_/chanx_left_in[18] cbx_3__0_/chanx_left_in[19]
+ cbx_3__0_/chanx_left_in[1] cbx_3__0_/chanx_left_in[2] cbx_3__0_/chanx_left_in[3]
+ cbx_3__0_/chanx_left_in[4] cbx_3__0_/chanx_left_in[5] cbx_3__0_/chanx_left_in[6]
+ cbx_3__0_/chanx_left_in[7] cbx_3__0_/chanx_left_in[8] cbx_3__0_/chanx_left_in[9]
+ sb_2__0_/chanx_right_in[0] sb_2__0_/chanx_right_in[10] sb_2__0_/chanx_right_in[11]
+ sb_2__0_/chanx_right_in[12] sb_2__0_/chanx_right_in[13] sb_2__0_/chanx_right_in[14]
+ sb_2__0_/chanx_right_in[15] sb_2__0_/chanx_right_in[16] sb_2__0_/chanx_right_in[17]
+ sb_2__0_/chanx_right_in[18] sb_2__0_/chanx_right_in[19] sb_2__0_/chanx_right_in[1]
+ sb_2__0_/chanx_right_in[2] sb_2__0_/chanx_right_in[3] sb_2__0_/chanx_right_in[4]
+ sb_2__0_/chanx_right_in[5] sb_2__0_/chanx_right_in[6] sb_2__0_/chanx_right_in[7]
+ sb_2__0_/chanx_right_in[8] sb_2__0_/chanx_right_in[9] sb_3__0_/chanx_left_out[0]
+ sb_3__0_/chanx_left_out[10] sb_3__0_/chanx_left_out[11] sb_3__0_/chanx_left_out[12]
+ sb_3__0_/chanx_left_out[13] sb_3__0_/chanx_left_out[14] sb_3__0_/chanx_left_out[15]
+ sb_3__0_/chanx_left_out[16] sb_3__0_/chanx_left_out[17] sb_3__0_/chanx_left_out[18]
+ sb_3__0_/chanx_left_out[19] sb_3__0_/chanx_left_out[1] sb_3__0_/chanx_left_out[2]
+ sb_3__0_/chanx_left_out[3] sb_3__0_/chanx_left_out[4] sb_3__0_/chanx_left_out[5]
+ sb_3__0_/chanx_left_out[6] sb_3__0_/chanx_left_out[7] sb_3__0_/chanx_left_out[8]
+ sb_3__0_/chanx_left_out[9] sb_3__0_/chanx_left_in[0] sb_3__0_/chanx_left_in[10]
+ sb_3__0_/chanx_left_in[11] sb_3__0_/chanx_left_in[12] sb_3__0_/chanx_left_in[13]
+ sb_3__0_/chanx_left_in[14] sb_3__0_/chanx_left_in[15] sb_3__0_/chanx_left_in[16]
+ sb_3__0_/chanx_left_in[17] sb_3__0_/chanx_left_in[18] sb_3__0_/chanx_left_in[19]
+ sb_3__0_/chanx_left_in[1] sb_3__0_/chanx_left_in[2] sb_3__0_/chanx_left_in[3] sb_3__0_/chanx_left_in[4]
+ sb_3__0_/chanx_left_in[5] sb_3__0_/chanx_left_in[6] sb_3__0_/chanx_left_in[7] sb_3__0_/chanx_left_in[8]
+ sb_3__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69] cbx_3__0_/prog_clk_0_N_in cbx_3__0_/prog_clk_0_W_out
+ cbx_3__0_/bottom_grid_pin_0_ cbx_3__0_/bottom_grid_pin_10_ sb_3__0_/left_bottom_grid_pin_11_
+ sb_2__0_/right_bottom_grid_pin_11_ cbx_3__0_/bottom_grid_pin_12_ sb_3__0_/left_bottom_grid_pin_13_
+ sb_2__0_/right_bottom_grid_pin_13_ cbx_3__0_/bottom_grid_pin_14_ sb_3__0_/left_bottom_grid_pin_15_
+ sb_2__0_/right_bottom_grid_pin_15_ cbx_3__0_/bottom_grid_pin_16_ sb_3__0_/left_bottom_grid_pin_17_
+ sb_2__0_/right_bottom_grid_pin_17_ sb_3__0_/left_bottom_grid_pin_1_ sb_2__0_/right_bottom_grid_pin_1_
+ cbx_3__0_/bottom_grid_pin_2_ sb_3__0_/left_bottom_grid_pin_3_ sb_2__0_/right_bottom_grid_pin_3_
+ cbx_3__0_/bottom_grid_pin_4_ sb_3__0_/left_bottom_grid_pin_5_ sb_2__0_/right_bottom_grid_pin_5_
+ cbx_3__0_/bottom_grid_pin_6_ sb_3__0_/left_bottom_grid_pin_7_ sb_2__0_/right_bottom_grid_pin_7_
+ cbx_3__0_/bottom_grid_pin_8_ sb_3__0_/left_bottom_grid_pin_9_ sb_2__0_/right_bottom_grid_pin_9_
+ cbx_1__0_
Xgrid_clb_5__3_ cbx_5__3_/SC_OUT_BOT cbx_5__2_/SC_IN_TOP grid_clb_5__3_/SC_OUT_TOP
+ cby_4__3_/Test_en_E_out cby_5__3_/Test_en_W_in cby_4__3_/Test_en_E_out grid_clb_5__3_/Test_en_W_out
+ VGND VPWR cbx_5__2_/REGIN_FEEDTHROUGH grid_clb_5__3_/bottom_width_0_height_0__pin_51_
+ cby_4__3_/ccff_tail cby_5__3_/ccff_head cbx_5__3_/clk_1_S_out cbx_5__3_/clk_1_S_out
+ cby_5__3_/prog_clk_0_W_in cbx_5__3_/prog_clk_1_S_out grid_clb_5__3_/prog_clk_0_N_out
+ cbx_5__3_/prog_clk_1_S_out cbx_5__2_/prog_clk_0_N_in grid_clb_5__3_/prog_clk_0_W_out
+ cby_5__3_/left_grid_pin_16_ cby_5__3_/left_grid_pin_17_ cby_5__3_/left_grid_pin_18_
+ cby_5__3_/left_grid_pin_19_ cby_5__3_/left_grid_pin_20_ cby_5__3_/left_grid_pin_21_
+ cby_5__3_/left_grid_pin_22_ cby_5__3_/left_grid_pin_23_ cby_5__3_/left_grid_pin_24_
+ cby_5__3_/left_grid_pin_25_ cby_5__3_/left_grid_pin_26_ cby_5__3_/left_grid_pin_27_
+ cby_5__3_/left_grid_pin_28_ cby_5__3_/left_grid_pin_29_ cby_5__3_/left_grid_pin_30_
+ cby_5__3_/left_grid_pin_31_ sb_5__2_/top_left_grid_pin_42_ sb_5__3_/bottom_left_grid_pin_42_
+ sb_5__2_/top_left_grid_pin_43_ sb_5__3_/bottom_left_grid_pin_43_ sb_5__2_/top_left_grid_pin_44_
+ sb_5__3_/bottom_left_grid_pin_44_ sb_5__2_/top_left_grid_pin_45_ sb_5__3_/bottom_left_grid_pin_45_
+ sb_5__2_/top_left_grid_pin_46_ sb_5__3_/bottom_left_grid_pin_46_ sb_5__2_/top_left_grid_pin_47_
+ sb_5__3_/bottom_left_grid_pin_47_ sb_5__2_/top_left_grid_pin_48_ sb_5__3_/bottom_left_grid_pin_48_
+ sb_5__2_/top_left_grid_pin_49_ sb_5__3_/bottom_left_grid_pin_49_ cbx_5__3_/bottom_grid_pin_0_
+ cbx_5__3_/bottom_grid_pin_10_ cbx_5__3_/bottom_grid_pin_11_ cbx_5__3_/bottom_grid_pin_12_
+ cbx_5__3_/bottom_grid_pin_13_ cbx_5__3_/bottom_grid_pin_14_ cbx_5__3_/bottom_grid_pin_15_
+ cbx_5__3_/bottom_grid_pin_1_ cbx_5__3_/bottom_grid_pin_2_ cbx_5__3_/REGOUT_FEEDTHROUGH
+ grid_clb_5__3_/top_width_0_height_0__pin_33_ sb_5__3_/left_bottom_grid_pin_34_ sb_4__3_/right_bottom_grid_pin_34_
+ sb_5__3_/left_bottom_grid_pin_35_ sb_4__3_/right_bottom_grid_pin_35_ sb_5__3_/left_bottom_grid_pin_36_
+ sb_4__3_/right_bottom_grid_pin_36_ sb_5__3_/left_bottom_grid_pin_37_ sb_4__3_/right_bottom_grid_pin_37_
+ sb_5__3_/left_bottom_grid_pin_38_ sb_4__3_/right_bottom_grid_pin_38_ sb_5__3_/left_bottom_grid_pin_39_
+ sb_4__3_/right_bottom_grid_pin_39_ cbx_5__3_/bottom_grid_pin_3_ sb_5__3_/left_bottom_grid_pin_40_
+ sb_4__3_/right_bottom_grid_pin_40_ sb_5__3_/left_bottom_grid_pin_41_ sb_4__3_/right_bottom_grid_pin_41_
+ cbx_5__3_/bottom_grid_pin_4_ cbx_5__3_/bottom_grid_pin_5_ cbx_5__3_/bottom_grid_pin_6_
+ cbx_5__3_/bottom_grid_pin_7_ cbx_5__3_/bottom_grid_pin_8_ cbx_5__3_/bottom_grid_pin_9_
+ grid_clb
Xsb_3__5_ sb_3__5_/Test_en_N_out sb_3__5_/Test_en_S_in VGND VPWR sb_3__5_/bottom_left_grid_pin_42_
+ sb_3__5_/bottom_left_grid_pin_43_ sb_3__5_/bottom_left_grid_pin_44_ sb_3__5_/bottom_left_grid_pin_45_
+ sb_3__5_/bottom_left_grid_pin_46_ sb_3__5_/bottom_left_grid_pin_47_ sb_3__5_/bottom_left_grid_pin_48_
+ sb_3__5_/bottom_left_grid_pin_49_ sb_3__5_/ccff_head sb_3__5_/ccff_tail sb_3__5_/chanx_left_in[0]
+ sb_3__5_/chanx_left_in[10] sb_3__5_/chanx_left_in[11] sb_3__5_/chanx_left_in[12]
+ sb_3__5_/chanx_left_in[13] sb_3__5_/chanx_left_in[14] sb_3__5_/chanx_left_in[15]
+ sb_3__5_/chanx_left_in[16] sb_3__5_/chanx_left_in[17] sb_3__5_/chanx_left_in[18]
+ sb_3__5_/chanx_left_in[19] sb_3__5_/chanx_left_in[1] sb_3__5_/chanx_left_in[2] sb_3__5_/chanx_left_in[3]
+ sb_3__5_/chanx_left_in[4] sb_3__5_/chanx_left_in[5] sb_3__5_/chanx_left_in[6] sb_3__5_/chanx_left_in[7]
+ sb_3__5_/chanx_left_in[8] sb_3__5_/chanx_left_in[9] sb_3__5_/chanx_left_out[0] sb_3__5_/chanx_left_out[10]
+ sb_3__5_/chanx_left_out[11] sb_3__5_/chanx_left_out[12] sb_3__5_/chanx_left_out[13]
+ sb_3__5_/chanx_left_out[14] sb_3__5_/chanx_left_out[15] sb_3__5_/chanx_left_out[16]
+ sb_3__5_/chanx_left_out[17] sb_3__5_/chanx_left_out[18] sb_3__5_/chanx_left_out[19]
+ sb_3__5_/chanx_left_out[1] sb_3__5_/chanx_left_out[2] sb_3__5_/chanx_left_out[3]
+ sb_3__5_/chanx_left_out[4] sb_3__5_/chanx_left_out[5] sb_3__5_/chanx_left_out[6]
+ sb_3__5_/chanx_left_out[7] sb_3__5_/chanx_left_out[8] sb_3__5_/chanx_left_out[9]
+ sb_3__5_/chanx_right_in[0] sb_3__5_/chanx_right_in[10] sb_3__5_/chanx_right_in[11]
+ sb_3__5_/chanx_right_in[12] sb_3__5_/chanx_right_in[13] sb_3__5_/chanx_right_in[14]
+ sb_3__5_/chanx_right_in[15] sb_3__5_/chanx_right_in[16] sb_3__5_/chanx_right_in[17]
+ sb_3__5_/chanx_right_in[18] sb_3__5_/chanx_right_in[19] sb_3__5_/chanx_right_in[1]
+ sb_3__5_/chanx_right_in[2] sb_3__5_/chanx_right_in[3] sb_3__5_/chanx_right_in[4]
+ sb_3__5_/chanx_right_in[5] sb_3__5_/chanx_right_in[6] sb_3__5_/chanx_right_in[7]
+ sb_3__5_/chanx_right_in[8] sb_3__5_/chanx_right_in[9] cbx_4__5_/chanx_left_in[0]
+ cbx_4__5_/chanx_left_in[10] cbx_4__5_/chanx_left_in[11] cbx_4__5_/chanx_left_in[12]
+ cbx_4__5_/chanx_left_in[13] cbx_4__5_/chanx_left_in[14] cbx_4__5_/chanx_left_in[15]
+ cbx_4__5_/chanx_left_in[16] cbx_4__5_/chanx_left_in[17] cbx_4__5_/chanx_left_in[18]
+ cbx_4__5_/chanx_left_in[19] cbx_4__5_/chanx_left_in[1] cbx_4__5_/chanx_left_in[2]
+ cbx_4__5_/chanx_left_in[3] cbx_4__5_/chanx_left_in[4] cbx_4__5_/chanx_left_in[5]
+ cbx_4__5_/chanx_left_in[6] cbx_4__5_/chanx_left_in[7] cbx_4__5_/chanx_left_in[8]
+ cbx_4__5_/chanx_left_in[9] cby_3__5_/chany_top_out[0] cby_3__5_/chany_top_out[10]
+ cby_3__5_/chany_top_out[11] cby_3__5_/chany_top_out[12] cby_3__5_/chany_top_out[13]
+ cby_3__5_/chany_top_out[14] cby_3__5_/chany_top_out[15] cby_3__5_/chany_top_out[16]
+ cby_3__5_/chany_top_out[17] cby_3__5_/chany_top_out[18] cby_3__5_/chany_top_out[19]
+ cby_3__5_/chany_top_out[1] cby_3__5_/chany_top_out[2] cby_3__5_/chany_top_out[3]
+ cby_3__5_/chany_top_out[4] cby_3__5_/chany_top_out[5] cby_3__5_/chany_top_out[6]
+ cby_3__5_/chany_top_out[7] cby_3__5_/chany_top_out[8] cby_3__5_/chany_top_out[9]
+ cby_3__5_/chany_top_in[0] cby_3__5_/chany_top_in[10] cby_3__5_/chany_top_in[11]
+ cby_3__5_/chany_top_in[12] cby_3__5_/chany_top_in[13] cby_3__5_/chany_top_in[14]
+ cby_3__5_/chany_top_in[15] cby_3__5_/chany_top_in[16] cby_3__5_/chany_top_in[17]
+ cby_3__5_/chany_top_in[18] cby_3__5_/chany_top_in[19] cby_3__5_/chany_top_in[1]
+ cby_3__5_/chany_top_in[2] cby_3__5_/chany_top_in[3] cby_3__5_/chany_top_in[4] cby_3__5_/chany_top_in[5]
+ cby_3__5_/chany_top_in[6] cby_3__5_/chany_top_in[7] cby_3__5_/chany_top_in[8] cby_3__5_/chany_top_in[9]
+ sb_3__5_/chany_top_in[0] sb_3__5_/chany_top_in[10] sb_3__5_/chany_top_in[11] sb_3__5_/chany_top_in[12]
+ sb_3__5_/chany_top_in[13] sb_3__5_/chany_top_in[14] sb_3__5_/chany_top_in[15] sb_3__5_/chany_top_in[16]
+ sb_3__5_/chany_top_in[17] sb_3__5_/chany_top_in[18] sb_3__5_/chany_top_in[19] sb_3__5_/chany_top_in[1]
+ sb_3__5_/chany_top_in[2] sb_3__5_/chany_top_in[3] sb_3__5_/chany_top_in[4] sb_3__5_/chany_top_in[5]
+ sb_3__5_/chany_top_in[6] sb_3__5_/chany_top_in[7] sb_3__5_/chany_top_in[8] sb_3__5_/chany_top_in[9]
+ sb_3__5_/chany_top_out[0] sb_3__5_/chany_top_out[10] sb_3__5_/chany_top_out[11]
+ sb_3__5_/chany_top_out[12] sb_3__5_/chany_top_out[13] sb_3__5_/chany_top_out[14]
+ sb_3__5_/chany_top_out[15] sb_3__5_/chany_top_out[16] sb_3__5_/chany_top_out[17]
+ sb_3__5_/chany_top_out[18] sb_3__5_/chany_top_out[19] sb_3__5_/chany_top_out[1]
+ sb_3__5_/chany_top_out[2] sb_3__5_/chany_top_out[3] sb_3__5_/chany_top_out[4] sb_3__5_/chany_top_out[5]
+ sb_3__5_/chany_top_out[6] sb_3__5_/chany_top_out[7] sb_3__5_/chany_top_out[8] sb_3__5_/chany_top_out[9]
+ sb_3__5_/clk_1_E_out sb_3__5_/clk_1_N_in sb_3__5_/clk_1_W_out sb_3__5_/clk_2_E_out
+ sb_3__5_/clk_2_N_in sb_3__5_/clk_2_N_out sb_3__5_/clk_2_S_out sb_3__5_/clk_2_W_out
+ sb_3__5_/clk_3_E_out sb_3__5_/clk_3_N_in sb_3__5_/clk_3_N_out sb_3__5_/clk_3_S_out
+ sb_3__5_/clk_3_W_out sb_3__5_/left_bottom_grid_pin_34_ sb_3__5_/left_bottom_grid_pin_35_
+ sb_3__5_/left_bottom_grid_pin_36_ sb_3__5_/left_bottom_grid_pin_37_ sb_3__5_/left_bottom_grid_pin_38_
+ sb_3__5_/left_bottom_grid_pin_39_ sb_3__5_/left_bottom_grid_pin_40_ sb_3__5_/left_bottom_grid_pin_41_
+ sb_3__5_/prog_clk_0_N_in sb_3__5_/prog_clk_1_E_out sb_3__5_/prog_clk_1_N_in sb_3__5_/prog_clk_1_W_out
+ sb_3__5_/prog_clk_2_E_out sb_3__5_/prog_clk_2_N_in sb_3__5_/prog_clk_2_N_out sb_3__5_/prog_clk_2_S_out
+ sb_3__5_/prog_clk_2_W_out sb_3__5_/prog_clk_3_E_out sb_3__5_/prog_clk_3_N_in sb_3__5_/prog_clk_3_N_out
+ sb_3__5_/prog_clk_3_S_out sb_3__5_/prog_clk_3_W_out sb_3__5_/right_bottom_grid_pin_34_
+ sb_3__5_/right_bottom_grid_pin_35_ sb_3__5_/right_bottom_grid_pin_36_ sb_3__5_/right_bottom_grid_pin_37_
+ sb_3__5_/right_bottom_grid_pin_38_ sb_3__5_/right_bottom_grid_pin_39_ sb_3__5_/right_bottom_grid_pin_40_
+ sb_3__5_/right_bottom_grid_pin_41_ sb_3__5_/top_left_grid_pin_42_ sb_3__5_/top_left_grid_pin_43_
+ sb_3__5_/top_left_grid_pin_44_ sb_3__5_/top_left_grid_pin_45_ sb_3__5_/top_left_grid_pin_46_
+ sb_3__5_/top_left_grid_pin_47_ sb_3__5_/top_left_grid_pin_48_ sb_3__5_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_0__2_ VGND VPWR sb_0__2_/bottom_left_grid_pin_1_ sb_0__2_/ccff_head sb_0__2_/ccff_tail
+ sb_0__2_/chanx_right_in[0] sb_0__2_/chanx_right_in[10] sb_0__2_/chanx_right_in[11]
+ sb_0__2_/chanx_right_in[12] sb_0__2_/chanx_right_in[13] sb_0__2_/chanx_right_in[14]
+ sb_0__2_/chanx_right_in[15] sb_0__2_/chanx_right_in[16] sb_0__2_/chanx_right_in[17]
+ sb_0__2_/chanx_right_in[18] sb_0__2_/chanx_right_in[19] sb_0__2_/chanx_right_in[1]
+ sb_0__2_/chanx_right_in[2] sb_0__2_/chanx_right_in[3] sb_0__2_/chanx_right_in[4]
+ sb_0__2_/chanx_right_in[5] sb_0__2_/chanx_right_in[6] sb_0__2_/chanx_right_in[7]
+ sb_0__2_/chanx_right_in[8] sb_0__2_/chanx_right_in[9] cbx_1__2_/chanx_left_in[0]
+ cbx_1__2_/chanx_left_in[10] cbx_1__2_/chanx_left_in[11] cbx_1__2_/chanx_left_in[12]
+ cbx_1__2_/chanx_left_in[13] cbx_1__2_/chanx_left_in[14] cbx_1__2_/chanx_left_in[15]
+ cbx_1__2_/chanx_left_in[16] cbx_1__2_/chanx_left_in[17] cbx_1__2_/chanx_left_in[18]
+ cbx_1__2_/chanx_left_in[19] cbx_1__2_/chanx_left_in[1] cbx_1__2_/chanx_left_in[2]
+ cbx_1__2_/chanx_left_in[3] cbx_1__2_/chanx_left_in[4] cbx_1__2_/chanx_left_in[5]
+ cbx_1__2_/chanx_left_in[6] cbx_1__2_/chanx_left_in[7] cbx_1__2_/chanx_left_in[8]
+ cbx_1__2_/chanx_left_in[9] cby_0__2_/chany_top_out[0] cby_0__2_/chany_top_out[10]
+ cby_0__2_/chany_top_out[11] cby_0__2_/chany_top_out[12] cby_0__2_/chany_top_out[13]
+ cby_0__2_/chany_top_out[14] cby_0__2_/chany_top_out[15] cby_0__2_/chany_top_out[16]
+ cby_0__2_/chany_top_out[17] cby_0__2_/chany_top_out[18] cby_0__2_/chany_top_out[19]
+ cby_0__2_/chany_top_out[1] cby_0__2_/chany_top_out[2] cby_0__2_/chany_top_out[3]
+ cby_0__2_/chany_top_out[4] cby_0__2_/chany_top_out[5] cby_0__2_/chany_top_out[6]
+ cby_0__2_/chany_top_out[7] cby_0__2_/chany_top_out[8] cby_0__2_/chany_top_out[9]
+ cby_0__2_/chany_top_in[0] cby_0__2_/chany_top_in[10] cby_0__2_/chany_top_in[11]
+ cby_0__2_/chany_top_in[12] cby_0__2_/chany_top_in[13] cby_0__2_/chany_top_in[14]
+ cby_0__2_/chany_top_in[15] cby_0__2_/chany_top_in[16] cby_0__2_/chany_top_in[17]
+ cby_0__2_/chany_top_in[18] cby_0__2_/chany_top_in[19] cby_0__2_/chany_top_in[1]
+ cby_0__2_/chany_top_in[2] cby_0__2_/chany_top_in[3] cby_0__2_/chany_top_in[4] cby_0__2_/chany_top_in[5]
+ cby_0__2_/chany_top_in[6] cby_0__2_/chany_top_in[7] cby_0__2_/chany_top_in[8] cby_0__2_/chany_top_in[9]
+ sb_0__2_/chany_top_in[0] sb_0__2_/chany_top_in[10] sb_0__2_/chany_top_in[11] sb_0__2_/chany_top_in[12]
+ sb_0__2_/chany_top_in[13] sb_0__2_/chany_top_in[14] sb_0__2_/chany_top_in[15] sb_0__2_/chany_top_in[16]
+ sb_0__2_/chany_top_in[17] sb_0__2_/chany_top_in[18] sb_0__2_/chany_top_in[19] sb_0__2_/chany_top_in[1]
+ sb_0__2_/chany_top_in[2] sb_0__2_/chany_top_in[3] sb_0__2_/chany_top_in[4] sb_0__2_/chany_top_in[5]
+ sb_0__2_/chany_top_in[6] sb_0__2_/chany_top_in[7] sb_0__2_/chany_top_in[8] sb_0__2_/chany_top_in[9]
+ sb_0__2_/chany_top_out[0] sb_0__2_/chany_top_out[10] sb_0__2_/chany_top_out[11]
+ sb_0__2_/chany_top_out[12] sb_0__2_/chany_top_out[13] sb_0__2_/chany_top_out[14]
+ sb_0__2_/chany_top_out[15] sb_0__2_/chany_top_out[16] sb_0__2_/chany_top_out[17]
+ sb_0__2_/chany_top_out[18] sb_0__2_/chany_top_out[19] sb_0__2_/chany_top_out[1]
+ sb_0__2_/chany_top_out[2] sb_0__2_/chany_top_out[3] sb_0__2_/chany_top_out[4] sb_0__2_/chany_top_out[5]
+ sb_0__2_/chany_top_out[6] sb_0__2_/chany_top_out[7] sb_0__2_/chany_top_out[8] sb_0__2_/chany_top_out[9]
+ sb_0__2_/prog_clk_0_E_in sb_0__2_/right_bottom_grid_pin_34_ sb_0__2_/right_bottom_grid_pin_35_
+ sb_0__2_/right_bottom_grid_pin_36_ sb_0__2_/right_bottom_grid_pin_37_ sb_0__2_/right_bottom_grid_pin_38_
+ sb_0__2_/right_bottom_grid_pin_39_ sb_0__2_/right_bottom_grid_pin_40_ sb_0__2_/right_bottom_grid_pin_41_
+ sb_0__2_/top_left_grid_pin_1_ sb_0__1_
Xcby_6__1_ cby_6__1_/Test_en_W_in cby_6__1_/Test_en_E_out cby_6__1_/Test_en_N_out
+ cby_6__1_/Test_en_W_in cby_6__1_/Test_en_W_in cby_6__1_/Test_en_W_out VGND VPWR
+ cby_6__1_/ccff_head cby_6__1_/ccff_tail sb_6__0_/chany_top_out[0] sb_6__0_/chany_top_out[10]
+ sb_6__0_/chany_top_out[11] sb_6__0_/chany_top_out[12] sb_6__0_/chany_top_out[13]
+ sb_6__0_/chany_top_out[14] sb_6__0_/chany_top_out[15] sb_6__0_/chany_top_out[16]
+ sb_6__0_/chany_top_out[17] sb_6__0_/chany_top_out[18] sb_6__0_/chany_top_out[19]
+ sb_6__0_/chany_top_out[1] sb_6__0_/chany_top_out[2] sb_6__0_/chany_top_out[3] sb_6__0_/chany_top_out[4]
+ sb_6__0_/chany_top_out[5] sb_6__0_/chany_top_out[6] sb_6__0_/chany_top_out[7] sb_6__0_/chany_top_out[8]
+ sb_6__0_/chany_top_out[9] sb_6__0_/chany_top_in[0] sb_6__0_/chany_top_in[10] sb_6__0_/chany_top_in[11]
+ sb_6__0_/chany_top_in[12] sb_6__0_/chany_top_in[13] sb_6__0_/chany_top_in[14] sb_6__0_/chany_top_in[15]
+ sb_6__0_/chany_top_in[16] sb_6__0_/chany_top_in[17] sb_6__0_/chany_top_in[18] sb_6__0_/chany_top_in[19]
+ sb_6__0_/chany_top_in[1] sb_6__0_/chany_top_in[2] sb_6__0_/chany_top_in[3] sb_6__0_/chany_top_in[4]
+ sb_6__0_/chany_top_in[5] sb_6__0_/chany_top_in[6] sb_6__0_/chany_top_in[7] sb_6__0_/chany_top_in[8]
+ sb_6__0_/chany_top_in[9] cby_6__1_/chany_top_in[0] cby_6__1_/chany_top_in[10] cby_6__1_/chany_top_in[11]
+ cby_6__1_/chany_top_in[12] cby_6__1_/chany_top_in[13] cby_6__1_/chany_top_in[14]
+ cby_6__1_/chany_top_in[15] cby_6__1_/chany_top_in[16] cby_6__1_/chany_top_in[17]
+ cby_6__1_/chany_top_in[18] cby_6__1_/chany_top_in[19] cby_6__1_/chany_top_in[1]
+ cby_6__1_/chany_top_in[2] cby_6__1_/chany_top_in[3] cby_6__1_/chany_top_in[4] cby_6__1_/chany_top_in[5]
+ cby_6__1_/chany_top_in[6] cby_6__1_/chany_top_in[7] cby_6__1_/chany_top_in[8] cby_6__1_/chany_top_in[9]
+ cby_6__1_/chany_top_out[0] cby_6__1_/chany_top_out[10] cby_6__1_/chany_top_out[11]
+ cby_6__1_/chany_top_out[12] cby_6__1_/chany_top_out[13] cby_6__1_/chany_top_out[14]
+ cby_6__1_/chany_top_out[15] cby_6__1_/chany_top_out[16] cby_6__1_/chany_top_out[17]
+ cby_6__1_/chany_top_out[18] cby_6__1_/chany_top_out[19] cby_6__1_/chany_top_out[1]
+ cby_6__1_/chany_top_out[2] cby_6__1_/chany_top_out[3] cby_6__1_/chany_top_out[4]
+ cby_6__1_/chany_top_out[5] cby_6__1_/chany_top_out[6] cby_6__1_/chany_top_out[7]
+ cby_6__1_/chany_top_out[8] cby_6__1_/chany_top_out[9] cby_6__1_/clk_2_N_out cby_6__1_/clk_2_S_in
+ cby_6__1_/clk_2_S_out cby_6__1_/clk_3_N_out cby_6__1_/clk_3_S_in cby_6__1_/clk_3_S_out
+ cby_6__1_/left_grid_pin_16_ cby_6__1_/left_grid_pin_17_ cby_6__1_/left_grid_pin_18_
+ cby_6__1_/left_grid_pin_19_ cby_6__1_/left_grid_pin_20_ cby_6__1_/left_grid_pin_21_
+ cby_6__1_/left_grid_pin_22_ cby_6__1_/left_grid_pin_23_ cby_6__1_/left_grid_pin_24_
+ cby_6__1_/left_grid_pin_25_ cby_6__1_/left_grid_pin_26_ cby_6__1_/left_grid_pin_27_
+ cby_6__1_/left_grid_pin_28_ cby_6__1_/left_grid_pin_29_ cby_6__1_/left_grid_pin_30_
+ cby_6__1_/left_grid_pin_31_ cby_6__1_/prog_clk_0_N_out sb_6__0_/prog_clk_0_N_in
+ cby_6__1_/prog_clk_0_W_in cby_6__1_/prog_clk_2_N_out cby_6__1_/prog_clk_2_S_in cby_6__1_/prog_clk_2_S_out
+ cby_6__1_/prog_clk_3_N_out cby_6__1_/prog_clk_3_S_in cby_6__1_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_8__5_ cbx_8__4_/SC_OUT_TOP grid_clb_8__5_/SC_OUT_BOT cbx_8__5_/SC_IN_BOT
+ cby_7__5_/Test_en_E_out grid_clb_8__5_/Test_en_E_out cby_7__5_/Test_en_E_out grid_clb_8__5_/Test_en_W_out
+ VGND VPWR cbx_8__4_/REGIN_FEEDTHROUGH grid_clb_8__5_/bottom_width_0_height_0__pin_51_
+ cby_7__5_/ccff_tail cby_8__5_/ccff_head cbx_8__5_/clk_1_S_out cbx_8__5_/clk_1_S_out
+ cby_8__5_/prog_clk_0_W_in cbx_8__5_/prog_clk_1_S_out grid_clb_8__5_/prog_clk_0_N_out
+ cbx_8__5_/prog_clk_1_S_out cbx_8__4_/prog_clk_0_N_in grid_clb_8__5_/prog_clk_0_W_out
+ cby_8__5_/left_grid_pin_16_ cby_8__5_/left_grid_pin_17_ cby_8__5_/left_grid_pin_18_
+ cby_8__5_/left_grid_pin_19_ cby_8__5_/left_grid_pin_20_ cby_8__5_/left_grid_pin_21_
+ cby_8__5_/left_grid_pin_22_ cby_8__5_/left_grid_pin_23_ cby_8__5_/left_grid_pin_24_
+ cby_8__5_/left_grid_pin_25_ cby_8__5_/left_grid_pin_26_ cby_8__5_/left_grid_pin_27_
+ cby_8__5_/left_grid_pin_28_ cby_8__5_/left_grid_pin_29_ cby_8__5_/left_grid_pin_30_
+ cby_8__5_/left_grid_pin_31_ sb_8__4_/top_left_grid_pin_42_ sb_8__5_/bottom_left_grid_pin_42_
+ sb_8__4_/top_left_grid_pin_43_ sb_8__5_/bottom_left_grid_pin_43_ sb_8__4_/top_left_grid_pin_44_
+ sb_8__5_/bottom_left_grid_pin_44_ sb_8__4_/top_left_grid_pin_45_ sb_8__5_/bottom_left_grid_pin_45_
+ sb_8__4_/top_left_grid_pin_46_ sb_8__5_/bottom_left_grid_pin_46_ sb_8__4_/top_left_grid_pin_47_
+ sb_8__5_/bottom_left_grid_pin_47_ sb_8__4_/top_left_grid_pin_48_ sb_8__5_/bottom_left_grid_pin_48_
+ sb_8__4_/top_left_grid_pin_49_ sb_8__5_/bottom_left_grid_pin_49_ cbx_8__5_/bottom_grid_pin_0_
+ cbx_8__5_/bottom_grid_pin_10_ cbx_8__5_/bottom_grid_pin_11_ cbx_8__5_/bottom_grid_pin_12_
+ cbx_8__5_/bottom_grid_pin_13_ cbx_8__5_/bottom_grid_pin_14_ cbx_8__5_/bottom_grid_pin_15_
+ cbx_8__5_/bottom_grid_pin_1_ cbx_8__5_/bottom_grid_pin_2_ cbx_8__5_/REGOUT_FEEDTHROUGH
+ grid_clb_8__5_/top_width_0_height_0__pin_33_ sb_8__5_/left_bottom_grid_pin_34_ sb_7__5_/right_bottom_grid_pin_34_
+ sb_8__5_/left_bottom_grid_pin_35_ sb_7__5_/right_bottom_grid_pin_35_ sb_8__5_/left_bottom_grid_pin_36_
+ sb_7__5_/right_bottom_grid_pin_36_ sb_8__5_/left_bottom_grid_pin_37_ sb_7__5_/right_bottom_grid_pin_37_
+ sb_8__5_/left_bottom_grid_pin_38_ sb_7__5_/right_bottom_grid_pin_38_ sb_8__5_/left_bottom_grid_pin_39_
+ sb_7__5_/right_bottom_grid_pin_39_ cbx_8__5_/bottom_grid_pin_3_ sb_8__5_/left_bottom_grid_pin_40_
+ sb_7__5_/right_bottom_grid_pin_40_ sb_8__5_/left_bottom_grid_pin_41_ sb_7__5_/right_bottom_grid_pin_41_
+ cbx_8__5_/bottom_grid_pin_4_ cbx_8__5_/bottom_grid_pin_5_ cbx_8__5_/bottom_grid_pin_6_
+ cbx_8__5_/bottom_grid_pin_7_ cbx_8__5_/bottom_grid_pin_8_ cbx_8__5_/bottom_grid_pin_9_
+ grid_clb
Xcbx_6__2_ cbx_6__2_/REGIN_FEEDTHROUGH cbx_6__2_/REGOUT_FEEDTHROUGH cbx_6__2_/SC_IN_BOT
+ cbx_6__2_/SC_IN_TOP cbx_6__2_/SC_OUT_BOT cbx_6__2_/SC_OUT_TOP VGND VPWR cbx_6__2_/bottom_grid_pin_0_
+ cbx_6__2_/bottom_grid_pin_10_ cbx_6__2_/bottom_grid_pin_11_ cbx_6__2_/bottom_grid_pin_12_
+ cbx_6__2_/bottom_grid_pin_13_ cbx_6__2_/bottom_grid_pin_14_ cbx_6__2_/bottom_grid_pin_15_
+ cbx_6__2_/bottom_grid_pin_1_ cbx_6__2_/bottom_grid_pin_2_ cbx_6__2_/bottom_grid_pin_3_
+ cbx_6__2_/bottom_grid_pin_4_ cbx_6__2_/bottom_grid_pin_5_ cbx_6__2_/bottom_grid_pin_6_
+ cbx_6__2_/bottom_grid_pin_7_ cbx_6__2_/bottom_grid_pin_8_ cbx_6__2_/bottom_grid_pin_9_
+ sb_6__2_/ccff_tail sb_5__2_/ccff_head cbx_6__2_/chanx_left_in[0] cbx_6__2_/chanx_left_in[10]
+ cbx_6__2_/chanx_left_in[11] cbx_6__2_/chanx_left_in[12] cbx_6__2_/chanx_left_in[13]
+ cbx_6__2_/chanx_left_in[14] cbx_6__2_/chanx_left_in[15] cbx_6__2_/chanx_left_in[16]
+ cbx_6__2_/chanx_left_in[17] cbx_6__2_/chanx_left_in[18] cbx_6__2_/chanx_left_in[19]
+ cbx_6__2_/chanx_left_in[1] cbx_6__2_/chanx_left_in[2] cbx_6__2_/chanx_left_in[3]
+ cbx_6__2_/chanx_left_in[4] cbx_6__2_/chanx_left_in[5] cbx_6__2_/chanx_left_in[6]
+ cbx_6__2_/chanx_left_in[7] cbx_6__2_/chanx_left_in[8] cbx_6__2_/chanx_left_in[9]
+ sb_5__2_/chanx_right_in[0] sb_5__2_/chanx_right_in[10] sb_5__2_/chanx_right_in[11]
+ sb_5__2_/chanx_right_in[12] sb_5__2_/chanx_right_in[13] sb_5__2_/chanx_right_in[14]
+ sb_5__2_/chanx_right_in[15] sb_5__2_/chanx_right_in[16] sb_5__2_/chanx_right_in[17]
+ sb_5__2_/chanx_right_in[18] sb_5__2_/chanx_right_in[19] sb_5__2_/chanx_right_in[1]
+ sb_5__2_/chanx_right_in[2] sb_5__2_/chanx_right_in[3] sb_5__2_/chanx_right_in[4]
+ sb_5__2_/chanx_right_in[5] sb_5__2_/chanx_right_in[6] sb_5__2_/chanx_right_in[7]
+ sb_5__2_/chanx_right_in[8] sb_5__2_/chanx_right_in[9] sb_6__2_/chanx_left_out[0]
+ sb_6__2_/chanx_left_out[10] sb_6__2_/chanx_left_out[11] sb_6__2_/chanx_left_out[12]
+ sb_6__2_/chanx_left_out[13] sb_6__2_/chanx_left_out[14] sb_6__2_/chanx_left_out[15]
+ sb_6__2_/chanx_left_out[16] sb_6__2_/chanx_left_out[17] sb_6__2_/chanx_left_out[18]
+ sb_6__2_/chanx_left_out[19] sb_6__2_/chanx_left_out[1] sb_6__2_/chanx_left_out[2]
+ sb_6__2_/chanx_left_out[3] sb_6__2_/chanx_left_out[4] sb_6__2_/chanx_left_out[5]
+ sb_6__2_/chanx_left_out[6] sb_6__2_/chanx_left_out[7] sb_6__2_/chanx_left_out[8]
+ sb_6__2_/chanx_left_out[9] sb_6__2_/chanx_left_in[0] sb_6__2_/chanx_left_in[10]
+ sb_6__2_/chanx_left_in[11] sb_6__2_/chanx_left_in[12] sb_6__2_/chanx_left_in[13]
+ sb_6__2_/chanx_left_in[14] sb_6__2_/chanx_left_in[15] sb_6__2_/chanx_left_in[16]
+ sb_6__2_/chanx_left_in[17] sb_6__2_/chanx_left_in[18] sb_6__2_/chanx_left_in[19]
+ sb_6__2_/chanx_left_in[1] sb_6__2_/chanx_left_in[2] sb_6__2_/chanx_left_in[3] sb_6__2_/chanx_left_in[4]
+ sb_6__2_/chanx_left_in[5] sb_6__2_/chanx_left_in[6] sb_6__2_/chanx_left_in[7] sb_6__2_/chanx_left_in[8]
+ sb_6__2_/chanx_left_in[9] cbx_6__2_/clk_1_N_out cbx_6__2_/clk_1_S_out cbx_6__2_/clk_1_W_in
+ cbx_6__2_/clk_2_E_out sb_6__2_/clk_2_W_out sb_5__2_/clk_2_N_in cbx_6__2_/clk_3_E_out
+ cbx_6__2_/clk_3_W_in cbx_6__2_/clk_3_W_out cbx_6__2_/prog_clk_0_N_in cbx_6__2_/prog_clk_0_W_out
+ cbx_6__2_/prog_clk_1_N_out cbx_6__2_/prog_clk_1_S_out cbx_6__2_/prog_clk_1_W_in
+ cbx_6__2_/prog_clk_2_E_out sb_6__2_/prog_clk_2_W_out sb_5__2_/prog_clk_2_N_in cbx_6__2_/prog_clk_3_E_out
+ cbx_6__2_/prog_clk_3_W_in cbx_6__2_/prog_clk_3_W_out cbx_1__1_
Xsb_6__7_ sb_6__7_/Test_en_N_out sb_6__7_/Test_en_S_in VGND VPWR sb_6__7_/bottom_left_grid_pin_42_
+ sb_6__7_/bottom_left_grid_pin_43_ sb_6__7_/bottom_left_grid_pin_44_ sb_6__7_/bottom_left_grid_pin_45_
+ sb_6__7_/bottom_left_grid_pin_46_ sb_6__7_/bottom_left_grid_pin_47_ sb_6__7_/bottom_left_grid_pin_48_
+ sb_6__7_/bottom_left_grid_pin_49_ sb_6__7_/ccff_head sb_6__7_/ccff_tail sb_6__7_/chanx_left_in[0]
+ sb_6__7_/chanx_left_in[10] sb_6__7_/chanx_left_in[11] sb_6__7_/chanx_left_in[12]
+ sb_6__7_/chanx_left_in[13] sb_6__7_/chanx_left_in[14] sb_6__7_/chanx_left_in[15]
+ sb_6__7_/chanx_left_in[16] sb_6__7_/chanx_left_in[17] sb_6__7_/chanx_left_in[18]
+ sb_6__7_/chanx_left_in[19] sb_6__7_/chanx_left_in[1] sb_6__7_/chanx_left_in[2] sb_6__7_/chanx_left_in[3]
+ sb_6__7_/chanx_left_in[4] sb_6__7_/chanx_left_in[5] sb_6__7_/chanx_left_in[6] sb_6__7_/chanx_left_in[7]
+ sb_6__7_/chanx_left_in[8] sb_6__7_/chanx_left_in[9] sb_6__7_/chanx_left_out[0] sb_6__7_/chanx_left_out[10]
+ sb_6__7_/chanx_left_out[11] sb_6__7_/chanx_left_out[12] sb_6__7_/chanx_left_out[13]
+ sb_6__7_/chanx_left_out[14] sb_6__7_/chanx_left_out[15] sb_6__7_/chanx_left_out[16]
+ sb_6__7_/chanx_left_out[17] sb_6__7_/chanx_left_out[18] sb_6__7_/chanx_left_out[19]
+ sb_6__7_/chanx_left_out[1] sb_6__7_/chanx_left_out[2] sb_6__7_/chanx_left_out[3]
+ sb_6__7_/chanx_left_out[4] sb_6__7_/chanx_left_out[5] sb_6__7_/chanx_left_out[6]
+ sb_6__7_/chanx_left_out[7] sb_6__7_/chanx_left_out[8] sb_6__7_/chanx_left_out[9]
+ sb_6__7_/chanx_right_in[0] sb_6__7_/chanx_right_in[10] sb_6__7_/chanx_right_in[11]
+ sb_6__7_/chanx_right_in[12] sb_6__7_/chanx_right_in[13] sb_6__7_/chanx_right_in[14]
+ sb_6__7_/chanx_right_in[15] sb_6__7_/chanx_right_in[16] sb_6__7_/chanx_right_in[17]
+ sb_6__7_/chanx_right_in[18] sb_6__7_/chanx_right_in[19] sb_6__7_/chanx_right_in[1]
+ sb_6__7_/chanx_right_in[2] sb_6__7_/chanx_right_in[3] sb_6__7_/chanx_right_in[4]
+ sb_6__7_/chanx_right_in[5] sb_6__7_/chanx_right_in[6] sb_6__7_/chanx_right_in[7]
+ sb_6__7_/chanx_right_in[8] sb_6__7_/chanx_right_in[9] cbx_7__7_/chanx_left_in[0]
+ cbx_7__7_/chanx_left_in[10] cbx_7__7_/chanx_left_in[11] cbx_7__7_/chanx_left_in[12]
+ cbx_7__7_/chanx_left_in[13] cbx_7__7_/chanx_left_in[14] cbx_7__7_/chanx_left_in[15]
+ cbx_7__7_/chanx_left_in[16] cbx_7__7_/chanx_left_in[17] cbx_7__7_/chanx_left_in[18]
+ cbx_7__7_/chanx_left_in[19] cbx_7__7_/chanx_left_in[1] cbx_7__7_/chanx_left_in[2]
+ cbx_7__7_/chanx_left_in[3] cbx_7__7_/chanx_left_in[4] cbx_7__7_/chanx_left_in[5]
+ cbx_7__7_/chanx_left_in[6] cbx_7__7_/chanx_left_in[7] cbx_7__7_/chanx_left_in[8]
+ cbx_7__7_/chanx_left_in[9] cby_6__7_/chany_top_out[0] cby_6__7_/chany_top_out[10]
+ cby_6__7_/chany_top_out[11] cby_6__7_/chany_top_out[12] cby_6__7_/chany_top_out[13]
+ cby_6__7_/chany_top_out[14] cby_6__7_/chany_top_out[15] cby_6__7_/chany_top_out[16]
+ cby_6__7_/chany_top_out[17] cby_6__7_/chany_top_out[18] cby_6__7_/chany_top_out[19]
+ cby_6__7_/chany_top_out[1] cby_6__7_/chany_top_out[2] cby_6__7_/chany_top_out[3]
+ cby_6__7_/chany_top_out[4] cby_6__7_/chany_top_out[5] cby_6__7_/chany_top_out[6]
+ cby_6__7_/chany_top_out[7] cby_6__7_/chany_top_out[8] cby_6__7_/chany_top_out[9]
+ cby_6__7_/chany_top_in[0] cby_6__7_/chany_top_in[10] cby_6__7_/chany_top_in[11]
+ cby_6__7_/chany_top_in[12] cby_6__7_/chany_top_in[13] cby_6__7_/chany_top_in[14]
+ cby_6__7_/chany_top_in[15] cby_6__7_/chany_top_in[16] cby_6__7_/chany_top_in[17]
+ cby_6__7_/chany_top_in[18] cby_6__7_/chany_top_in[19] cby_6__7_/chany_top_in[1]
+ cby_6__7_/chany_top_in[2] cby_6__7_/chany_top_in[3] cby_6__7_/chany_top_in[4] cby_6__7_/chany_top_in[5]
+ cby_6__7_/chany_top_in[6] cby_6__7_/chany_top_in[7] cby_6__7_/chany_top_in[8] cby_6__7_/chany_top_in[9]
+ sb_6__7_/chany_top_in[0] sb_6__7_/chany_top_in[10] sb_6__7_/chany_top_in[11] sb_6__7_/chany_top_in[12]
+ sb_6__7_/chany_top_in[13] sb_6__7_/chany_top_in[14] sb_6__7_/chany_top_in[15] sb_6__7_/chany_top_in[16]
+ sb_6__7_/chany_top_in[17] sb_6__7_/chany_top_in[18] sb_6__7_/chany_top_in[19] sb_6__7_/chany_top_in[1]
+ sb_6__7_/chany_top_in[2] sb_6__7_/chany_top_in[3] sb_6__7_/chany_top_in[4] sb_6__7_/chany_top_in[5]
+ sb_6__7_/chany_top_in[6] sb_6__7_/chany_top_in[7] sb_6__7_/chany_top_in[8] sb_6__7_/chany_top_in[9]
+ sb_6__7_/chany_top_out[0] sb_6__7_/chany_top_out[10] sb_6__7_/chany_top_out[11]
+ sb_6__7_/chany_top_out[12] sb_6__7_/chany_top_out[13] sb_6__7_/chany_top_out[14]
+ sb_6__7_/chany_top_out[15] sb_6__7_/chany_top_out[16] sb_6__7_/chany_top_out[17]
+ sb_6__7_/chany_top_out[18] sb_6__7_/chany_top_out[19] sb_6__7_/chany_top_out[1]
+ sb_6__7_/chany_top_out[2] sb_6__7_/chany_top_out[3] sb_6__7_/chany_top_out[4] sb_6__7_/chany_top_out[5]
+ sb_6__7_/chany_top_out[6] sb_6__7_/chany_top_out[7] sb_6__7_/chany_top_out[8] sb_6__7_/chany_top_out[9]
+ sb_6__7_/clk_1_E_out sb_6__7_/clk_1_N_in sb_6__7_/clk_1_W_out sb_6__7_/clk_2_E_out
+ sb_6__7_/clk_2_N_in sb_6__7_/clk_2_N_out sb_6__7_/clk_2_S_out sb_6__7_/clk_2_W_out
+ sb_6__7_/clk_3_E_out sb_6__7_/clk_3_N_in sb_6__7_/clk_3_N_out sb_6__7_/clk_3_S_out
+ sb_6__7_/clk_3_W_out sb_6__7_/left_bottom_grid_pin_34_ sb_6__7_/left_bottom_grid_pin_35_
+ sb_6__7_/left_bottom_grid_pin_36_ sb_6__7_/left_bottom_grid_pin_37_ sb_6__7_/left_bottom_grid_pin_38_
+ sb_6__7_/left_bottom_grid_pin_39_ sb_6__7_/left_bottom_grid_pin_40_ sb_6__7_/left_bottom_grid_pin_41_
+ sb_6__7_/prog_clk_0_N_in sb_6__7_/prog_clk_1_E_out sb_6__7_/prog_clk_1_N_in sb_6__7_/prog_clk_1_W_out
+ sb_6__7_/prog_clk_2_E_out sb_6__7_/prog_clk_2_N_in sb_6__7_/prog_clk_2_N_out sb_6__7_/prog_clk_2_S_out
+ sb_6__7_/prog_clk_2_W_out sb_6__7_/prog_clk_3_E_out sb_6__7_/prog_clk_3_N_in sb_6__7_/prog_clk_3_N_out
+ sb_6__7_/prog_clk_3_S_out sb_6__7_/prog_clk_3_W_out sb_6__7_/right_bottom_grid_pin_34_
+ sb_6__7_/right_bottom_grid_pin_35_ sb_6__7_/right_bottom_grid_pin_36_ sb_6__7_/right_bottom_grid_pin_37_
+ sb_6__7_/right_bottom_grid_pin_38_ sb_6__7_/right_bottom_grid_pin_39_ sb_6__7_/right_bottom_grid_pin_40_
+ sb_6__7_/right_bottom_grid_pin_41_ sb_6__7_/top_left_grid_pin_42_ sb_6__7_/top_left_grid_pin_43_
+ sb_6__7_/top_left_grid_pin_44_ sb_6__7_/top_left_grid_pin_45_ sb_6__7_/top_left_grid_pin_46_
+ sb_6__7_/top_left_grid_pin_47_ sb_6__7_/top_left_grid_pin_48_ sb_6__7_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_3__4_ sb_3__4_/Test_en_N_out sb_3__4_/Test_en_S_in VGND VPWR sb_3__4_/bottom_left_grid_pin_42_
+ sb_3__4_/bottom_left_grid_pin_43_ sb_3__4_/bottom_left_grid_pin_44_ sb_3__4_/bottom_left_grid_pin_45_
+ sb_3__4_/bottom_left_grid_pin_46_ sb_3__4_/bottom_left_grid_pin_47_ sb_3__4_/bottom_left_grid_pin_48_
+ sb_3__4_/bottom_left_grid_pin_49_ sb_3__4_/ccff_head sb_3__4_/ccff_tail sb_3__4_/chanx_left_in[0]
+ sb_3__4_/chanx_left_in[10] sb_3__4_/chanx_left_in[11] sb_3__4_/chanx_left_in[12]
+ sb_3__4_/chanx_left_in[13] sb_3__4_/chanx_left_in[14] sb_3__4_/chanx_left_in[15]
+ sb_3__4_/chanx_left_in[16] sb_3__4_/chanx_left_in[17] sb_3__4_/chanx_left_in[18]
+ sb_3__4_/chanx_left_in[19] sb_3__4_/chanx_left_in[1] sb_3__4_/chanx_left_in[2] sb_3__4_/chanx_left_in[3]
+ sb_3__4_/chanx_left_in[4] sb_3__4_/chanx_left_in[5] sb_3__4_/chanx_left_in[6] sb_3__4_/chanx_left_in[7]
+ sb_3__4_/chanx_left_in[8] sb_3__4_/chanx_left_in[9] sb_3__4_/chanx_left_out[0] sb_3__4_/chanx_left_out[10]
+ sb_3__4_/chanx_left_out[11] sb_3__4_/chanx_left_out[12] sb_3__4_/chanx_left_out[13]
+ sb_3__4_/chanx_left_out[14] sb_3__4_/chanx_left_out[15] sb_3__4_/chanx_left_out[16]
+ sb_3__4_/chanx_left_out[17] sb_3__4_/chanx_left_out[18] sb_3__4_/chanx_left_out[19]
+ sb_3__4_/chanx_left_out[1] sb_3__4_/chanx_left_out[2] sb_3__4_/chanx_left_out[3]
+ sb_3__4_/chanx_left_out[4] sb_3__4_/chanx_left_out[5] sb_3__4_/chanx_left_out[6]
+ sb_3__4_/chanx_left_out[7] sb_3__4_/chanx_left_out[8] sb_3__4_/chanx_left_out[9]
+ sb_3__4_/chanx_right_in[0] sb_3__4_/chanx_right_in[10] sb_3__4_/chanx_right_in[11]
+ sb_3__4_/chanx_right_in[12] sb_3__4_/chanx_right_in[13] sb_3__4_/chanx_right_in[14]
+ sb_3__4_/chanx_right_in[15] sb_3__4_/chanx_right_in[16] sb_3__4_/chanx_right_in[17]
+ sb_3__4_/chanx_right_in[18] sb_3__4_/chanx_right_in[19] sb_3__4_/chanx_right_in[1]
+ sb_3__4_/chanx_right_in[2] sb_3__4_/chanx_right_in[3] sb_3__4_/chanx_right_in[4]
+ sb_3__4_/chanx_right_in[5] sb_3__4_/chanx_right_in[6] sb_3__4_/chanx_right_in[7]
+ sb_3__4_/chanx_right_in[8] sb_3__4_/chanx_right_in[9] cbx_4__4_/chanx_left_in[0]
+ cbx_4__4_/chanx_left_in[10] cbx_4__4_/chanx_left_in[11] cbx_4__4_/chanx_left_in[12]
+ cbx_4__4_/chanx_left_in[13] cbx_4__4_/chanx_left_in[14] cbx_4__4_/chanx_left_in[15]
+ cbx_4__4_/chanx_left_in[16] cbx_4__4_/chanx_left_in[17] cbx_4__4_/chanx_left_in[18]
+ cbx_4__4_/chanx_left_in[19] cbx_4__4_/chanx_left_in[1] cbx_4__4_/chanx_left_in[2]
+ cbx_4__4_/chanx_left_in[3] cbx_4__4_/chanx_left_in[4] cbx_4__4_/chanx_left_in[5]
+ cbx_4__4_/chanx_left_in[6] cbx_4__4_/chanx_left_in[7] cbx_4__4_/chanx_left_in[8]
+ cbx_4__4_/chanx_left_in[9] cby_3__4_/chany_top_out[0] cby_3__4_/chany_top_out[10]
+ cby_3__4_/chany_top_out[11] cby_3__4_/chany_top_out[12] cby_3__4_/chany_top_out[13]
+ cby_3__4_/chany_top_out[14] cby_3__4_/chany_top_out[15] cby_3__4_/chany_top_out[16]
+ cby_3__4_/chany_top_out[17] cby_3__4_/chany_top_out[18] cby_3__4_/chany_top_out[19]
+ cby_3__4_/chany_top_out[1] cby_3__4_/chany_top_out[2] cby_3__4_/chany_top_out[3]
+ cby_3__4_/chany_top_out[4] cby_3__4_/chany_top_out[5] cby_3__4_/chany_top_out[6]
+ cby_3__4_/chany_top_out[7] cby_3__4_/chany_top_out[8] cby_3__4_/chany_top_out[9]
+ cby_3__4_/chany_top_in[0] cby_3__4_/chany_top_in[10] cby_3__4_/chany_top_in[11]
+ cby_3__4_/chany_top_in[12] cby_3__4_/chany_top_in[13] cby_3__4_/chany_top_in[14]
+ cby_3__4_/chany_top_in[15] cby_3__4_/chany_top_in[16] cby_3__4_/chany_top_in[17]
+ cby_3__4_/chany_top_in[18] cby_3__4_/chany_top_in[19] cby_3__4_/chany_top_in[1]
+ cby_3__4_/chany_top_in[2] cby_3__4_/chany_top_in[3] cby_3__4_/chany_top_in[4] cby_3__4_/chany_top_in[5]
+ cby_3__4_/chany_top_in[6] cby_3__4_/chany_top_in[7] cby_3__4_/chany_top_in[8] cby_3__4_/chany_top_in[9]
+ sb_3__4_/chany_top_in[0] sb_3__4_/chany_top_in[10] sb_3__4_/chany_top_in[11] sb_3__4_/chany_top_in[12]
+ sb_3__4_/chany_top_in[13] sb_3__4_/chany_top_in[14] sb_3__4_/chany_top_in[15] sb_3__4_/chany_top_in[16]
+ sb_3__4_/chany_top_in[17] sb_3__4_/chany_top_in[18] sb_3__4_/chany_top_in[19] sb_3__4_/chany_top_in[1]
+ sb_3__4_/chany_top_in[2] sb_3__4_/chany_top_in[3] sb_3__4_/chany_top_in[4] sb_3__4_/chany_top_in[5]
+ sb_3__4_/chany_top_in[6] sb_3__4_/chany_top_in[7] sb_3__4_/chany_top_in[8] sb_3__4_/chany_top_in[9]
+ sb_3__4_/chany_top_out[0] sb_3__4_/chany_top_out[10] sb_3__4_/chany_top_out[11]
+ sb_3__4_/chany_top_out[12] sb_3__4_/chany_top_out[13] sb_3__4_/chany_top_out[14]
+ sb_3__4_/chany_top_out[15] sb_3__4_/chany_top_out[16] sb_3__4_/chany_top_out[17]
+ sb_3__4_/chany_top_out[18] sb_3__4_/chany_top_out[19] sb_3__4_/chany_top_out[1]
+ sb_3__4_/chany_top_out[2] sb_3__4_/chany_top_out[3] sb_3__4_/chany_top_out[4] sb_3__4_/chany_top_out[5]
+ sb_3__4_/chany_top_out[6] sb_3__4_/chany_top_out[7] sb_3__4_/chany_top_out[8] sb_3__4_/chany_top_out[9]
+ sb_3__4_/clk_1_E_out sb_3__4_/clk_1_N_in sb_3__4_/clk_1_W_out sb_3__4_/clk_2_E_out
+ sb_3__4_/clk_2_N_in sb_3__4_/clk_2_N_out sb_3__4_/clk_2_S_out sb_3__4_/clk_2_W_out
+ sb_3__4_/clk_3_E_out sb_3__4_/clk_3_N_in sb_3__4_/clk_3_N_out sb_3__4_/clk_3_S_out
+ sb_3__4_/clk_3_W_out sb_3__4_/left_bottom_grid_pin_34_ sb_3__4_/left_bottom_grid_pin_35_
+ sb_3__4_/left_bottom_grid_pin_36_ sb_3__4_/left_bottom_grid_pin_37_ sb_3__4_/left_bottom_grid_pin_38_
+ sb_3__4_/left_bottom_grid_pin_39_ sb_3__4_/left_bottom_grid_pin_40_ sb_3__4_/left_bottom_grid_pin_41_
+ sb_3__4_/prog_clk_0_N_in sb_3__4_/prog_clk_1_E_out sb_3__4_/prog_clk_1_N_in sb_3__4_/prog_clk_1_W_out
+ sb_3__4_/prog_clk_2_E_out sb_3__4_/prog_clk_2_N_in sb_3__4_/prog_clk_2_N_out sb_3__4_/prog_clk_2_S_out
+ sb_3__4_/prog_clk_2_W_out sb_3__4_/prog_clk_3_E_out sb_3__4_/prog_clk_3_N_in sb_3__4_/prog_clk_3_N_out
+ sb_3__4_/prog_clk_3_S_out sb_3__4_/prog_clk_3_W_out sb_3__4_/right_bottom_grid_pin_34_
+ sb_3__4_/right_bottom_grid_pin_35_ sb_3__4_/right_bottom_grid_pin_36_ sb_3__4_/right_bottom_grid_pin_37_
+ sb_3__4_/right_bottom_grid_pin_38_ sb_3__4_/right_bottom_grid_pin_39_ sb_3__4_/right_bottom_grid_pin_40_
+ sb_3__4_/right_bottom_grid_pin_41_ sb_3__4_/top_left_grid_pin_42_ sb_3__4_/top_left_grid_pin_43_
+ sb_3__4_/top_left_grid_pin_44_ sb_3__4_/top_left_grid_pin_45_ sb_3__4_/top_left_grid_pin_46_
+ sb_3__4_/top_left_grid_pin_47_ sb_3__4_/top_left_grid_pin_48_ sb_3__4_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_5__2_ cbx_5__2_/SC_OUT_BOT cbx_5__1_/SC_IN_TOP grid_clb_5__2_/SC_OUT_TOP
+ cby_4__2_/Test_en_E_out cby_5__2_/Test_en_W_in cby_4__2_/Test_en_E_out grid_clb_5__2_/Test_en_W_out
+ VGND VPWR cbx_5__1_/REGIN_FEEDTHROUGH grid_clb_5__2_/bottom_width_0_height_0__pin_51_
+ cby_4__2_/ccff_tail cby_5__2_/ccff_head cbx_5__1_/clk_1_N_out cbx_5__1_/clk_1_N_out
+ cby_5__2_/prog_clk_0_W_in cbx_5__1_/prog_clk_1_N_out grid_clb_5__2_/prog_clk_0_N_out
+ cbx_5__1_/prog_clk_1_N_out cbx_5__1_/prog_clk_0_N_in grid_clb_5__2_/prog_clk_0_W_out
+ cby_5__2_/left_grid_pin_16_ cby_5__2_/left_grid_pin_17_ cby_5__2_/left_grid_pin_18_
+ cby_5__2_/left_grid_pin_19_ cby_5__2_/left_grid_pin_20_ cby_5__2_/left_grid_pin_21_
+ cby_5__2_/left_grid_pin_22_ cby_5__2_/left_grid_pin_23_ cby_5__2_/left_grid_pin_24_
+ cby_5__2_/left_grid_pin_25_ cby_5__2_/left_grid_pin_26_ cby_5__2_/left_grid_pin_27_
+ cby_5__2_/left_grid_pin_28_ cby_5__2_/left_grid_pin_29_ cby_5__2_/left_grid_pin_30_
+ cby_5__2_/left_grid_pin_31_ sb_5__1_/top_left_grid_pin_42_ sb_5__2_/bottom_left_grid_pin_42_
+ sb_5__1_/top_left_grid_pin_43_ sb_5__2_/bottom_left_grid_pin_43_ sb_5__1_/top_left_grid_pin_44_
+ sb_5__2_/bottom_left_grid_pin_44_ sb_5__1_/top_left_grid_pin_45_ sb_5__2_/bottom_left_grid_pin_45_
+ sb_5__1_/top_left_grid_pin_46_ sb_5__2_/bottom_left_grid_pin_46_ sb_5__1_/top_left_grid_pin_47_
+ sb_5__2_/bottom_left_grid_pin_47_ sb_5__1_/top_left_grid_pin_48_ sb_5__2_/bottom_left_grid_pin_48_
+ sb_5__1_/top_left_grid_pin_49_ sb_5__2_/bottom_left_grid_pin_49_ cbx_5__2_/bottom_grid_pin_0_
+ cbx_5__2_/bottom_grid_pin_10_ cbx_5__2_/bottom_grid_pin_11_ cbx_5__2_/bottom_grid_pin_12_
+ cbx_5__2_/bottom_grid_pin_13_ cbx_5__2_/bottom_grid_pin_14_ cbx_5__2_/bottom_grid_pin_15_
+ cbx_5__2_/bottom_grid_pin_1_ cbx_5__2_/bottom_grid_pin_2_ cbx_5__2_/REGOUT_FEEDTHROUGH
+ grid_clb_5__2_/top_width_0_height_0__pin_33_ sb_5__2_/left_bottom_grid_pin_34_ sb_4__2_/right_bottom_grid_pin_34_
+ sb_5__2_/left_bottom_grid_pin_35_ sb_4__2_/right_bottom_grid_pin_35_ sb_5__2_/left_bottom_grid_pin_36_
+ sb_4__2_/right_bottom_grid_pin_36_ sb_5__2_/left_bottom_grid_pin_37_ sb_4__2_/right_bottom_grid_pin_37_
+ sb_5__2_/left_bottom_grid_pin_38_ sb_4__2_/right_bottom_grid_pin_38_ sb_5__2_/left_bottom_grid_pin_39_
+ sb_4__2_/right_bottom_grid_pin_39_ cbx_5__2_/bottom_grid_pin_3_ sb_5__2_/left_bottom_grid_pin_40_
+ sb_4__2_/right_bottom_grid_pin_40_ sb_5__2_/left_bottom_grid_pin_41_ sb_4__2_/right_bottom_grid_pin_41_
+ cbx_5__2_/bottom_grid_pin_4_ cbx_5__2_/bottom_grid_pin_5_ cbx_5__2_/bottom_grid_pin_6_
+ cbx_5__2_/bottom_grid_pin_7_ cbx_5__2_/bottom_grid_pin_8_ cbx_5__2_/bottom_grid_pin_9_
+ grid_clb
Xsb_0__1_ VGND VPWR sb_0__1_/bottom_left_grid_pin_1_ sb_0__1_/ccff_head sb_0__1_/ccff_tail
+ sb_0__1_/chanx_right_in[0] sb_0__1_/chanx_right_in[10] sb_0__1_/chanx_right_in[11]
+ sb_0__1_/chanx_right_in[12] sb_0__1_/chanx_right_in[13] sb_0__1_/chanx_right_in[14]
+ sb_0__1_/chanx_right_in[15] sb_0__1_/chanx_right_in[16] sb_0__1_/chanx_right_in[17]
+ sb_0__1_/chanx_right_in[18] sb_0__1_/chanx_right_in[19] sb_0__1_/chanx_right_in[1]
+ sb_0__1_/chanx_right_in[2] sb_0__1_/chanx_right_in[3] sb_0__1_/chanx_right_in[4]
+ sb_0__1_/chanx_right_in[5] sb_0__1_/chanx_right_in[6] sb_0__1_/chanx_right_in[7]
+ sb_0__1_/chanx_right_in[8] sb_0__1_/chanx_right_in[9] cbx_1__1_/chanx_left_in[0]
+ cbx_1__1_/chanx_left_in[10] cbx_1__1_/chanx_left_in[11] cbx_1__1_/chanx_left_in[12]
+ cbx_1__1_/chanx_left_in[13] cbx_1__1_/chanx_left_in[14] cbx_1__1_/chanx_left_in[15]
+ cbx_1__1_/chanx_left_in[16] cbx_1__1_/chanx_left_in[17] cbx_1__1_/chanx_left_in[18]
+ cbx_1__1_/chanx_left_in[19] cbx_1__1_/chanx_left_in[1] cbx_1__1_/chanx_left_in[2]
+ cbx_1__1_/chanx_left_in[3] cbx_1__1_/chanx_left_in[4] cbx_1__1_/chanx_left_in[5]
+ cbx_1__1_/chanx_left_in[6] cbx_1__1_/chanx_left_in[7] cbx_1__1_/chanx_left_in[8]
+ cbx_1__1_/chanx_left_in[9] cby_0__1_/chany_top_out[0] cby_0__1_/chany_top_out[10]
+ cby_0__1_/chany_top_out[11] cby_0__1_/chany_top_out[12] cby_0__1_/chany_top_out[13]
+ cby_0__1_/chany_top_out[14] cby_0__1_/chany_top_out[15] cby_0__1_/chany_top_out[16]
+ cby_0__1_/chany_top_out[17] cby_0__1_/chany_top_out[18] cby_0__1_/chany_top_out[19]
+ cby_0__1_/chany_top_out[1] cby_0__1_/chany_top_out[2] cby_0__1_/chany_top_out[3]
+ cby_0__1_/chany_top_out[4] cby_0__1_/chany_top_out[5] cby_0__1_/chany_top_out[6]
+ cby_0__1_/chany_top_out[7] cby_0__1_/chany_top_out[8] cby_0__1_/chany_top_out[9]
+ cby_0__1_/chany_top_in[0] cby_0__1_/chany_top_in[10] cby_0__1_/chany_top_in[11]
+ cby_0__1_/chany_top_in[12] cby_0__1_/chany_top_in[13] cby_0__1_/chany_top_in[14]
+ cby_0__1_/chany_top_in[15] cby_0__1_/chany_top_in[16] cby_0__1_/chany_top_in[17]
+ cby_0__1_/chany_top_in[18] cby_0__1_/chany_top_in[19] cby_0__1_/chany_top_in[1]
+ cby_0__1_/chany_top_in[2] cby_0__1_/chany_top_in[3] cby_0__1_/chany_top_in[4] cby_0__1_/chany_top_in[5]
+ cby_0__1_/chany_top_in[6] cby_0__1_/chany_top_in[7] cby_0__1_/chany_top_in[8] cby_0__1_/chany_top_in[9]
+ sb_0__1_/chany_top_in[0] sb_0__1_/chany_top_in[10] sb_0__1_/chany_top_in[11] sb_0__1_/chany_top_in[12]
+ sb_0__1_/chany_top_in[13] sb_0__1_/chany_top_in[14] sb_0__1_/chany_top_in[15] sb_0__1_/chany_top_in[16]
+ sb_0__1_/chany_top_in[17] sb_0__1_/chany_top_in[18] sb_0__1_/chany_top_in[19] sb_0__1_/chany_top_in[1]
+ sb_0__1_/chany_top_in[2] sb_0__1_/chany_top_in[3] sb_0__1_/chany_top_in[4] sb_0__1_/chany_top_in[5]
+ sb_0__1_/chany_top_in[6] sb_0__1_/chany_top_in[7] sb_0__1_/chany_top_in[8] sb_0__1_/chany_top_in[9]
+ sb_0__1_/chany_top_out[0] sb_0__1_/chany_top_out[10] sb_0__1_/chany_top_out[11]
+ sb_0__1_/chany_top_out[12] sb_0__1_/chany_top_out[13] sb_0__1_/chany_top_out[14]
+ sb_0__1_/chany_top_out[15] sb_0__1_/chany_top_out[16] sb_0__1_/chany_top_out[17]
+ sb_0__1_/chany_top_out[18] sb_0__1_/chany_top_out[19] sb_0__1_/chany_top_out[1]
+ sb_0__1_/chany_top_out[2] sb_0__1_/chany_top_out[3] sb_0__1_/chany_top_out[4] sb_0__1_/chany_top_out[5]
+ sb_0__1_/chany_top_out[6] sb_0__1_/chany_top_out[7] sb_0__1_/chany_top_out[8] sb_0__1_/chany_top_out[9]
+ sb_0__1_/prog_clk_0_E_in sb_0__1_/right_bottom_grid_pin_34_ sb_0__1_/right_bottom_grid_pin_35_
+ sb_0__1_/right_bottom_grid_pin_36_ sb_0__1_/right_bottom_grid_pin_37_ sb_0__1_/right_bottom_grid_pin_38_
+ sb_0__1_/right_bottom_grid_pin_39_ sb_0__1_/right_bottom_grid_pin_40_ sb_0__1_/right_bottom_grid_pin_41_
+ sb_0__1_/top_left_grid_pin_1_ sb_0__1_
Xcby_2__8_ cby_2__8_/Test_en_W_in cby_2__8_/Test_en_E_out cby_2__8_/Test_en_N_out
+ cby_2__8_/Test_en_W_in cby_2__8_/Test_en_W_in cby_2__8_/Test_en_W_out VGND VPWR
+ cby_2__8_/ccff_head cby_2__8_/ccff_tail sb_2__7_/chany_top_out[0] sb_2__7_/chany_top_out[10]
+ sb_2__7_/chany_top_out[11] sb_2__7_/chany_top_out[12] sb_2__7_/chany_top_out[13]
+ sb_2__7_/chany_top_out[14] sb_2__7_/chany_top_out[15] sb_2__7_/chany_top_out[16]
+ sb_2__7_/chany_top_out[17] sb_2__7_/chany_top_out[18] sb_2__7_/chany_top_out[19]
+ sb_2__7_/chany_top_out[1] sb_2__7_/chany_top_out[2] sb_2__7_/chany_top_out[3] sb_2__7_/chany_top_out[4]
+ sb_2__7_/chany_top_out[5] sb_2__7_/chany_top_out[6] sb_2__7_/chany_top_out[7] sb_2__7_/chany_top_out[8]
+ sb_2__7_/chany_top_out[9] sb_2__7_/chany_top_in[0] sb_2__7_/chany_top_in[10] sb_2__7_/chany_top_in[11]
+ sb_2__7_/chany_top_in[12] sb_2__7_/chany_top_in[13] sb_2__7_/chany_top_in[14] sb_2__7_/chany_top_in[15]
+ sb_2__7_/chany_top_in[16] sb_2__7_/chany_top_in[17] sb_2__7_/chany_top_in[18] sb_2__7_/chany_top_in[19]
+ sb_2__7_/chany_top_in[1] sb_2__7_/chany_top_in[2] sb_2__7_/chany_top_in[3] sb_2__7_/chany_top_in[4]
+ sb_2__7_/chany_top_in[5] sb_2__7_/chany_top_in[6] sb_2__7_/chany_top_in[7] sb_2__7_/chany_top_in[8]
+ sb_2__7_/chany_top_in[9] cby_2__8_/chany_top_in[0] cby_2__8_/chany_top_in[10] cby_2__8_/chany_top_in[11]
+ cby_2__8_/chany_top_in[12] cby_2__8_/chany_top_in[13] cby_2__8_/chany_top_in[14]
+ cby_2__8_/chany_top_in[15] cby_2__8_/chany_top_in[16] cby_2__8_/chany_top_in[17]
+ cby_2__8_/chany_top_in[18] cby_2__8_/chany_top_in[19] cby_2__8_/chany_top_in[1]
+ cby_2__8_/chany_top_in[2] cby_2__8_/chany_top_in[3] cby_2__8_/chany_top_in[4] cby_2__8_/chany_top_in[5]
+ cby_2__8_/chany_top_in[6] cby_2__8_/chany_top_in[7] cby_2__8_/chany_top_in[8] cby_2__8_/chany_top_in[9]
+ cby_2__8_/chany_top_out[0] cby_2__8_/chany_top_out[10] cby_2__8_/chany_top_out[11]
+ cby_2__8_/chany_top_out[12] cby_2__8_/chany_top_out[13] cby_2__8_/chany_top_out[14]
+ cby_2__8_/chany_top_out[15] cby_2__8_/chany_top_out[16] cby_2__8_/chany_top_out[17]
+ cby_2__8_/chany_top_out[18] cby_2__8_/chany_top_out[19] cby_2__8_/chany_top_out[1]
+ cby_2__8_/chany_top_out[2] cby_2__8_/chany_top_out[3] cby_2__8_/chany_top_out[4]
+ cby_2__8_/chany_top_out[5] cby_2__8_/chany_top_out[6] cby_2__8_/chany_top_out[7]
+ cby_2__8_/chany_top_out[8] cby_2__8_/chany_top_out[9] cby_2__8_/clk_2_N_out cby_2__8_/clk_2_S_in
+ cby_2__8_/clk_2_S_out cby_2__8_/clk_3_N_out cby_2__8_/clk_3_S_in cby_2__8_/clk_3_S_out
+ cby_2__8_/left_grid_pin_16_ cby_2__8_/left_grid_pin_17_ cby_2__8_/left_grid_pin_18_
+ cby_2__8_/left_grid_pin_19_ cby_2__8_/left_grid_pin_20_ cby_2__8_/left_grid_pin_21_
+ cby_2__8_/left_grid_pin_22_ cby_2__8_/left_grid_pin_23_ cby_2__8_/left_grid_pin_24_
+ cby_2__8_/left_grid_pin_25_ cby_2__8_/left_grid_pin_26_ cby_2__8_/left_grid_pin_27_
+ cby_2__8_/left_grid_pin_28_ cby_2__8_/left_grid_pin_29_ cby_2__8_/left_grid_pin_30_
+ cby_2__8_/left_grid_pin_31_ sb_2__8_/prog_clk_0_S_in sb_2__7_/prog_clk_0_N_in cby_2__8_/prog_clk_0_W_in
+ cby_2__8_/prog_clk_2_N_out cby_2__8_/prog_clk_2_S_in cby_2__8_/prog_clk_2_S_out
+ cby_2__8_/prog_clk_3_N_out cby_2__8_/prog_clk_3_S_in cby_2__8_/prog_clk_3_S_out
+ cby_1__1_
Xsb_6__6_ sb_6__6_/Test_en_N_out sb_6__6_/Test_en_S_in VGND VPWR sb_6__6_/bottom_left_grid_pin_42_
+ sb_6__6_/bottom_left_grid_pin_43_ sb_6__6_/bottom_left_grid_pin_44_ sb_6__6_/bottom_left_grid_pin_45_
+ sb_6__6_/bottom_left_grid_pin_46_ sb_6__6_/bottom_left_grid_pin_47_ sb_6__6_/bottom_left_grid_pin_48_
+ sb_6__6_/bottom_left_grid_pin_49_ sb_6__6_/ccff_head sb_6__6_/ccff_tail sb_6__6_/chanx_left_in[0]
+ sb_6__6_/chanx_left_in[10] sb_6__6_/chanx_left_in[11] sb_6__6_/chanx_left_in[12]
+ sb_6__6_/chanx_left_in[13] sb_6__6_/chanx_left_in[14] sb_6__6_/chanx_left_in[15]
+ sb_6__6_/chanx_left_in[16] sb_6__6_/chanx_left_in[17] sb_6__6_/chanx_left_in[18]
+ sb_6__6_/chanx_left_in[19] sb_6__6_/chanx_left_in[1] sb_6__6_/chanx_left_in[2] sb_6__6_/chanx_left_in[3]
+ sb_6__6_/chanx_left_in[4] sb_6__6_/chanx_left_in[5] sb_6__6_/chanx_left_in[6] sb_6__6_/chanx_left_in[7]
+ sb_6__6_/chanx_left_in[8] sb_6__6_/chanx_left_in[9] sb_6__6_/chanx_left_out[0] sb_6__6_/chanx_left_out[10]
+ sb_6__6_/chanx_left_out[11] sb_6__6_/chanx_left_out[12] sb_6__6_/chanx_left_out[13]
+ sb_6__6_/chanx_left_out[14] sb_6__6_/chanx_left_out[15] sb_6__6_/chanx_left_out[16]
+ sb_6__6_/chanx_left_out[17] sb_6__6_/chanx_left_out[18] sb_6__6_/chanx_left_out[19]
+ sb_6__6_/chanx_left_out[1] sb_6__6_/chanx_left_out[2] sb_6__6_/chanx_left_out[3]
+ sb_6__6_/chanx_left_out[4] sb_6__6_/chanx_left_out[5] sb_6__6_/chanx_left_out[6]
+ sb_6__6_/chanx_left_out[7] sb_6__6_/chanx_left_out[8] sb_6__6_/chanx_left_out[9]
+ sb_6__6_/chanx_right_in[0] sb_6__6_/chanx_right_in[10] sb_6__6_/chanx_right_in[11]
+ sb_6__6_/chanx_right_in[12] sb_6__6_/chanx_right_in[13] sb_6__6_/chanx_right_in[14]
+ sb_6__6_/chanx_right_in[15] sb_6__6_/chanx_right_in[16] sb_6__6_/chanx_right_in[17]
+ sb_6__6_/chanx_right_in[18] sb_6__6_/chanx_right_in[19] sb_6__6_/chanx_right_in[1]
+ sb_6__6_/chanx_right_in[2] sb_6__6_/chanx_right_in[3] sb_6__6_/chanx_right_in[4]
+ sb_6__6_/chanx_right_in[5] sb_6__6_/chanx_right_in[6] sb_6__6_/chanx_right_in[7]
+ sb_6__6_/chanx_right_in[8] sb_6__6_/chanx_right_in[9] cbx_7__6_/chanx_left_in[0]
+ cbx_7__6_/chanx_left_in[10] cbx_7__6_/chanx_left_in[11] cbx_7__6_/chanx_left_in[12]
+ cbx_7__6_/chanx_left_in[13] cbx_7__6_/chanx_left_in[14] cbx_7__6_/chanx_left_in[15]
+ cbx_7__6_/chanx_left_in[16] cbx_7__6_/chanx_left_in[17] cbx_7__6_/chanx_left_in[18]
+ cbx_7__6_/chanx_left_in[19] cbx_7__6_/chanx_left_in[1] cbx_7__6_/chanx_left_in[2]
+ cbx_7__6_/chanx_left_in[3] cbx_7__6_/chanx_left_in[4] cbx_7__6_/chanx_left_in[5]
+ cbx_7__6_/chanx_left_in[6] cbx_7__6_/chanx_left_in[7] cbx_7__6_/chanx_left_in[8]
+ cbx_7__6_/chanx_left_in[9] cby_6__6_/chany_top_out[0] cby_6__6_/chany_top_out[10]
+ cby_6__6_/chany_top_out[11] cby_6__6_/chany_top_out[12] cby_6__6_/chany_top_out[13]
+ cby_6__6_/chany_top_out[14] cby_6__6_/chany_top_out[15] cby_6__6_/chany_top_out[16]
+ cby_6__6_/chany_top_out[17] cby_6__6_/chany_top_out[18] cby_6__6_/chany_top_out[19]
+ cby_6__6_/chany_top_out[1] cby_6__6_/chany_top_out[2] cby_6__6_/chany_top_out[3]
+ cby_6__6_/chany_top_out[4] cby_6__6_/chany_top_out[5] cby_6__6_/chany_top_out[6]
+ cby_6__6_/chany_top_out[7] cby_6__6_/chany_top_out[8] cby_6__6_/chany_top_out[9]
+ cby_6__6_/chany_top_in[0] cby_6__6_/chany_top_in[10] cby_6__6_/chany_top_in[11]
+ cby_6__6_/chany_top_in[12] cby_6__6_/chany_top_in[13] cby_6__6_/chany_top_in[14]
+ cby_6__6_/chany_top_in[15] cby_6__6_/chany_top_in[16] cby_6__6_/chany_top_in[17]
+ cby_6__6_/chany_top_in[18] cby_6__6_/chany_top_in[19] cby_6__6_/chany_top_in[1]
+ cby_6__6_/chany_top_in[2] cby_6__6_/chany_top_in[3] cby_6__6_/chany_top_in[4] cby_6__6_/chany_top_in[5]
+ cby_6__6_/chany_top_in[6] cby_6__6_/chany_top_in[7] cby_6__6_/chany_top_in[8] cby_6__6_/chany_top_in[9]
+ sb_6__6_/chany_top_in[0] sb_6__6_/chany_top_in[10] sb_6__6_/chany_top_in[11] sb_6__6_/chany_top_in[12]
+ sb_6__6_/chany_top_in[13] sb_6__6_/chany_top_in[14] sb_6__6_/chany_top_in[15] sb_6__6_/chany_top_in[16]
+ sb_6__6_/chany_top_in[17] sb_6__6_/chany_top_in[18] sb_6__6_/chany_top_in[19] sb_6__6_/chany_top_in[1]
+ sb_6__6_/chany_top_in[2] sb_6__6_/chany_top_in[3] sb_6__6_/chany_top_in[4] sb_6__6_/chany_top_in[5]
+ sb_6__6_/chany_top_in[6] sb_6__6_/chany_top_in[7] sb_6__6_/chany_top_in[8] sb_6__6_/chany_top_in[9]
+ sb_6__6_/chany_top_out[0] sb_6__6_/chany_top_out[10] sb_6__6_/chany_top_out[11]
+ sb_6__6_/chany_top_out[12] sb_6__6_/chany_top_out[13] sb_6__6_/chany_top_out[14]
+ sb_6__6_/chany_top_out[15] sb_6__6_/chany_top_out[16] sb_6__6_/chany_top_out[17]
+ sb_6__6_/chany_top_out[18] sb_6__6_/chany_top_out[19] sb_6__6_/chany_top_out[1]
+ sb_6__6_/chany_top_out[2] sb_6__6_/chany_top_out[3] sb_6__6_/chany_top_out[4] sb_6__6_/chany_top_out[5]
+ sb_6__6_/chany_top_out[6] sb_6__6_/chany_top_out[7] sb_6__6_/chany_top_out[8] sb_6__6_/chany_top_out[9]
+ sb_6__6_/clk_1_E_out sb_6__6_/clk_1_N_in sb_6__6_/clk_1_W_out sb_6__6_/clk_2_E_out
+ sb_6__6_/clk_2_N_in sb_6__6_/clk_2_N_out sb_6__6_/clk_2_S_out sb_6__6_/clk_2_W_out
+ sb_6__6_/clk_3_E_out sb_6__6_/clk_3_N_in sb_6__6_/clk_3_N_out sb_6__6_/clk_3_S_out
+ sb_6__6_/clk_3_W_out sb_6__6_/left_bottom_grid_pin_34_ sb_6__6_/left_bottom_grid_pin_35_
+ sb_6__6_/left_bottom_grid_pin_36_ sb_6__6_/left_bottom_grid_pin_37_ sb_6__6_/left_bottom_grid_pin_38_
+ sb_6__6_/left_bottom_grid_pin_39_ sb_6__6_/left_bottom_grid_pin_40_ sb_6__6_/left_bottom_grid_pin_41_
+ sb_6__6_/prog_clk_0_N_in sb_6__6_/prog_clk_1_E_out sb_6__6_/prog_clk_1_N_in sb_6__6_/prog_clk_1_W_out
+ sb_6__6_/prog_clk_2_E_out sb_6__6_/prog_clk_2_N_in sb_6__6_/prog_clk_2_N_out sb_6__6_/prog_clk_2_S_out
+ sb_6__6_/prog_clk_2_W_out sb_6__6_/prog_clk_3_E_out sb_6__6_/prog_clk_3_N_in sb_6__6_/prog_clk_3_N_out
+ sb_6__6_/prog_clk_3_S_out sb_6__6_/prog_clk_3_W_out sb_6__6_/right_bottom_grid_pin_34_
+ sb_6__6_/right_bottom_grid_pin_35_ sb_6__6_/right_bottom_grid_pin_36_ sb_6__6_/right_bottom_grid_pin_37_
+ sb_6__6_/right_bottom_grid_pin_38_ sb_6__6_/right_bottom_grid_pin_39_ sb_6__6_/right_bottom_grid_pin_40_
+ sb_6__6_/right_bottom_grid_pin_41_ sb_6__6_/top_left_grid_pin_42_ sb_6__6_/top_left_grid_pin_43_
+ sb_6__6_/top_left_grid_pin_44_ sb_6__6_/top_left_grid_pin_45_ sb_6__6_/top_left_grid_pin_46_
+ sb_6__6_/top_left_grid_pin_47_ sb_6__6_/top_left_grid_pin_48_ sb_6__6_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_8__4_ cbx_8__3_/SC_OUT_TOP grid_clb_8__4_/SC_OUT_BOT cbx_8__4_/SC_IN_BOT
+ cby_7__4_/Test_en_E_out grid_clb_8__4_/Test_en_E_out cby_7__4_/Test_en_E_out grid_clb_8__4_/Test_en_W_out
+ VGND VPWR cbx_8__3_/REGIN_FEEDTHROUGH grid_clb_8__4_/bottom_width_0_height_0__pin_51_
+ cby_7__4_/ccff_tail cby_8__4_/ccff_head cbx_8__3_/clk_1_N_out cbx_8__3_/clk_1_N_out
+ cby_8__4_/prog_clk_0_W_in cbx_8__3_/prog_clk_1_N_out grid_clb_8__4_/prog_clk_0_N_out
+ cbx_8__3_/prog_clk_1_N_out cbx_8__3_/prog_clk_0_N_in grid_clb_8__4_/prog_clk_0_W_out
+ cby_8__4_/left_grid_pin_16_ cby_8__4_/left_grid_pin_17_ cby_8__4_/left_grid_pin_18_
+ cby_8__4_/left_grid_pin_19_ cby_8__4_/left_grid_pin_20_ cby_8__4_/left_grid_pin_21_
+ cby_8__4_/left_grid_pin_22_ cby_8__4_/left_grid_pin_23_ cby_8__4_/left_grid_pin_24_
+ cby_8__4_/left_grid_pin_25_ cby_8__4_/left_grid_pin_26_ cby_8__4_/left_grid_pin_27_
+ cby_8__4_/left_grid_pin_28_ cby_8__4_/left_grid_pin_29_ cby_8__4_/left_grid_pin_30_
+ cby_8__4_/left_grid_pin_31_ sb_8__3_/top_left_grid_pin_42_ sb_8__4_/bottom_left_grid_pin_42_
+ sb_8__3_/top_left_grid_pin_43_ sb_8__4_/bottom_left_grid_pin_43_ sb_8__3_/top_left_grid_pin_44_
+ sb_8__4_/bottom_left_grid_pin_44_ sb_8__3_/top_left_grid_pin_45_ sb_8__4_/bottom_left_grid_pin_45_
+ sb_8__3_/top_left_grid_pin_46_ sb_8__4_/bottom_left_grid_pin_46_ sb_8__3_/top_left_grid_pin_47_
+ sb_8__4_/bottom_left_grid_pin_47_ sb_8__3_/top_left_grid_pin_48_ sb_8__4_/bottom_left_grid_pin_48_
+ sb_8__3_/top_left_grid_pin_49_ sb_8__4_/bottom_left_grid_pin_49_ cbx_8__4_/bottom_grid_pin_0_
+ cbx_8__4_/bottom_grid_pin_10_ cbx_8__4_/bottom_grid_pin_11_ cbx_8__4_/bottom_grid_pin_12_
+ cbx_8__4_/bottom_grid_pin_13_ cbx_8__4_/bottom_grid_pin_14_ cbx_8__4_/bottom_grid_pin_15_
+ cbx_8__4_/bottom_grid_pin_1_ cbx_8__4_/bottom_grid_pin_2_ cbx_8__4_/REGOUT_FEEDTHROUGH
+ grid_clb_8__4_/top_width_0_height_0__pin_33_ sb_8__4_/left_bottom_grid_pin_34_ sb_7__4_/right_bottom_grid_pin_34_
+ sb_8__4_/left_bottom_grid_pin_35_ sb_7__4_/right_bottom_grid_pin_35_ sb_8__4_/left_bottom_grid_pin_36_
+ sb_7__4_/right_bottom_grid_pin_36_ sb_8__4_/left_bottom_grid_pin_37_ sb_7__4_/right_bottom_grid_pin_37_
+ sb_8__4_/left_bottom_grid_pin_38_ sb_7__4_/right_bottom_grid_pin_38_ sb_8__4_/left_bottom_grid_pin_39_
+ sb_7__4_/right_bottom_grid_pin_39_ cbx_8__4_/bottom_grid_pin_3_ sb_8__4_/left_bottom_grid_pin_40_
+ sb_7__4_/right_bottom_grid_pin_40_ sb_8__4_/left_bottom_grid_pin_41_ sb_7__4_/right_bottom_grid_pin_41_
+ cbx_8__4_/bottom_grid_pin_4_ cbx_8__4_/bottom_grid_pin_5_ cbx_8__4_/bottom_grid_pin_6_
+ cbx_8__4_/bottom_grid_pin_7_ cbx_8__4_/bottom_grid_pin_8_ cbx_8__4_/bottom_grid_pin_9_
+ grid_clb
Xgrid_clb_5__1_ cbx_5__1_/SC_OUT_BOT cbx_5__0_/SC_IN_TOP grid_clb_5__1_/SC_OUT_TOP
+ cby_4__1_/Test_en_E_out cby_5__1_/Test_en_W_in cby_4__1_/Test_en_E_out grid_clb_5__1_/Test_en_W_out
+ VGND VPWR grid_clb_5__1_/bottom_width_0_height_0__pin_50_ grid_clb_5__1_/bottom_width_0_height_0__pin_51_
+ cby_4__1_/ccff_tail cby_5__1_/ccff_head cbx_5__1_/clk_1_S_out cbx_5__1_/clk_1_S_out
+ cby_5__1_/prog_clk_0_W_in cbx_5__1_/prog_clk_1_S_out grid_clb_5__1_/prog_clk_0_N_out
+ cbx_5__1_/prog_clk_1_S_out cbx_5__0_/prog_clk_0_N_in grid_clb_5__1_/prog_clk_0_W_out
+ cby_5__1_/left_grid_pin_16_ cby_5__1_/left_grid_pin_17_ cby_5__1_/left_grid_pin_18_
+ cby_5__1_/left_grid_pin_19_ cby_5__1_/left_grid_pin_20_ cby_5__1_/left_grid_pin_21_
+ cby_5__1_/left_grid_pin_22_ cby_5__1_/left_grid_pin_23_ cby_5__1_/left_grid_pin_24_
+ cby_5__1_/left_grid_pin_25_ cby_5__1_/left_grid_pin_26_ cby_5__1_/left_grid_pin_27_
+ cby_5__1_/left_grid_pin_28_ cby_5__1_/left_grid_pin_29_ cby_5__1_/left_grid_pin_30_
+ cby_5__1_/left_grid_pin_31_ sb_5__0_/top_left_grid_pin_42_ sb_5__1_/bottom_left_grid_pin_42_
+ sb_5__0_/top_left_grid_pin_43_ sb_5__1_/bottom_left_grid_pin_43_ sb_5__0_/top_left_grid_pin_44_
+ sb_5__1_/bottom_left_grid_pin_44_ sb_5__0_/top_left_grid_pin_45_ sb_5__1_/bottom_left_grid_pin_45_
+ sb_5__0_/top_left_grid_pin_46_ sb_5__1_/bottom_left_grid_pin_46_ sb_5__0_/top_left_grid_pin_47_
+ sb_5__1_/bottom_left_grid_pin_47_ sb_5__0_/top_left_grid_pin_48_ sb_5__1_/bottom_left_grid_pin_48_
+ sb_5__0_/top_left_grid_pin_49_ sb_5__1_/bottom_left_grid_pin_49_ cbx_5__1_/bottom_grid_pin_0_
+ cbx_5__1_/bottom_grid_pin_10_ cbx_5__1_/bottom_grid_pin_11_ cbx_5__1_/bottom_grid_pin_12_
+ cbx_5__1_/bottom_grid_pin_13_ cbx_5__1_/bottom_grid_pin_14_ cbx_5__1_/bottom_grid_pin_15_
+ cbx_5__1_/bottom_grid_pin_1_ cbx_5__1_/bottom_grid_pin_2_ cbx_5__1_/REGOUT_FEEDTHROUGH
+ grid_clb_5__1_/top_width_0_height_0__pin_33_ sb_5__1_/left_bottom_grid_pin_34_ sb_4__1_/right_bottom_grid_pin_34_
+ sb_5__1_/left_bottom_grid_pin_35_ sb_4__1_/right_bottom_grid_pin_35_ sb_5__1_/left_bottom_grid_pin_36_
+ sb_4__1_/right_bottom_grid_pin_36_ sb_5__1_/left_bottom_grid_pin_37_ sb_4__1_/right_bottom_grid_pin_37_
+ sb_5__1_/left_bottom_grid_pin_38_ sb_4__1_/right_bottom_grid_pin_38_ sb_5__1_/left_bottom_grid_pin_39_
+ sb_4__1_/right_bottom_grid_pin_39_ cbx_5__1_/bottom_grid_pin_3_ sb_5__1_/left_bottom_grid_pin_40_
+ sb_4__1_/right_bottom_grid_pin_40_ sb_5__1_/left_bottom_grid_pin_41_ sb_4__1_/right_bottom_grid_pin_41_
+ cbx_5__1_/bottom_grid_pin_4_ cbx_5__1_/bottom_grid_pin_5_ cbx_5__1_/bottom_grid_pin_6_
+ cbx_5__1_/bottom_grid_pin_7_ cbx_5__1_/bottom_grid_pin_8_ cbx_5__1_/bottom_grid_pin_9_
+ grid_clb
Xcbx_6__1_ cbx_6__1_/REGIN_FEEDTHROUGH cbx_6__1_/REGOUT_FEEDTHROUGH cbx_6__1_/SC_IN_BOT
+ cbx_6__1_/SC_IN_TOP cbx_6__1_/SC_OUT_BOT cbx_6__1_/SC_OUT_TOP VGND VPWR cbx_6__1_/bottom_grid_pin_0_
+ cbx_6__1_/bottom_grid_pin_10_ cbx_6__1_/bottom_grid_pin_11_ cbx_6__1_/bottom_grid_pin_12_
+ cbx_6__1_/bottom_grid_pin_13_ cbx_6__1_/bottom_grid_pin_14_ cbx_6__1_/bottom_grid_pin_15_
+ cbx_6__1_/bottom_grid_pin_1_ cbx_6__1_/bottom_grid_pin_2_ cbx_6__1_/bottom_grid_pin_3_
+ cbx_6__1_/bottom_grid_pin_4_ cbx_6__1_/bottom_grid_pin_5_ cbx_6__1_/bottom_grid_pin_6_
+ cbx_6__1_/bottom_grid_pin_7_ cbx_6__1_/bottom_grid_pin_8_ cbx_6__1_/bottom_grid_pin_9_
+ sb_6__1_/ccff_tail sb_5__1_/ccff_head cbx_6__1_/chanx_left_in[0] cbx_6__1_/chanx_left_in[10]
+ cbx_6__1_/chanx_left_in[11] cbx_6__1_/chanx_left_in[12] cbx_6__1_/chanx_left_in[13]
+ cbx_6__1_/chanx_left_in[14] cbx_6__1_/chanx_left_in[15] cbx_6__1_/chanx_left_in[16]
+ cbx_6__1_/chanx_left_in[17] cbx_6__1_/chanx_left_in[18] cbx_6__1_/chanx_left_in[19]
+ cbx_6__1_/chanx_left_in[1] cbx_6__1_/chanx_left_in[2] cbx_6__1_/chanx_left_in[3]
+ cbx_6__1_/chanx_left_in[4] cbx_6__1_/chanx_left_in[5] cbx_6__1_/chanx_left_in[6]
+ cbx_6__1_/chanx_left_in[7] cbx_6__1_/chanx_left_in[8] cbx_6__1_/chanx_left_in[9]
+ sb_5__1_/chanx_right_in[0] sb_5__1_/chanx_right_in[10] sb_5__1_/chanx_right_in[11]
+ sb_5__1_/chanx_right_in[12] sb_5__1_/chanx_right_in[13] sb_5__1_/chanx_right_in[14]
+ sb_5__1_/chanx_right_in[15] sb_5__1_/chanx_right_in[16] sb_5__1_/chanx_right_in[17]
+ sb_5__1_/chanx_right_in[18] sb_5__1_/chanx_right_in[19] sb_5__1_/chanx_right_in[1]
+ sb_5__1_/chanx_right_in[2] sb_5__1_/chanx_right_in[3] sb_5__1_/chanx_right_in[4]
+ sb_5__1_/chanx_right_in[5] sb_5__1_/chanx_right_in[6] sb_5__1_/chanx_right_in[7]
+ sb_5__1_/chanx_right_in[8] sb_5__1_/chanx_right_in[9] sb_6__1_/chanx_left_out[0]
+ sb_6__1_/chanx_left_out[10] sb_6__1_/chanx_left_out[11] sb_6__1_/chanx_left_out[12]
+ sb_6__1_/chanx_left_out[13] sb_6__1_/chanx_left_out[14] sb_6__1_/chanx_left_out[15]
+ sb_6__1_/chanx_left_out[16] sb_6__1_/chanx_left_out[17] sb_6__1_/chanx_left_out[18]
+ sb_6__1_/chanx_left_out[19] sb_6__1_/chanx_left_out[1] sb_6__1_/chanx_left_out[2]
+ sb_6__1_/chanx_left_out[3] sb_6__1_/chanx_left_out[4] sb_6__1_/chanx_left_out[5]
+ sb_6__1_/chanx_left_out[6] sb_6__1_/chanx_left_out[7] sb_6__1_/chanx_left_out[8]
+ sb_6__1_/chanx_left_out[9] sb_6__1_/chanx_left_in[0] sb_6__1_/chanx_left_in[10]
+ sb_6__1_/chanx_left_in[11] sb_6__1_/chanx_left_in[12] sb_6__1_/chanx_left_in[13]
+ sb_6__1_/chanx_left_in[14] sb_6__1_/chanx_left_in[15] sb_6__1_/chanx_left_in[16]
+ sb_6__1_/chanx_left_in[17] sb_6__1_/chanx_left_in[18] sb_6__1_/chanx_left_in[19]
+ sb_6__1_/chanx_left_in[1] sb_6__1_/chanx_left_in[2] sb_6__1_/chanx_left_in[3] sb_6__1_/chanx_left_in[4]
+ sb_6__1_/chanx_left_in[5] sb_6__1_/chanx_left_in[6] sb_6__1_/chanx_left_in[7] sb_6__1_/chanx_left_in[8]
+ sb_6__1_/chanx_left_in[9] cbx_6__1_/clk_1_N_out cbx_6__1_/clk_1_S_out sb_5__1_/clk_1_E_out
+ cbx_6__1_/clk_2_E_out cbx_6__1_/clk_2_W_in cbx_6__1_/clk_2_W_out cbx_6__1_/clk_3_E_out
+ cbx_6__1_/clk_3_W_in cbx_6__1_/clk_3_W_out cbx_6__1_/prog_clk_0_N_in cbx_6__1_/prog_clk_0_W_out
+ cbx_6__1_/prog_clk_1_N_out cbx_6__1_/prog_clk_1_S_out sb_5__1_/prog_clk_1_E_out
+ cbx_6__1_/prog_clk_2_E_out cbx_6__1_/prog_clk_2_W_in cbx_6__1_/prog_clk_2_W_out
+ cbx_6__1_/prog_clk_3_E_out cbx_6__1_/prog_clk_3_W_in cbx_6__1_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_3__3_ sb_3__3_/Test_en_N_out sb_3__3_/Test_en_S_in VGND VPWR sb_3__3_/bottom_left_grid_pin_42_
+ sb_3__3_/bottom_left_grid_pin_43_ sb_3__3_/bottom_left_grid_pin_44_ sb_3__3_/bottom_left_grid_pin_45_
+ sb_3__3_/bottom_left_grid_pin_46_ sb_3__3_/bottom_left_grid_pin_47_ sb_3__3_/bottom_left_grid_pin_48_
+ sb_3__3_/bottom_left_grid_pin_49_ sb_3__3_/ccff_head sb_3__3_/ccff_tail sb_3__3_/chanx_left_in[0]
+ sb_3__3_/chanx_left_in[10] sb_3__3_/chanx_left_in[11] sb_3__3_/chanx_left_in[12]
+ sb_3__3_/chanx_left_in[13] sb_3__3_/chanx_left_in[14] sb_3__3_/chanx_left_in[15]
+ sb_3__3_/chanx_left_in[16] sb_3__3_/chanx_left_in[17] sb_3__3_/chanx_left_in[18]
+ sb_3__3_/chanx_left_in[19] sb_3__3_/chanx_left_in[1] sb_3__3_/chanx_left_in[2] sb_3__3_/chanx_left_in[3]
+ sb_3__3_/chanx_left_in[4] sb_3__3_/chanx_left_in[5] sb_3__3_/chanx_left_in[6] sb_3__3_/chanx_left_in[7]
+ sb_3__3_/chanx_left_in[8] sb_3__3_/chanx_left_in[9] sb_3__3_/chanx_left_out[0] sb_3__3_/chanx_left_out[10]
+ sb_3__3_/chanx_left_out[11] sb_3__3_/chanx_left_out[12] sb_3__3_/chanx_left_out[13]
+ sb_3__3_/chanx_left_out[14] sb_3__3_/chanx_left_out[15] sb_3__3_/chanx_left_out[16]
+ sb_3__3_/chanx_left_out[17] sb_3__3_/chanx_left_out[18] sb_3__3_/chanx_left_out[19]
+ sb_3__3_/chanx_left_out[1] sb_3__3_/chanx_left_out[2] sb_3__3_/chanx_left_out[3]
+ sb_3__3_/chanx_left_out[4] sb_3__3_/chanx_left_out[5] sb_3__3_/chanx_left_out[6]
+ sb_3__3_/chanx_left_out[7] sb_3__3_/chanx_left_out[8] sb_3__3_/chanx_left_out[9]
+ sb_3__3_/chanx_right_in[0] sb_3__3_/chanx_right_in[10] sb_3__3_/chanx_right_in[11]
+ sb_3__3_/chanx_right_in[12] sb_3__3_/chanx_right_in[13] sb_3__3_/chanx_right_in[14]
+ sb_3__3_/chanx_right_in[15] sb_3__3_/chanx_right_in[16] sb_3__3_/chanx_right_in[17]
+ sb_3__3_/chanx_right_in[18] sb_3__3_/chanx_right_in[19] sb_3__3_/chanx_right_in[1]
+ sb_3__3_/chanx_right_in[2] sb_3__3_/chanx_right_in[3] sb_3__3_/chanx_right_in[4]
+ sb_3__3_/chanx_right_in[5] sb_3__3_/chanx_right_in[6] sb_3__3_/chanx_right_in[7]
+ sb_3__3_/chanx_right_in[8] sb_3__3_/chanx_right_in[9] cbx_4__3_/chanx_left_in[0]
+ cbx_4__3_/chanx_left_in[10] cbx_4__3_/chanx_left_in[11] cbx_4__3_/chanx_left_in[12]
+ cbx_4__3_/chanx_left_in[13] cbx_4__3_/chanx_left_in[14] cbx_4__3_/chanx_left_in[15]
+ cbx_4__3_/chanx_left_in[16] cbx_4__3_/chanx_left_in[17] cbx_4__3_/chanx_left_in[18]
+ cbx_4__3_/chanx_left_in[19] cbx_4__3_/chanx_left_in[1] cbx_4__3_/chanx_left_in[2]
+ cbx_4__3_/chanx_left_in[3] cbx_4__3_/chanx_left_in[4] cbx_4__3_/chanx_left_in[5]
+ cbx_4__3_/chanx_left_in[6] cbx_4__3_/chanx_left_in[7] cbx_4__3_/chanx_left_in[8]
+ cbx_4__3_/chanx_left_in[9] cby_3__3_/chany_top_out[0] cby_3__3_/chany_top_out[10]
+ cby_3__3_/chany_top_out[11] cby_3__3_/chany_top_out[12] cby_3__3_/chany_top_out[13]
+ cby_3__3_/chany_top_out[14] cby_3__3_/chany_top_out[15] cby_3__3_/chany_top_out[16]
+ cby_3__3_/chany_top_out[17] cby_3__3_/chany_top_out[18] cby_3__3_/chany_top_out[19]
+ cby_3__3_/chany_top_out[1] cby_3__3_/chany_top_out[2] cby_3__3_/chany_top_out[3]
+ cby_3__3_/chany_top_out[4] cby_3__3_/chany_top_out[5] cby_3__3_/chany_top_out[6]
+ cby_3__3_/chany_top_out[7] cby_3__3_/chany_top_out[8] cby_3__3_/chany_top_out[9]
+ cby_3__3_/chany_top_in[0] cby_3__3_/chany_top_in[10] cby_3__3_/chany_top_in[11]
+ cby_3__3_/chany_top_in[12] cby_3__3_/chany_top_in[13] cby_3__3_/chany_top_in[14]
+ cby_3__3_/chany_top_in[15] cby_3__3_/chany_top_in[16] cby_3__3_/chany_top_in[17]
+ cby_3__3_/chany_top_in[18] cby_3__3_/chany_top_in[19] cby_3__3_/chany_top_in[1]
+ cby_3__3_/chany_top_in[2] cby_3__3_/chany_top_in[3] cby_3__3_/chany_top_in[4] cby_3__3_/chany_top_in[5]
+ cby_3__3_/chany_top_in[6] cby_3__3_/chany_top_in[7] cby_3__3_/chany_top_in[8] cby_3__3_/chany_top_in[9]
+ sb_3__3_/chany_top_in[0] sb_3__3_/chany_top_in[10] sb_3__3_/chany_top_in[11] sb_3__3_/chany_top_in[12]
+ sb_3__3_/chany_top_in[13] sb_3__3_/chany_top_in[14] sb_3__3_/chany_top_in[15] sb_3__3_/chany_top_in[16]
+ sb_3__3_/chany_top_in[17] sb_3__3_/chany_top_in[18] sb_3__3_/chany_top_in[19] sb_3__3_/chany_top_in[1]
+ sb_3__3_/chany_top_in[2] sb_3__3_/chany_top_in[3] sb_3__3_/chany_top_in[4] sb_3__3_/chany_top_in[5]
+ sb_3__3_/chany_top_in[6] sb_3__3_/chany_top_in[7] sb_3__3_/chany_top_in[8] sb_3__3_/chany_top_in[9]
+ sb_3__3_/chany_top_out[0] sb_3__3_/chany_top_out[10] sb_3__3_/chany_top_out[11]
+ sb_3__3_/chany_top_out[12] sb_3__3_/chany_top_out[13] sb_3__3_/chany_top_out[14]
+ sb_3__3_/chany_top_out[15] sb_3__3_/chany_top_out[16] sb_3__3_/chany_top_out[17]
+ sb_3__3_/chany_top_out[18] sb_3__3_/chany_top_out[19] sb_3__3_/chany_top_out[1]
+ sb_3__3_/chany_top_out[2] sb_3__3_/chany_top_out[3] sb_3__3_/chany_top_out[4] sb_3__3_/chany_top_out[5]
+ sb_3__3_/chany_top_out[6] sb_3__3_/chany_top_out[7] sb_3__3_/chany_top_out[8] sb_3__3_/chany_top_out[9]
+ sb_3__3_/clk_1_E_out sb_3__3_/clk_1_N_in sb_3__3_/clk_1_W_out sb_3__3_/clk_2_E_out
+ sb_3__3_/clk_2_N_in sb_3__3_/clk_2_N_out sb_3__3_/clk_2_S_out sb_3__3_/clk_2_W_out
+ sb_3__3_/clk_3_E_out sb_3__3_/clk_3_N_in sb_3__3_/clk_3_N_out sb_3__3_/clk_3_S_out
+ sb_3__3_/clk_3_W_out sb_3__3_/left_bottom_grid_pin_34_ sb_3__3_/left_bottom_grid_pin_35_
+ sb_3__3_/left_bottom_grid_pin_36_ sb_3__3_/left_bottom_grid_pin_37_ sb_3__3_/left_bottom_grid_pin_38_
+ sb_3__3_/left_bottom_grid_pin_39_ sb_3__3_/left_bottom_grid_pin_40_ sb_3__3_/left_bottom_grid_pin_41_
+ sb_3__3_/prog_clk_0_N_in sb_3__3_/prog_clk_1_E_out sb_3__3_/prog_clk_1_N_in sb_3__3_/prog_clk_1_W_out
+ sb_3__3_/prog_clk_2_E_out sb_3__3_/prog_clk_2_N_in sb_3__3_/prog_clk_2_N_out sb_3__3_/prog_clk_2_S_out
+ sb_3__3_/prog_clk_2_W_out sb_3__3_/prog_clk_3_E_out sb_3__3_/prog_clk_3_N_in sb_3__3_/prog_clk_3_N_out
+ sb_3__3_/prog_clk_3_S_out sb_3__3_/prog_clk_3_W_out sb_3__3_/right_bottom_grid_pin_34_
+ sb_3__3_/right_bottom_grid_pin_35_ sb_3__3_/right_bottom_grid_pin_36_ sb_3__3_/right_bottom_grid_pin_37_
+ sb_3__3_/right_bottom_grid_pin_38_ sb_3__3_/right_bottom_grid_pin_39_ sb_3__3_/right_bottom_grid_pin_40_
+ sb_3__3_/right_bottom_grid_pin_41_ sb_3__3_/top_left_grid_pin_42_ sb_3__3_/top_left_grid_pin_43_
+ sb_3__3_/top_left_grid_pin_44_ sb_3__3_/top_left_grid_pin_45_ sb_3__3_/top_left_grid_pin_46_
+ sb_3__3_/top_left_grid_pin_47_ sb_3__3_/top_left_grid_pin_48_ sb_3__3_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_0__0_ VGND VPWR sb_0__0_/ccff_head ccff_tail sb_0__0_/chanx_right_in[0] sb_0__0_/chanx_right_in[10]
+ sb_0__0_/chanx_right_in[11] sb_0__0_/chanx_right_in[12] sb_0__0_/chanx_right_in[13]
+ sb_0__0_/chanx_right_in[14] sb_0__0_/chanx_right_in[15] sb_0__0_/chanx_right_in[16]
+ sb_0__0_/chanx_right_in[17] sb_0__0_/chanx_right_in[18] sb_0__0_/chanx_right_in[19]
+ sb_0__0_/chanx_right_in[1] sb_0__0_/chanx_right_in[2] sb_0__0_/chanx_right_in[3]
+ sb_0__0_/chanx_right_in[4] sb_0__0_/chanx_right_in[5] sb_0__0_/chanx_right_in[6]
+ sb_0__0_/chanx_right_in[7] sb_0__0_/chanx_right_in[8] sb_0__0_/chanx_right_in[9]
+ cbx_1__0_/chanx_left_in[0] cbx_1__0_/chanx_left_in[10] cbx_1__0_/chanx_left_in[11]
+ cbx_1__0_/chanx_left_in[12] cbx_1__0_/chanx_left_in[13] cbx_1__0_/chanx_left_in[14]
+ cbx_1__0_/chanx_left_in[15] cbx_1__0_/chanx_left_in[16] cbx_1__0_/chanx_left_in[17]
+ cbx_1__0_/chanx_left_in[18] cbx_1__0_/chanx_left_in[19] cbx_1__0_/chanx_left_in[1]
+ cbx_1__0_/chanx_left_in[2] cbx_1__0_/chanx_left_in[3] cbx_1__0_/chanx_left_in[4]
+ cbx_1__0_/chanx_left_in[5] cbx_1__0_/chanx_left_in[6] cbx_1__0_/chanx_left_in[7]
+ cbx_1__0_/chanx_left_in[8] cbx_1__0_/chanx_left_in[9] sb_0__0_/chany_top_in[0] sb_0__0_/chany_top_in[10]
+ sb_0__0_/chany_top_in[11] sb_0__0_/chany_top_in[12] sb_0__0_/chany_top_in[13] sb_0__0_/chany_top_in[14]
+ sb_0__0_/chany_top_in[15] sb_0__0_/chany_top_in[16] sb_0__0_/chany_top_in[17] sb_0__0_/chany_top_in[18]
+ sb_0__0_/chany_top_in[19] sb_0__0_/chany_top_in[1] sb_0__0_/chany_top_in[2] sb_0__0_/chany_top_in[3]
+ sb_0__0_/chany_top_in[4] sb_0__0_/chany_top_in[5] sb_0__0_/chany_top_in[6] sb_0__0_/chany_top_in[7]
+ sb_0__0_/chany_top_in[8] sb_0__0_/chany_top_in[9] sb_0__0_/chany_top_out[0] sb_0__0_/chany_top_out[10]
+ sb_0__0_/chany_top_out[11] sb_0__0_/chany_top_out[12] sb_0__0_/chany_top_out[13]
+ sb_0__0_/chany_top_out[14] sb_0__0_/chany_top_out[15] sb_0__0_/chany_top_out[16]
+ sb_0__0_/chany_top_out[17] sb_0__0_/chany_top_out[18] sb_0__0_/chany_top_out[19]
+ sb_0__0_/chany_top_out[1] sb_0__0_/chany_top_out[2] sb_0__0_/chany_top_out[3] sb_0__0_/chany_top_out[4]
+ sb_0__0_/chany_top_out[5] sb_0__0_/chany_top_out[6] sb_0__0_/chany_top_out[7] sb_0__0_/chany_top_out[8]
+ sb_0__0_/chany_top_out[9] sb_0__0_/prog_clk_0_E_in sb_0__0_/right_bottom_grid_pin_11_
+ sb_0__0_/right_bottom_grid_pin_13_ sb_0__0_/right_bottom_grid_pin_15_ sb_0__0_/right_bottom_grid_pin_17_
+ sb_0__0_/right_bottom_grid_pin_1_ sb_0__0_/right_bottom_grid_pin_3_ sb_0__0_/right_bottom_grid_pin_5_
+ sb_0__0_/right_bottom_grid_pin_7_ sb_0__0_/right_bottom_grid_pin_9_ sb_0__0_/top_left_grid_pin_1_
+ sb_0__0_
Xcby_2__7_ cby_2__7_/Test_en_W_in cby_2__7_/Test_en_E_out cby_2__7_/Test_en_N_out
+ cby_2__7_/Test_en_W_in cby_2__7_/Test_en_W_in cby_2__7_/Test_en_W_out VGND VPWR
+ cby_2__7_/ccff_head cby_2__7_/ccff_tail sb_2__6_/chany_top_out[0] sb_2__6_/chany_top_out[10]
+ sb_2__6_/chany_top_out[11] sb_2__6_/chany_top_out[12] sb_2__6_/chany_top_out[13]
+ sb_2__6_/chany_top_out[14] sb_2__6_/chany_top_out[15] sb_2__6_/chany_top_out[16]
+ sb_2__6_/chany_top_out[17] sb_2__6_/chany_top_out[18] sb_2__6_/chany_top_out[19]
+ sb_2__6_/chany_top_out[1] sb_2__6_/chany_top_out[2] sb_2__6_/chany_top_out[3] sb_2__6_/chany_top_out[4]
+ sb_2__6_/chany_top_out[5] sb_2__6_/chany_top_out[6] sb_2__6_/chany_top_out[7] sb_2__6_/chany_top_out[8]
+ sb_2__6_/chany_top_out[9] sb_2__6_/chany_top_in[0] sb_2__6_/chany_top_in[10] sb_2__6_/chany_top_in[11]
+ sb_2__6_/chany_top_in[12] sb_2__6_/chany_top_in[13] sb_2__6_/chany_top_in[14] sb_2__6_/chany_top_in[15]
+ sb_2__6_/chany_top_in[16] sb_2__6_/chany_top_in[17] sb_2__6_/chany_top_in[18] sb_2__6_/chany_top_in[19]
+ sb_2__6_/chany_top_in[1] sb_2__6_/chany_top_in[2] sb_2__6_/chany_top_in[3] sb_2__6_/chany_top_in[4]
+ sb_2__6_/chany_top_in[5] sb_2__6_/chany_top_in[6] sb_2__6_/chany_top_in[7] sb_2__6_/chany_top_in[8]
+ sb_2__6_/chany_top_in[9] cby_2__7_/chany_top_in[0] cby_2__7_/chany_top_in[10] cby_2__7_/chany_top_in[11]
+ cby_2__7_/chany_top_in[12] cby_2__7_/chany_top_in[13] cby_2__7_/chany_top_in[14]
+ cby_2__7_/chany_top_in[15] cby_2__7_/chany_top_in[16] cby_2__7_/chany_top_in[17]
+ cby_2__7_/chany_top_in[18] cby_2__7_/chany_top_in[19] cby_2__7_/chany_top_in[1]
+ cby_2__7_/chany_top_in[2] cby_2__7_/chany_top_in[3] cby_2__7_/chany_top_in[4] cby_2__7_/chany_top_in[5]
+ cby_2__7_/chany_top_in[6] cby_2__7_/chany_top_in[7] cby_2__7_/chany_top_in[8] cby_2__7_/chany_top_in[9]
+ cby_2__7_/chany_top_out[0] cby_2__7_/chany_top_out[10] cby_2__7_/chany_top_out[11]
+ cby_2__7_/chany_top_out[12] cby_2__7_/chany_top_out[13] cby_2__7_/chany_top_out[14]
+ cby_2__7_/chany_top_out[15] cby_2__7_/chany_top_out[16] cby_2__7_/chany_top_out[17]
+ cby_2__7_/chany_top_out[18] cby_2__7_/chany_top_out[19] cby_2__7_/chany_top_out[1]
+ cby_2__7_/chany_top_out[2] cby_2__7_/chany_top_out[3] cby_2__7_/chany_top_out[4]
+ cby_2__7_/chany_top_out[5] cby_2__7_/chany_top_out[6] cby_2__7_/chany_top_out[7]
+ cby_2__7_/chany_top_out[8] cby_2__7_/chany_top_out[9] cby_2__7_/clk_2_N_out cby_2__7_/clk_2_S_in
+ cby_2__7_/clk_2_S_out cby_2__7_/clk_3_N_out cby_2__7_/clk_3_S_in cby_2__7_/clk_3_S_out
+ cby_2__7_/left_grid_pin_16_ cby_2__7_/left_grid_pin_17_ cby_2__7_/left_grid_pin_18_
+ cby_2__7_/left_grid_pin_19_ cby_2__7_/left_grid_pin_20_ cby_2__7_/left_grid_pin_21_
+ cby_2__7_/left_grid_pin_22_ cby_2__7_/left_grid_pin_23_ cby_2__7_/left_grid_pin_24_
+ cby_2__7_/left_grid_pin_25_ cby_2__7_/left_grid_pin_26_ cby_2__7_/left_grid_pin_27_
+ cby_2__7_/left_grid_pin_28_ cby_2__7_/left_grid_pin_29_ cby_2__7_/left_grid_pin_30_
+ cby_2__7_/left_grid_pin_31_ cby_2__7_/prog_clk_0_N_out sb_2__6_/prog_clk_0_N_in
+ cby_2__7_/prog_clk_0_W_in cby_2__7_/prog_clk_2_N_out cby_2__7_/prog_clk_2_S_in cby_2__7_/prog_clk_2_S_out
+ cby_2__7_/prog_clk_3_N_out cby_2__7_/prog_clk_3_S_in cby_2__7_/prog_clk_3_S_out
+ cby_1__1_
Xgrid_clb_8__3_ cbx_8__2_/SC_OUT_TOP grid_clb_8__3_/SC_OUT_BOT cbx_8__3_/SC_IN_BOT
+ cby_7__3_/Test_en_E_out grid_clb_8__3_/Test_en_E_out cby_7__3_/Test_en_E_out grid_clb_8__3_/Test_en_W_out
+ VGND VPWR cbx_8__2_/REGIN_FEEDTHROUGH grid_clb_8__3_/bottom_width_0_height_0__pin_51_
+ cby_7__3_/ccff_tail cby_8__3_/ccff_head cbx_8__3_/clk_1_S_out cbx_8__3_/clk_1_S_out
+ cby_8__3_/prog_clk_0_W_in cbx_8__3_/prog_clk_1_S_out grid_clb_8__3_/prog_clk_0_N_out
+ cbx_8__3_/prog_clk_1_S_out cbx_8__2_/prog_clk_0_N_in grid_clb_8__3_/prog_clk_0_W_out
+ cby_8__3_/left_grid_pin_16_ cby_8__3_/left_grid_pin_17_ cby_8__3_/left_grid_pin_18_
+ cby_8__3_/left_grid_pin_19_ cby_8__3_/left_grid_pin_20_ cby_8__3_/left_grid_pin_21_
+ cby_8__3_/left_grid_pin_22_ cby_8__3_/left_grid_pin_23_ cby_8__3_/left_grid_pin_24_
+ cby_8__3_/left_grid_pin_25_ cby_8__3_/left_grid_pin_26_ cby_8__3_/left_grid_pin_27_
+ cby_8__3_/left_grid_pin_28_ cby_8__3_/left_grid_pin_29_ cby_8__3_/left_grid_pin_30_
+ cby_8__3_/left_grid_pin_31_ sb_8__2_/top_left_grid_pin_42_ sb_8__3_/bottom_left_grid_pin_42_
+ sb_8__2_/top_left_grid_pin_43_ sb_8__3_/bottom_left_grid_pin_43_ sb_8__2_/top_left_grid_pin_44_
+ sb_8__3_/bottom_left_grid_pin_44_ sb_8__2_/top_left_grid_pin_45_ sb_8__3_/bottom_left_grid_pin_45_
+ sb_8__2_/top_left_grid_pin_46_ sb_8__3_/bottom_left_grid_pin_46_ sb_8__2_/top_left_grid_pin_47_
+ sb_8__3_/bottom_left_grid_pin_47_ sb_8__2_/top_left_grid_pin_48_ sb_8__3_/bottom_left_grid_pin_48_
+ sb_8__2_/top_left_grid_pin_49_ sb_8__3_/bottom_left_grid_pin_49_ cbx_8__3_/bottom_grid_pin_0_
+ cbx_8__3_/bottom_grid_pin_10_ cbx_8__3_/bottom_grid_pin_11_ cbx_8__3_/bottom_grid_pin_12_
+ cbx_8__3_/bottom_grid_pin_13_ cbx_8__3_/bottom_grid_pin_14_ cbx_8__3_/bottom_grid_pin_15_
+ cbx_8__3_/bottom_grid_pin_1_ cbx_8__3_/bottom_grid_pin_2_ cbx_8__3_/REGOUT_FEEDTHROUGH
+ grid_clb_8__3_/top_width_0_height_0__pin_33_ sb_8__3_/left_bottom_grid_pin_34_ sb_7__3_/right_bottom_grid_pin_34_
+ sb_8__3_/left_bottom_grid_pin_35_ sb_7__3_/right_bottom_grid_pin_35_ sb_8__3_/left_bottom_grid_pin_36_
+ sb_7__3_/right_bottom_grid_pin_36_ sb_8__3_/left_bottom_grid_pin_37_ sb_7__3_/right_bottom_grid_pin_37_
+ sb_8__3_/left_bottom_grid_pin_38_ sb_7__3_/right_bottom_grid_pin_38_ sb_8__3_/left_bottom_grid_pin_39_
+ sb_7__3_/right_bottom_grid_pin_39_ cbx_8__3_/bottom_grid_pin_3_ sb_8__3_/left_bottom_grid_pin_40_
+ sb_7__3_/right_bottom_grid_pin_40_ sb_8__3_/left_bottom_grid_pin_41_ sb_7__3_/right_bottom_grid_pin_41_
+ cbx_8__3_/bottom_grid_pin_4_ cbx_8__3_/bottom_grid_pin_5_ cbx_8__3_/bottom_grid_pin_6_
+ cbx_8__3_/bottom_grid_pin_7_ cbx_8__3_/bottom_grid_pin_8_ cbx_8__3_/bottom_grid_pin_9_
+ grid_clb
Xcbx_6__0_ IO_ISOL_N sb_5__0_/SC_OUT_TOP cbx_6__0_/SC_IN_TOP cbx_6__0_/SC_OUT_BOT
+ cbx_6__0_/SC_OUT_TOP VGND VPWR cbx_6__0_/bottom_grid_pin_0_ cbx_6__0_/bottom_grid_pin_10_
+ cbx_6__0_/bottom_grid_pin_12_ cbx_6__0_/bottom_grid_pin_14_ cbx_6__0_/bottom_grid_pin_16_
+ cbx_6__0_/bottom_grid_pin_2_ cbx_6__0_/bottom_grid_pin_4_ cbx_6__0_/bottom_grid_pin_6_
+ cbx_6__0_/bottom_grid_pin_8_ sb_6__0_/ccff_tail sb_5__0_/ccff_head cbx_6__0_/chanx_left_in[0]
+ cbx_6__0_/chanx_left_in[10] cbx_6__0_/chanx_left_in[11] cbx_6__0_/chanx_left_in[12]
+ cbx_6__0_/chanx_left_in[13] cbx_6__0_/chanx_left_in[14] cbx_6__0_/chanx_left_in[15]
+ cbx_6__0_/chanx_left_in[16] cbx_6__0_/chanx_left_in[17] cbx_6__0_/chanx_left_in[18]
+ cbx_6__0_/chanx_left_in[19] cbx_6__0_/chanx_left_in[1] cbx_6__0_/chanx_left_in[2]
+ cbx_6__0_/chanx_left_in[3] cbx_6__0_/chanx_left_in[4] cbx_6__0_/chanx_left_in[5]
+ cbx_6__0_/chanx_left_in[6] cbx_6__0_/chanx_left_in[7] cbx_6__0_/chanx_left_in[8]
+ cbx_6__0_/chanx_left_in[9] sb_5__0_/chanx_right_in[0] sb_5__0_/chanx_right_in[10]
+ sb_5__0_/chanx_right_in[11] sb_5__0_/chanx_right_in[12] sb_5__0_/chanx_right_in[13]
+ sb_5__0_/chanx_right_in[14] sb_5__0_/chanx_right_in[15] sb_5__0_/chanx_right_in[16]
+ sb_5__0_/chanx_right_in[17] sb_5__0_/chanx_right_in[18] sb_5__0_/chanx_right_in[19]
+ sb_5__0_/chanx_right_in[1] sb_5__0_/chanx_right_in[2] sb_5__0_/chanx_right_in[3]
+ sb_5__0_/chanx_right_in[4] sb_5__0_/chanx_right_in[5] sb_5__0_/chanx_right_in[6]
+ sb_5__0_/chanx_right_in[7] sb_5__0_/chanx_right_in[8] sb_5__0_/chanx_right_in[9]
+ sb_6__0_/chanx_left_out[0] sb_6__0_/chanx_left_out[10] sb_6__0_/chanx_left_out[11]
+ sb_6__0_/chanx_left_out[12] sb_6__0_/chanx_left_out[13] sb_6__0_/chanx_left_out[14]
+ sb_6__0_/chanx_left_out[15] sb_6__0_/chanx_left_out[16] sb_6__0_/chanx_left_out[17]
+ sb_6__0_/chanx_left_out[18] sb_6__0_/chanx_left_out[19] sb_6__0_/chanx_left_out[1]
+ sb_6__0_/chanx_left_out[2] sb_6__0_/chanx_left_out[3] sb_6__0_/chanx_left_out[4]
+ sb_6__0_/chanx_left_out[5] sb_6__0_/chanx_left_out[6] sb_6__0_/chanx_left_out[7]
+ sb_6__0_/chanx_left_out[8] sb_6__0_/chanx_left_out[9] sb_6__0_/chanx_left_in[0]
+ sb_6__0_/chanx_left_in[10] sb_6__0_/chanx_left_in[11] sb_6__0_/chanx_left_in[12]
+ sb_6__0_/chanx_left_in[13] sb_6__0_/chanx_left_in[14] sb_6__0_/chanx_left_in[15]
+ sb_6__0_/chanx_left_in[16] sb_6__0_/chanx_left_in[17] sb_6__0_/chanx_left_in[18]
+ sb_6__0_/chanx_left_in[19] sb_6__0_/chanx_left_in[1] sb_6__0_/chanx_left_in[2] sb_6__0_/chanx_left_in[3]
+ sb_6__0_/chanx_left_in[4] sb_6__0_/chanx_left_in[5] sb_6__0_/chanx_left_in[6] sb_6__0_/chanx_left_in[7]
+ sb_6__0_/chanx_left_in[8] sb_6__0_/chanx_left_in[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42] cbx_6__0_/prog_clk_0_N_in
+ cbx_6__0_/prog_clk_0_W_out cbx_6__0_/bottom_grid_pin_0_ cbx_6__0_/bottom_grid_pin_10_
+ sb_6__0_/left_bottom_grid_pin_11_ sb_5__0_/right_bottom_grid_pin_11_ cbx_6__0_/bottom_grid_pin_12_
+ sb_6__0_/left_bottom_grid_pin_13_ sb_5__0_/right_bottom_grid_pin_13_ cbx_6__0_/bottom_grid_pin_14_
+ sb_6__0_/left_bottom_grid_pin_15_ sb_5__0_/right_bottom_grid_pin_15_ cbx_6__0_/bottom_grid_pin_16_
+ sb_6__0_/left_bottom_grid_pin_17_ sb_5__0_/right_bottom_grid_pin_17_ sb_6__0_/left_bottom_grid_pin_1_
+ sb_5__0_/right_bottom_grid_pin_1_ cbx_6__0_/bottom_grid_pin_2_ sb_6__0_/left_bottom_grid_pin_3_
+ sb_5__0_/right_bottom_grid_pin_3_ cbx_6__0_/bottom_grid_pin_4_ sb_6__0_/left_bottom_grid_pin_5_
+ sb_5__0_/right_bottom_grid_pin_5_ cbx_6__0_/bottom_grid_pin_6_ sb_6__0_/left_bottom_grid_pin_7_
+ sb_5__0_/right_bottom_grid_pin_7_ cbx_6__0_/bottom_grid_pin_8_ sb_6__0_/left_bottom_grid_pin_9_
+ sb_5__0_/right_bottom_grid_pin_9_ cbx_1__0_
Xcbx_2__8_ IO_ISOL_N cbx_2__8_/SC_IN_BOT cbx_2__8_/SC_IN_TOP cbx_2__8_/SC_OUT_BOT
+ sb_2__8_/SC_IN_BOT VGND VPWR cbx_2__8_/bottom_grid_pin_0_ cbx_2__8_/bottom_grid_pin_10_
+ cbx_2__8_/bottom_grid_pin_11_ cbx_2__8_/bottom_grid_pin_12_ cbx_2__8_/bottom_grid_pin_13_
+ cbx_2__8_/bottom_grid_pin_14_ cbx_2__8_/bottom_grid_pin_15_ cbx_2__8_/bottom_grid_pin_1_
+ cbx_2__8_/bottom_grid_pin_2_ cbx_2__8_/bottom_grid_pin_3_ cbx_2__8_/bottom_grid_pin_4_
+ cbx_2__8_/bottom_grid_pin_5_ cbx_2__8_/bottom_grid_pin_6_ cbx_2__8_/bottom_grid_pin_7_
+ cbx_2__8_/bottom_grid_pin_8_ cbx_2__8_/bottom_grid_pin_9_ cbx_2__8_/top_grid_pin_0_
+ sb_2__8_/left_top_grid_pin_1_ sb_1__8_/right_top_grid_pin_1_ sb_2__8_/ccff_tail
+ sb_1__8_/ccff_head cbx_2__8_/chanx_left_in[0] cbx_2__8_/chanx_left_in[10] cbx_2__8_/chanx_left_in[11]
+ cbx_2__8_/chanx_left_in[12] cbx_2__8_/chanx_left_in[13] cbx_2__8_/chanx_left_in[14]
+ cbx_2__8_/chanx_left_in[15] cbx_2__8_/chanx_left_in[16] cbx_2__8_/chanx_left_in[17]
+ cbx_2__8_/chanx_left_in[18] cbx_2__8_/chanx_left_in[19] cbx_2__8_/chanx_left_in[1]
+ cbx_2__8_/chanx_left_in[2] cbx_2__8_/chanx_left_in[3] cbx_2__8_/chanx_left_in[4]
+ cbx_2__8_/chanx_left_in[5] cbx_2__8_/chanx_left_in[6] cbx_2__8_/chanx_left_in[7]
+ cbx_2__8_/chanx_left_in[8] cbx_2__8_/chanx_left_in[9] sb_1__8_/chanx_right_in[0]
+ sb_1__8_/chanx_right_in[10] sb_1__8_/chanx_right_in[11] sb_1__8_/chanx_right_in[12]
+ sb_1__8_/chanx_right_in[13] sb_1__8_/chanx_right_in[14] sb_1__8_/chanx_right_in[15]
+ sb_1__8_/chanx_right_in[16] sb_1__8_/chanx_right_in[17] sb_1__8_/chanx_right_in[18]
+ sb_1__8_/chanx_right_in[19] sb_1__8_/chanx_right_in[1] sb_1__8_/chanx_right_in[2]
+ sb_1__8_/chanx_right_in[3] sb_1__8_/chanx_right_in[4] sb_1__8_/chanx_right_in[5]
+ sb_1__8_/chanx_right_in[6] sb_1__8_/chanx_right_in[7] sb_1__8_/chanx_right_in[8]
+ sb_1__8_/chanx_right_in[9] sb_2__8_/chanx_left_out[0] sb_2__8_/chanx_left_out[10]
+ sb_2__8_/chanx_left_out[11] sb_2__8_/chanx_left_out[12] sb_2__8_/chanx_left_out[13]
+ sb_2__8_/chanx_left_out[14] sb_2__8_/chanx_left_out[15] sb_2__8_/chanx_left_out[16]
+ sb_2__8_/chanx_left_out[17] sb_2__8_/chanx_left_out[18] sb_2__8_/chanx_left_out[19]
+ sb_2__8_/chanx_left_out[1] sb_2__8_/chanx_left_out[2] sb_2__8_/chanx_left_out[3]
+ sb_2__8_/chanx_left_out[4] sb_2__8_/chanx_left_out[5] sb_2__8_/chanx_left_out[6]
+ sb_2__8_/chanx_left_out[7] sb_2__8_/chanx_left_out[8] sb_2__8_/chanx_left_out[9]
+ sb_2__8_/chanx_left_in[0] sb_2__8_/chanx_left_in[10] sb_2__8_/chanx_left_in[11]
+ sb_2__8_/chanx_left_in[12] sb_2__8_/chanx_left_in[13] sb_2__8_/chanx_left_in[14]
+ sb_2__8_/chanx_left_in[15] sb_2__8_/chanx_left_in[16] sb_2__8_/chanx_left_in[17]
+ sb_2__8_/chanx_left_in[18] sb_2__8_/chanx_left_in[19] sb_2__8_/chanx_left_in[1]
+ sb_2__8_/chanx_left_in[2] sb_2__8_/chanx_left_in[3] sb_2__8_/chanx_left_in[4] sb_2__8_/chanx_left_in[5]
+ sb_2__8_/chanx_left_in[6] sb_2__8_/chanx_left_in[7] sb_2__8_/chanx_left_in[8] sb_2__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
+ cbx_2__8_/prog_clk_0_S_in cbx_2__8_/prog_clk_0_W_out cbx_2__8_/top_grid_pin_0_ cbx_1__2_
Xgrid_clb_1__8_ cbx_1__8_/SC_OUT_BOT cbx_1__7_/SC_IN_TOP grid_clb_1__8_/SC_OUT_TOP
+ cby_1__8_/Test_en_W_out grid_clb_1__8_/Test_en_E_out cby_1__8_/Test_en_W_out grid_clb_1__8_/Test_en_W_out
+ VGND VPWR cbx_1__7_/REGIN_FEEDTHROUGH grid_clb_1__8_/bottom_width_0_height_0__pin_51_
+ cby_0__8_/ccff_tail cby_1__8_/ccff_head cbx_1__7_/clk_1_N_out cbx_1__7_/clk_1_N_out
+ cby_1__8_/prog_clk_0_W_in cbx_1__7_/prog_clk_1_N_out cbx_1__8_/prog_clk_0_S_in cbx_1__7_/prog_clk_1_N_out
+ cbx_1__7_/prog_clk_0_N_in cby_0__8_/prog_clk_0_E_in cby_1__8_/left_grid_pin_16_
+ cby_1__8_/left_grid_pin_17_ cby_1__8_/left_grid_pin_18_ cby_1__8_/left_grid_pin_19_
+ cby_1__8_/left_grid_pin_20_ cby_1__8_/left_grid_pin_21_ cby_1__8_/left_grid_pin_22_
+ cby_1__8_/left_grid_pin_23_ cby_1__8_/left_grid_pin_24_ cby_1__8_/left_grid_pin_25_
+ cby_1__8_/left_grid_pin_26_ cby_1__8_/left_grid_pin_27_ cby_1__8_/left_grid_pin_28_
+ cby_1__8_/left_grid_pin_29_ cby_1__8_/left_grid_pin_30_ cby_1__8_/left_grid_pin_31_
+ sb_1__7_/top_left_grid_pin_42_ sb_1__8_/bottom_left_grid_pin_42_ sb_1__7_/top_left_grid_pin_43_
+ sb_1__8_/bottom_left_grid_pin_43_ sb_1__7_/top_left_grid_pin_44_ sb_1__8_/bottom_left_grid_pin_44_
+ sb_1__7_/top_left_grid_pin_45_ sb_1__8_/bottom_left_grid_pin_45_ sb_1__7_/top_left_grid_pin_46_
+ sb_1__8_/bottom_left_grid_pin_46_ sb_1__7_/top_left_grid_pin_47_ sb_1__8_/bottom_left_grid_pin_47_
+ sb_1__7_/top_left_grid_pin_48_ sb_1__8_/bottom_left_grid_pin_48_ sb_1__7_/top_left_grid_pin_49_
+ sb_1__8_/bottom_left_grid_pin_49_ cbx_1__8_/bottom_grid_pin_0_ cbx_1__8_/bottom_grid_pin_10_
+ cbx_1__8_/bottom_grid_pin_11_ cbx_1__8_/bottom_grid_pin_12_ cbx_1__8_/bottom_grid_pin_13_
+ cbx_1__8_/bottom_grid_pin_14_ cbx_1__8_/bottom_grid_pin_15_ cbx_1__8_/bottom_grid_pin_1_
+ cbx_1__8_/bottom_grid_pin_2_ tie_array/x[0] grid_clb_1__8_/top_width_0_height_0__pin_33_
+ sb_1__8_/left_bottom_grid_pin_34_ sb_0__8_/right_bottom_grid_pin_34_ sb_1__8_/left_bottom_grid_pin_35_
+ sb_0__8_/right_bottom_grid_pin_35_ sb_1__8_/left_bottom_grid_pin_36_ sb_0__8_/right_bottom_grid_pin_36_
+ sb_1__8_/left_bottom_grid_pin_37_ sb_0__8_/right_bottom_grid_pin_37_ sb_1__8_/left_bottom_grid_pin_38_
+ sb_0__8_/right_bottom_grid_pin_38_ sb_1__8_/left_bottom_grid_pin_39_ sb_0__8_/right_bottom_grid_pin_39_
+ cbx_1__8_/bottom_grid_pin_3_ sb_1__8_/left_bottom_grid_pin_40_ sb_0__8_/right_bottom_grid_pin_40_
+ sb_1__8_/left_bottom_grid_pin_41_ sb_0__8_/right_bottom_grid_pin_41_ cbx_1__8_/bottom_grid_pin_4_
+ cbx_1__8_/bottom_grid_pin_5_ cbx_1__8_/bottom_grid_pin_6_ cbx_1__8_/bottom_grid_pin_7_
+ cbx_1__8_/bottom_grid_pin_8_ cbx_1__8_/bottom_grid_pin_9_ grid_clb
Xsb_6__5_ sb_6__5_/Test_en_N_out sb_6__5_/Test_en_S_in VGND VPWR sb_6__5_/bottom_left_grid_pin_42_
+ sb_6__5_/bottom_left_grid_pin_43_ sb_6__5_/bottom_left_grid_pin_44_ sb_6__5_/bottom_left_grid_pin_45_
+ sb_6__5_/bottom_left_grid_pin_46_ sb_6__5_/bottom_left_grid_pin_47_ sb_6__5_/bottom_left_grid_pin_48_
+ sb_6__5_/bottom_left_grid_pin_49_ sb_6__5_/ccff_head sb_6__5_/ccff_tail sb_6__5_/chanx_left_in[0]
+ sb_6__5_/chanx_left_in[10] sb_6__5_/chanx_left_in[11] sb_6__5_/chanx_left_in[12]
+ sb_6__5_/chanx_left_in[13] sb_6__5_/chanx_left_in[14] sb_6__5_/chanx_left_in[15]
+ sb_6__5_/chanx_left_in[16] sb_6__5_/chanx_left_in[17] sb_6__5_/chanx_left_in[18]
+ sb_6__5_/chanx_left_in[19] sb_6__5_/chanx_left_in[1] sb_6__5_/chanx_left_in[2] sb_6__5_/chanx_left_in[3]
+ sb_6__5_/chanx_left_in[4] sb_6__5_/chanx_left_in[5] sb_6__5_/chanx_left_in[6] sb_6__5_/chanx_left_in[7]
+ sb_6__5_/chanx_left_in[8] sb_6__5_/chanx_left_in[9] sb_6__5_/chanx_left_out[0] sb_6__5_/chanx_left_out[10]
+ sb_6__5_/chanx_left_out[11] sb_6__5_/chanx_left_out[12] sb_6__5_/chanx_left_out[13]
+ sb_6__5_/chanx_left_out[14] sb_6__5_/chanx_left_out[15] sb_6__5_/chanx_left_out[16]
+ sb_6__5_/chanx_left_out[17] sb_6__5_/chanx_left_out[18] sb_6__5_/chanx_left_out[19]
+ sb_6__5_/chanx_left_out[1] sb_6__5_/chanx_left_out[2] sb_6__5_/chanx_left_out[3]
+ sb_6__5_/chanx_left_out[4] sb_6__5_/chanx_left_out[5] sb_6__5_/chanx_left_out[6]
+ sb_6__5_/chanx_left_out[7] sb_6__5_/chanx_left_out[8] sb_6__5_/chanx_left_out[9]
+ sb_6__5_/chanx_right_in[0] sb_6__5_/chanx_right_in[10] sb_6__5_/chanx_right_in[11]
+ sb_6__5_/chanx_right_in[12] sb_6__5_/chanx_right_in[13] sb_6__5_/chanx_right_in[14]
+ sb_6__5_/chanx_right_in[15] sb_6__5_/chanx_right_in[16] sb_6__5_/chanx_right_in[17]
+ sb_6__5_/chanx_right_in[18] sb_6__5_/chanx_right_in[19] sb_6__5_/chanx_right_in[1]
+ sb_6__5_/chanx_right_in[2] sb_6__5_/chanx_right_in[3] sb_6__5_/chanx_right_in[4]
+ sb_6__5_/chanx_right_in[5] sb_6__5_/chanx_right_in[6] sb_6__5_/chanx_right_in[7]
+ sb_6__5_/chanx_right_in[8] sb_6__5_/chanx_right_in[9] cbx_7__5_/chanx_left_in[0]
+ cbx_7__5_/chanx_left_in[10] cbx_7__5_/chanx_left_in[11] cbx_7__5_/chanx_left_in[12]
+ cbx_7__5_/chanx_left_in[13] cbx_7__5_/chanx_left_in[14] cbx_7__5_/chanx_left_in[15]
+ cbx_7__5_/chanx_left_in[16] cbx_7__5_/chanx_left_in[17] cbx_7__5_/chanx_left_in[18]
+ cbx_7__5_/chanx_left_in[19] cbx_7__5_/chanx_left_in[1] cbx_7__5_/chanx_left_in[2]
+ cbx_7__5_/chanx_left_in[3] cbx_7__5_/chanx_left_in[4] cbx_7__5_/chanx_left_in[5]
+ cbx_7__5_/chanx_left_in[6] cbx_7__5_/chanx_left_in[7] cbx_7__5_/chanx_left_in[8]
+ cbx_7__5_/chanx_left_in[9] cby_6__5_/chany_top_out[0] cby_6__5_/chany_top_out[10]
+ cby_6__5_/chany_top_out[11] cby_6__5_/chany_top_out[12] cby_6__5_/chany_top_out[13]
+ cby_6__5_/chany_top_out[14] cby_6__5_/chany_top_out[15] cby_6__5_/chany_top_out[16]
+ cby_6__5_/chany_top_out[17] cby_6__5_/chany_top_out[18] cby_6__5_/chany_top_out[19]
+ cby_6__5_/chany_top_out[1] cby_6__5_/chany_top_out[2] cby_6__5_/chany_top_out[3]
+ cby_6__5_/chany_top_out[4] cby_6__5_/chany_top_out[5] cby_6__5_/chany_top_out[6]
+ cby_6__5_/chany_top_out[7] cby_6__5_/chany_top_out[8] cby_6__5_/chany_top_out[9]
+ cby_6__5_/chany_top_in[0] cby_6__5_/chany_top_in[10] cby_6__5_/chany_top_in[11]
+ cby_6__5_/chany_top_in[12] cby_6__5_/chany_top_in[13] cby_6__5_/chany_top_in[14]
+ cby_6__5_/chany_top_in[15] cby_6__5_/chany_top_in[16] cby_6__5_/chany_top_in[17]
+ cby_6__5_/chany_top_in[18] cby_6__5_/chany_top_in[19] cby_6__5_/chany_top_in[1]
+ cby_6__5_/chany_top_in[2] cby_6__5_/chany_top_in[3] cby_6__5_/chany_top_in[4] cby_6__5_/chany_top_in[5]
+ cby_6__5_/chany_top_in[6] cby_6__5_/chany_top_in[7] cby_6__5_/chany_top_in[8] cby_6__5_/chany_top_in[9]
+ sb_6__5_/chany_top_in[0] sb_6__5_/chany_top_in[10] sb_6__5_/chany_top_in[11] sb_6__5_/chany_top_in[12]
+ sb_6__5_/chany_top_in[13] sb_6__5_/chany_top_in[14] sb_6__5_/chany_top_in[15] sb_6__5_/chany_top_in[16]
+ sb_6__5_/chany_top_in[17] sb_6__5_/chany_top_in[18] sb_6__5_/chany_top_in[19] sb_6__5_/chany_top_in[1]
+ sb_6__5_/chany_top_in[2] sb_6__5_/chany_top_in[3] sb_6__5_/chany_top_in[4] sb_6__5_/chany_top_in[5]
+ sb_6__5_/chany_top_in[6] sb_6__5_/chany_top_in[7] sb_6__5_/chany_top_in[8] sb_6__5_/chany_top_in[9]
+ sb_6__5_/chany_top_out[0] sb_6__5_/chany_top_out[10] sb_6__5_/chany_top_out[11]
+ sb_6__5_/chany_top_out[12] sb_6__5_/chany_top_out[13] sb_6__5_/chany_top_out[14]
+ sb_6__5_/chany_top_out[15] sb_6__5_/chany_top_out[16] sb_6__5_/chany_top_out[17]
+ sb_6__5_/chany_top_out[18] sb_6__5_/chany_top_out[19] sb_6__5_/chany_top_out[1]
+ sb_6__5_/chany_top_out[2] sb_6__5_/chany_top_out[3] sb_6__5_/chany_top_out[4] sb_6__5_/chany_top_out[5]
+ sb_6__5_/chany_top_out[6] sb_6__5_/chany_top_out[7] sb_6__5_/chany_top_out[8] sb_6__5_/chany_top_out[9]
+ sb_6__5_/clk_1_E_out sb_6__5_/clk_1_N_in sb_6__5_/clk_1_W_out sb_6__5_/clk_2_E_out
+ sb_6__5_/clk_2_N_in sb_6__5_/clk_2_N_out sb_6__5_/clk_2_S_out sb_6__5_/clk_2_W_out
+ sb_6__5_/clk_3_E_out sb_6__5_/clk_3_N_in sb_6__5_/clk_3_N_out sb_6__5_/clk_3_S_out
+ sb_6__5_/clk_3_W_out sb_6__5_/left_bottom_grid_pin_34_ sb_6__5_/left_bottom_grid_pin_35_
+ sb_6__5_/left_bottom_grid_pin_36_ sb_6__5_/left_bottom_grid_pin_37_ sb_6__5_/left_bottom_grid_pin_38_
+ sb_6__5_/left_bottom_grid_pin_39_ sb_6__5_/left_bottom_grid_pin_40_ sb_6__5_/left_bottom_grid_pin_41_
+ sb_6__5_/prog_clk_0_N_in sb_6__5_/prog_clk_1_E_out sb_6__5_/prog_clk_1_N_in sb_6__5_/prog_clk_1_W_out
+ sb_6__5_/prog_clk_2_E_out sb_6__5_/prog_clk_2_N_in sb_6__5_/prog_clk_2_N_out sb_6__5_/prog_clk_2_S_out
+ sb_6__5_/prog_clk_2_W_out sb_6__5_/prog_clk_3_E_out sb_6__5_/prog_clk_3_N_in sb_6__5_/prog_clk_3_N_out
+ sb_6__5_/prog_clk_3_S_out sb_6__5_/prog_clk_3_W_out sb_6__5_/right_bottom_grid_pin_34_
+ sb_6__5_/right_bottom_grid_pin_35_ sb_6__5_/right_bottom_grid_pin_36_ sb_6__5_/right_bottom_grid_pin_37_
+ sb_6__5_/right_bottom_grid_pin_38_ sb_6__5_/right_bottom_grid_pin_39_ sb_6__5_/right_bottom_grid_pin_40_
+ sb_6__5_/right_bottom_grid_pin_41_ sb_6__5_/top_left_grid_pin_42_ sb_6__5_/top_left_grid_pin_43_
+ sb_6__5_/top_left_grid_pin_44_ sb_6__5_/top_left_grid_pin_45_ sb_6__5_/top_left_grid_pin_46_
+ sb_6__5_/top_left_grid_pin_47_ sb_6__5_/top_left_grid_pin_48_ sb_6__5_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_3__2_ sb_3__2_/Test_en_N_out sb_3__2_/Test_en_S_in VGND VPWR sb_3__2_/bottom_left_grid_pin_42_
+ sb_3__2_/bottom_left_grid_pin_43_ sb_3__2_/bottom_left_grid_pin_44_ sb_3__2_/bottom_left_grid_pin_45_
+ sb_3__2_/bottom_left_grid_pin_46_ sb_3__2_/bottom_left_grid_pin_47_ sb_3__2_/bottom_left_grid_pin_48_
+ sb_3__2_/bottom_left_grid_pin_49_ sb_3__2_/ccff_head sb_3__2_/ccff_tail sb_3__2_/chanx_left_in[0]
+ sb_3__2_/chanx_left_in[10] sb_3__2_/chanx_left_in[11] sb_3__2_/chanx_left_in[12]
+ sb_3__2_/chanx_left_in[13] sb_3__2_/chanx_left_in[14] sb_3__2_/chanx_left_in[15]
+ sb_3__2_/chanx_left_in[16] sb_3__2_/chanx_left_in[17] sb_3__2_/chanx_left_in[18]
+ sb_3__2_/chanx_left_in[19] sb_3__2_/chanx_left_in[1] sb_3__2_/chanx_left_in[2] sb_3__2_/chanx_left_in[3]
+ sb_3__2_/chanx_left_in[4] sb_3__2_/chanx_left_in[5] sb_3__2_/chanx_left_in[6] sb_3__2_/chanx_left_in[7]
+ sb_3__2_/chanx_left_in[8] sb_3__2_/chanx_left_in[9] sb_3__2_/chanx_left_out[0] sb_3__2_/chanx_left_out[10]
+ sb_3__2_/chanx_left_out[11] sb_3__2_/chanx_left_out[12] sb_3__2_/chanx_left_out[13]
+ sb_3__2_/chanx_left_out[14] sb_3__2_/chanx_left_out[15] sb_3__2_/chanx_left_out[16]
+ sb_3__2_/chanx_left_out[17] sb_3__2_/chanx_left_out[18] sb_3__2_/chanx_left_out[19]
+ sb_3__2_/chanx_left_out[1] sb_3__2_/chanx_left_out[2] sb_3__2_/chanx_left_out[3]
+ sb_3__2_/chanx_left_out[4] sb_3__2_/chanx_left_out[5] sb_3__2_/chanx_left_out[6]
+ sb_3__2_/chanx_left_out[7] sb_3__2_/chanx_left_out[8] sb_3__2_/chanx_left_out[9]
+ sb_3__2_/chanx_right_in[0] sb_3__2_/chanx_right_in[10] sb_3__2_/chanx_right_in[11]
+ sb_3__2_/chanx_right_in[12] sb_3__2_/chanx_right_in[13] sb_3__2_/chanx_right_in[14]
+ sb_3__2_/chanx_right_in[15] sb_3__2_/chanx_right_in[16] sb_3__2_/chanx_right_in[17]
+ sb_3__2_/chanx_right_in[18] sb_3__2_/chanx_right_in[19] sb_3__2_/chanx_right_in[1]
+ sb_3__2_/chanx_right_in[2] sb_3__2_/chanx_right_in[3] sb_3__2_/chanx_right_in[4]
+ sb_3__2_/chanx_right_in[5] sb_3__2_/chanx_right_in[6] sb_3__2_/chanx_right_in[7]
+ sb_3__2_/chanx_right_in[8] sb_3__2_/chanx_right_in[9] cbx_4__2_/chanx_left_in[0]
+ cbx_4__2_/chanx_left_in[10] cbx_4__2_/chanx_left_in[11] cbx_4__2_/chanx_left_in[12]
+ cbx_4__2_/chanx_left_in[13] cbx_4__2_/chanx_left_in[14] cbx_4__2_/chanx_left_in[15]
+ cbx_4__2_/chanx_left_in[16] cbx_4__2_/chanx_left_in[17] cbx_4__2_/chanx_left_in[18]
+ cbx_4__2_/chanx_left_in[19] cbx_4__2_/chanx_left_in[1] cbx_4__2_/chanx_left_in[2]
+ cbx_4__2_/chanx_left_in[3] cbx_4__2_/chanx_left_in[4] cbx_4__2_/chanx_left_in[5]
+ cbx_4__2_/chanx_left_in[6] cbx_4__2_/chanx_left_in[7] cbx_4__2_/chanx_left_in[8]
+ cbx_4__2_/chanx_left_in[9] cby_3__2_/chany_top_out[0] cby_3__2_/chany_top_out[10]
+ cby_3__2_/chany_top_out[11] cby_3__2_/chany_top_out[12] cby_3__2_/chany_top_out[13]
+ cby_3__2_/chany_top_out[14] cby_3__2_/chany_top_out[15] cby_3__2_/chany_top_out[16]
+ cby_3__2_/chany_top_out[17] cby_3__2_/chany_top_out[18] cby_3__2_/chany_top_out[19]
+ cby_3__2_/chany_top_out[1] cby_3__2_/chany_top_out[2] cby_3__2_/chany_top_out[3]
+ cby_3__2_/chany_top_out[4] cby_3__2_/chany_top_out[5] cby_3__2_/chany_top_out[6]
+ cby_3__2_/chany_top_out[7] cby_3__2_/chany_top_out[8] cby_3__2_/chany_top_out[9]
+ cby_3__2_/chany_top_in[0] cby_3__2_/chany_top_in[10] cby_3__2_/chany_top_in[11]
+ cby_3__2_/chany_top_in[12] cby_3__2_/chany_top_in[13] cby_3__2_/chany_top_in[14]
+ cby_3__2_/chany_top_in[15] cby_3__2_/chany_top_in[16] cby_3__2_/chany_top_in[17]
+ cby_3__2_/chany_top_in[18] cby_3__2_/chany_top_in[19] cby_3__2_/chany_top_in[1]
+ cby_3__2_/chany_top_in[2] cby_3__2_/chany_top_in[3] cby_3__2_/chany_top_in[4] cby_3__2_/chany_top_in[5]
+ cby_3__2_/chany_top_in[6] cby_3__2_/chany_top_in[7] cby_3__2_/chany_top_in[8] cby_3__2_/chany_top_in[9]
+ sb_3__2_/chany_top_in[0] sb_3__2_/chany_top_in[10] sb_3__2_/chany_top_in[11] sb_3__2_/chany_top_in[12]
+ sb_3__2_/chany_top_in[13] sb_3__2_/chany_top_in[14] sb_3__2_/chany_top_in[15] sb_3__2_/chany_top_in[16]
+ sb_3__2_/chany_top_in[17] sb_3__2_/chany_top_in[18] sb_3__2_/chany_top_in[19] sb_3__2_/chany_top_in[1]
+ sb_3__2_/chany_top_in[2] sb_3__2_/chany_top_in[3] sb_3__2_/chany_top_in[4] sb_3__2_/chany_top_in[5]
+ sb_3__2_/chany_top_in[6] sb_3__2_/chany_top_in[7] sb_3__2_/chany_top_in[8] sb_3__2_/chany_top_in[9]
+ sb_3__2_/chany_top_out[0] sb_3__2_/chany_top_out[10] sb_3__2_/chany_top_out[11]
+ sb_3__2_/chany_top_out[12] sb_3__2_/chany_top_out[13] sb_3__2_/chany_top_out[14]
+ sb_3__2_/chany_top_out[15] sb_3__2_/chany_top_out[16] sb_3__2_/chany_top_out[17]
+ sb_3__2_/chany_top_out[18] sb_3__2_/chany_top_out[19] sb_3__2_/chany_top_out[1]
+ sb_3__2_/chany_top_out[2] sb_3__2_/chany_top_out[3] sb_3__2_/chany_top_out[4] sb_3__2_/chany_top_out[5]
+ sb_3__2_/chany_top_out[6] sb_3__2_/chany_top_out[7] sb_3__2_/chany_top_out[8] sb_3__2_/chany_top_out[9]
+ sb_3__2_/clk_1_E_out sb_3__2_/clk_1_N_in sb_3__2_/clk_1_W_out sb_3__2_/clk_2_E_out
+ sb_3__2_/clk_2_N_in sb_3__2_/clk_2_N_out sb_3__2_/clk_2_S_out sb_3__2_/clk_2_W_out
+ sb_3__2_/clk_3_E_out sb_3__2_/clk_3_N_in sb_3__2_/clk_3_N_out sb_3__2_/clk_3_S_out
+ sb_3__2_/clk_3_W_out sb_3__2_/left_bottom_grid_pin_34_ sb_3__2_/left_bottom_grid_pin_35_
+ sb_3__2_/left_bottom_grid_pin_36_ sb_3__2_/left_bottom_grid_pin_37_ sb_3__2_/left_bottom_grid_pin_38_
+ sb_3__2_/left_bottom_grid_pin_39_ sb_3__2_/left_bottom_grid_pin_40_ sb_3__2_/left_bottom_grid_pin_41_
+ sb_3__2_/prog_clk_0_N_in sb_3__2_/prog_clk_1_E_out sb_3__2_/prog_clk_1_N_in sb_3__2_/prog_clk_1_W_out
+ sb_3__2_/prog_clk_2_E_out sb_3__2_/prog_clk_2_N_in sb_3__2_/prog_clk_2_N_out sb_3__2_/prog_clk_2_S_out
+ sb_3__2_/prog_clk_2_W_out sb_3__2_/prog_clk_3_E_out sb_3__2_/prog_clk_3_N_in sb_3__2_/prog_clk_3_N_out
+ sb_3__2_/prog_clk_3_S_out sb_3__2_/prog_clk_3_W_out sb_3__2_/right_bottom_grid_pin_34_
+ sb_3__2_/right_bottom_grid_pin_35_ sb_3__2_/right_bottom_grid_pin_36_ sb_3__2_/right_bottom_grid_pin_37_
+ sb_3__2_/right_bottom_grid_pin_38_ sb_3__2_/right_bottom_grid_pin_39_ sb_3__2_/right_bottom_grid_pin_40_
+ sb_3__2_/right_bottom_grid_pin_41_ sb_3__2_/top_left_grid_pin_42_ sb_3__2_/top_left_grid_pin_43_
+ sb_3__2_/top_left_grid_pin_44_ sb_3__2_/top_left_grid_pin_45_ sb_3__2_/top_left_grid_pin_46_
+ sb_3__2_/top_left_grid_pin_47_ sb_3__2_/top_left_grid_pin_48_ sb_3__2_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_2__6_ cby_2__6_/Test_en_W_in cby_2__6_/Test_en_E_out cby_2__6_/Test_en_N_out
+ cby_2__6_/Test_en_W_in cby_2__6_/Test_en_W_in cby_2__6_/Test_en_W_out VGND VPWR
+ cby_2__6_/ccff_head cby_2__6_/ccff_tail sb_2__5_/chany_top_out[0] sb_2__5_/chany_top_out[10]
+ sb_2__5_/chany_top_out[11] sb_2__5_/chany_top_out[12] sb_2__5_/chany_top_out[13]
+ sb_2__5_/chany_top_out[14] sb_2__5_/chany_top_out[15] sb_2__5_/chany_top_out[16]
+ sb_2__5_/chany_top_out[17] sb_2__5_/chany_top_out[18] sb_2__5_/chany_top_out[19]
+ sb_2__5_/chany_top_out[1] sb_2__5_/chany_top_out[2] sb_2__5_/chany_top_out[3] sb_2__5_/chany_top_out[4]
+ sb_2__5_/chany_top_out[5] sb_2__5_/chany_top_out[6] sb_2__5_/chany_top_out[7] sb_2__5_/chany_top_out[8]
+ sb_2__5_/chany_top_out[9] sb_2__5_/chany_top_in[0] sb_2__5_/chany_top_in[10] sb_2__5_/chany_top_in[11]
+ sb_2__5_/chany_top_in[12] sb_2__5_/chany_top_in[13] sb_2__5_/chany_top_in[14] sb_2__5_/chany_top_in[15]
+ sb_2__5_/chany_top_in[16] sb_2__5_/chany_top_in[17] sb_2__5_/chany_top_in[18] sb_2__5_/chany_top_in[19]
+ sb_2__5_/chany_top_in[1] sb_2__5_/chany_top_in[2] sb_2__5_/chany_top_in[3] sb_2__5_/chany_top_in[4]
+ sb_2__5_/chany_top_in[5] sb_2__5_/chany_top_in[6] sb_2__5_/chany_top_in[7] sb_2__5_/chany_top_in[8]
+ sb_2__5_/chany_top_in[9] cby_2__6_/chany_top_in[0] cby_2__6_/chany_top_in[10] cby_2__6_/chany_top_in[11]
+ cby_2__6_/chany_top_in[12] cby_2__6_/chany_top_in[13] cby_2__6_/chany_top_in[14]
+ cby_2__6_/chany_top_in[15] cby_2__6_/chany_top_in[16] cby_2__6_/chany_top_in[17]
+ cby_2__6_/chany_top_in[18] cby_2__6_/chany_top_in[19] cby_2__6_/chany_top_in[1]
+ cby_2__6_/chany_top_in[2] cby_2__6_/chany_top_in[3] cby_2__6_/chany_top_in[4] cby_2__6_/chany_top_in[5]
+ cby_2__6_/chany_top_in[6] cby_2__6_/chany_top_in[7] cby_2__6_/chany_top_in[8] cby_2__6_/chany_top_in[9]
+ cby_2__6_/chany_top_out[0] cby_2__6_/chany_top_out[10] cby_2__6_/chany_top_out[11]
+ cby_2__6_/chany_top_out[12] cby_2__6_/chany_top_out[13] cby_2__6_/chany_top_out[14]
+ cby_2__6_/chany_top_out[15] cby_2__6_/chany_top_out[16] cby_2__6_/chany_top_out[17]
+ cby_2__6_/chany_top_out[18] cby_2__6_/chany_top_out[19] cby_2__6_/chany_top_out[1]
+ cby_2__6_/chany_top_out[2] cby_2__6_/chany_top_out[3] cby_2__6_/chany_top_out[4]
+ cby_2__6_/chany_top_out[5] cby_2__6_/chany_top_out[6] cby_2__6_/chany_top_out[7]
+ cby_2__6_/chany_top_out[8] cby_2__6_/chany_top_out[9] cby_2__6_/clk_2_N_out cby_2__6_/clk_2_S_in
+ cby_2__6_/clk_2_S_out sb_2__6_/clk_2_N_in sb_2__5_/clk_3_N_out cby_2__6_/clk_3_S_out
+ cby_2__6_/left_grid_pin_16_ cby_2__6_/left_grid_pin_17_ cby_2__6_/left_grid_pin_18_
+ cby_2__6_/left_grid_pin_19_ cby_2__6_/left_grid_pin_20_ cby_2__6_/left_grid_pin_21_
+ cby_2__6_/left_grid_pin_22_ cby_2__6_/left_grid_pin_23_ cby_2__6_/left_grid_pin_24_
+ cby_2__6_/left_grid_pin_25_ cby_2__6_/left_grid_pin_26_ cby_2__6_/left_grid_pin_27_
+ cby_2__6_/left_grid_pin_28_ cby_2__6_/left_grid_pin_29_ cby_2__6_/left_grid_pin_30_
+ cby_2__6_/left_grid_pin_31_ cby_2__6_/prog_clk_0_N_out sb_2__5_/prog_clk_0_N_in
+ cby_2__6_/prog_clk_0_W_in cby_2__6_/prog_clk_2_N_out cby_2__6_/prog_clk_2_S_in cby_2__6_/prog_clk_2_S_out
+ sb_2__6_/prog_clk_2_N_in sb_2__5_/prog_clk_3_N_out cby_2__6_/prog_clk_3_S_out cby_1__1_
Xcbx_2__7_ cbx_2__7_/REGIN_FEEDTHROUGH cbx_2__7_/REGOUT_FEEDTHROUGH cbx_2__7_/SC_IN_BOT
+ cbx_2__7_/SC_IN_TOP cbx_2__7_/SC_OUT_BOT cbx_2__7_/SC_OUT_TOP VGND VPWR cbx_2__7_/bottom_grid_pin_0_
+ cbx_2__7_/bottom_grid_pin_10_ cbx_2__7_/bottom_grid_pin_11_ cbx_2__7_/bottom_grid_pin_12_
+ cbx_2__7_/bottom_grid_pin_13_ cbx_2__7_/bottom_grid_pin_14_ cbx_2__7_/bottom_grid_pin_15_
+ cbx_2__7_/bottom_grid_pin_1_ cbx_2__7_/bottom_grid_pin_2_ cbx_2__7_/bottom_grid_pin_3_
+ cbx_2__7_/bottom_grid_pin_4_ cbx_2__7_/bottom_grid_pin_5_ cbx_2__7_/bottom_grid_pin_6_
+ cbx_2__7_/bottom_grid_pin_7_ cbx_2__7_/bottom_grid_pin_8_ cbx_2__7_/bottom_grid_pin_9_
+ sb_2__7_/ccff_tail sb_1__7_/ccff_head cbx_2__7_/chanx_left_in[0] cbx_2__7_/chanx_left_in[10]
+ cbx_2__7_/chanx_left_in[11] cbx_2__7_/chanx_left_in[12] cbx_2__7_/chanx_left_in[13]
+ cbx_2__7_/chanx_left_in[14] cbx_2__7_/chanx_left_in[15] cbx_2__7_/chanx_left_in[16]
+ cbx_2__7_/chanx_left_in[17] cbx_2__7_/chanx_left_in[18] cbx_2__7_/chanx_left_in[19]
+ cbx_2__7_/chanx_left_in[1] cbx_2__7_/chanx_left_in[2] cbx_2__7_/chanx_left_in[3]
+ cbx_2__7_/chanx_left_in[4] cbx_2__7_/chanx_left_in[5] cbx_2__7_/chanx_left_in[6]
+ cbx_2__7_/chanx_left_in[7] cbx_2__7_/chanx_left_in[8] cbx_2__7_/chanx_left_in[9]
+ sb_1__7_/chanx_right_in[0] sb_1__7_/chanx_right_in[10] sb_1__7_/chanx_right_in[11]
+ sb_1__7_/chanx_right_in[12] sb_1__7_/chanx_right_in[13] sb_1__7_/chanx_right_in[14]
+ sb_1__7_/chanx_right_in[15] sb_1__7_/chanx_right_in[16] sb_1__7_/chanx_right_in[17]
+ sb_1__7_/chanx_right_in[18] sb_1__7_/chanx_right_in[19] sb_1__7_/chanx_right_in[1]
+ sb_1__7_/chanx_right_in[2] sb_1__7_/chanx_right_in[3] sb_1__7_/chanx_right_in[4]
+ sb_1__7_/chanx_right_in[5] sb_1__7_/chanx_right_in[6] sb_1__7_/chanx_right_in[7]
+ sb_1__7_/chanx_right_in[8] sb_1__7_/chanx_right_in[9] sb_2__7_/chanx_left_out[0]
+ sb_2__7_/chanx_left_out[10] sb_2__7_/chanx_left_out[11] sb_2__7_/chanx_left_out[12]
+ sb_2__7_/chanx_left_out[13] sb_2__7_/chanx_left_out[14] sb_2__7_/chanx_left_out[15]
+ sb_2__7_/chanx_left_out[16] sb_2__7_/chanx_left_out[17] sb_2__7_/chanx_left_out[18]
+ sb_2__7_/chanx_left_out[19] sb_2__7_/chanx_left_out[1] sb_2__7_/chanx_left_out[2]
+ sb_2__7_/chanx_left_out[3] sb_2__7_/chanx_left_out[4] sb_2__7_/chanx_left_out[5]
+ sb_2__7_/chanx_left_out[6] sb_2__7_/chanx_left_out[7] sb_2__7_/chanx_left_out[8]
+ sb_2__7_/chanx_left_out[9] sb_2__7_/chanx_left_in[0] sb_2__7_/chanx_left_in[10]
+ sb_2__7_/chanx_left_in[11] sb_2__7_/chanx_left_in[12] sb_2__7_/chanx_left_in[13]
+ sb_2__7_/chanx_left_in[14] sb_2__7_/chanx_left_in[15] sb_2__7_/chanx_left_in[16]
+ sb_2__7_/chanx_left_in[17] sb_2__7_/chanx_left_in[18] sb_2__7_/chanx_left_in[19]
+ sb_2__7_/chanx_left_in[1] sb_2__7_/chanx_left_in[2] sb_2__7_/chanx_left_in[3] sb_2__7_/chanx_left_in[4]
+ sb_2__7_/chanx_left_in[5] sb_2__7_/chanx_left_in[6] sb_2__7_/chanx_left_in[7] sb_2__7_/chanx_left_in[8]
+ sb_2__7_/chanx_left_in[9] cbx_2__7_/clk_1_N_out cbx_2__7_/clk_1_S_out sb_1__7_/clk_1_E_out
+ cbx_2__7_/clk_2_E_out cbx_2__7_/clk_2_W_in cbx_2__7_/clk_2_W_out cbx_2__7_/clk_3_E_out
+ cbx_2__7_/clk_3_W_in cbx_2__7_/clk_3_W_out cbx_2__7_/prog_clk_0_N_in cbx_2__7_/prog_clk_0_W_out
+ cbx_2__7_/prog_clk_1_N_out cbx_2__7_/prog_clk_1_S_out sb_1__7_/prog_clk_1_E_out
+ cbx_2__7_/prog_clk_2_E_out cbx_2__7_/prog_clk_2_W_in cbx_2__7_/prog_clk_2_W_out
+ cbx_2__7_/prog_clk_3_E_out cbx_2__7_/prog_clk_3_W_in cbx_2__7_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_6__4_ sb_6__4_/Test_en_N_out sb_6__4_/Test_en_S_in VGND VPWR sb_6__4_/bottom_left_grid_pin_42_
+ sb_6__4_/bottom_left_grid_pin_43_ sb_6__4_/bottom_left_grid_pin_44_ sb_6__4_/bottom_left_grid_pin_45_
+ sb_6__4_/bottom_left_grid_pin_46_ sb_6__4_/bottom_left_grid_pin_47_ sb_6__4_/bottom_left_grid_pin_48_
+ sb_6__4_/bottom_left_grid_pin_49_ sb_6__4_/ccff_head sb_6__4_/ccff_tail sb_6__4_/chanx_left_in[0]
+ sb_6__4_/chanx_left_in[10] sb_6__4_/chanx_left_in[11] sb_6__4_/chanx_left_in[12]
+ sb_6__4_/chanx_left_in[13] sb_6__4_/chanx_left_in[14] sb_6__4_/chanx_left_in[15]
+ sb_6__4_/chanx_left_in[16] sb_6__4_/chanx_left_in[17] sb_6__4_/chanx_left_in[18]
+ sb_6__4_/chanx_left_in[19] sb_6__4_/chanx_left_in[1] sb_6__4_/chanx_left_in[2] sb_6__4_/chanx_left_in[3]
+ sb_6__4_/chanx_left_in[4] sb_6__4_/chanx_left_in[5] sb_6__4_/chanx_left_in[6] sb_6__4_/chanx_left_in[7]
+ sb_6__4_/chanx_left_in[8] sb_6__4_/chanx_left_in[9] sb_6__4_/chanx_left_out[0] sb_6__4_/chanx_left_out[10]
+ sb_6__4_/chanx_left_out[11] sb_6__4_/chanx_left_out[12] sb_6__4_/chanx_left_out[13]
+ sb_6__4_/chanx_left_out[14] sb_6__4_/chanx_left_out[15] sb_6__4_/chanx_left_out[16]
+ sb_6__4_/chanx_left_out[17] sb_6__4_/chanx_left_out[18] sb_6__4_/chanx_left_out[19]
+ sb_6__4_/chanx_left_out[1] sb_6__4_/chanx_left_out[2] sb_6__4_/chanx_left_out[3]
+ sb_6__4_/chanx_left_out[4] sb_6__4_/chanx_left_out[5] sb_6__4_/chanx_left_out[6]
+ sb_6__4_/chanx_left_out[7] sb_6__4_/chanx_left_out[8] sb_6__4_/chanx_left_out[9]
+ sb_6__4_/chanx_right_in[0] sb_6__4_/chanx_right_in[10] sb_6__4_/chanx_right_in[11]
+ sb_6__4_/chanx_right_in[12] sb_6__4_/chanx_right_in[13] sb_6__4_/chanx_right_in[14]
+ sb_6__4_/chanx_right_in[15] sb_6__4_/chanx_right_in[16] sb_6__4_/chanx_right_in[17]
+ sb_6__4_/chanx_right_in[18] sb_6__4_/chanx_right_in[19] sb_6__4_/chanx_right_in[1]
+ sb_6__4_/chanx_right_in[2] sb_6__4_/chanx_right_in[3] sb_6__4_/chanx_right_in[4]
+ sb_6__4_/chanx_right_in[5] sb_6__4_/chanx_right_in[6] sb_6__4_/chanx_right_in[7]
+ sb_6__4_/chanx_right_in[8] sb_6__4_/chanx_right_in[9] cbx_7__4_/chanx_left_in[0]
+ cbx_7__4_/chanx_left_in[10] cbx_7__4_/chanx_left_in[11] cbx_7__4_/chanx_left_in[12]
+ cbx_7__4_/chanx_left_in[13] cbx_7__4_/chanx_left_in[14] cbx_7__4_/chanx_left_in[15]
+ cbx_7__4_/chanx_left_in[16] cbx_7__4_/chanx_left_in[17] cbx_7__4_/chanx_left_in[18]
+ cbx_7__4_/chanx_left_in[19] cbx_7__4_/chanx_left_in[1] cbx_7__4_/chanx_left_in[2]
+ cbx_7__4_/chanx_left_in[3] cbx_7__4_/chanx_left_in[4] cbx_7__4_/chanx_left_in[5]
+ cbx_7__4_/chanx_left_in[6] cbx_7__4_/chanx_left_in[7] cbx_7__4_/chanx_left_in[8]
+ cbx_7__4_/chanx_left_in[9] cby_6__4_/chany_top_out[0] cby_6__4_/chany_top_out[10]
+ cby_6__4_/chany_top_out[11] cby_6__4_/chany_top_out[12] cby_6__4_/chany_top_out[13]
+ cby_6__4_/chany_top_out[14] cby_6__4_/chany_top_out[15] cby_6__4_/chany_top_out[16]
+ cby_6__4_/chany_top_out[17] cby_6__4_/chany_top_out[18] cby_6__4_/chany_top_out[19]
+ cby_6__4_/chany_top_out[1] cby_6__4_/chany_top_out[2] cby_6__4_/chany_top_out[3]
+ cby_6__4_/chany_top_out[4] cby_6__4_/chany_top_out[5] cby_6__4_/chany_top_out[6]
+ cby_6__4_/chany_top_out[7] cby_6__4_/chany_top_out[8] cby_6__4_/chany_top_out[9]
+ cby_6__4_/chany_top_in[0] cby_6__4_/chany_top_in[10] cby_6__4_/chany_top_in[11]
+ cby_6__4_/chany_top_in[12] cby_6__4_/chany_top_in[13] cby_6__4_/chany_top_in[14]
+ cby_6__4_/chany_top_in[15] cby_6__4_/chany_top_in[16] cby_6__4_/chany_top_in[17]
+ cby_6__4_/chany_top_in[18] cby_6__4_/chany_top_in[19] cby_6__4_/chany_top_in[1]
+ cby_6__4_/chany_top_in[2] cby_6__4_/chany_top_in[3] cby_6__4_/chany_top_in[4] cby_6__4_/chany_top_in[5]
+ cby_6__4_/chany_top_in[6] cby_6__4_/chany_top_in[7] cby_6__4_/chany_top_in[8] cby_6__4_/chany_top_in[9]
+ sb_6__4_/chany_top_in[0] sb_6__4_/chany_top_in[10] sb_6__4_/chany_top_in[11] sb_6__4_/chany_top_in[12]
+ sb_6__4_/chany_top_in[13] sb_6__4_/chany_top_in[14] sb_6__4_/chany_top_in[15] sb_6__4_/chany_top_in[16]
+ sb_6__4_/chany_top_in[17] sb_6__4_/chany_top_in[18] sb_6__4_/chany_top_in[19] sb_6__4_/chany_top_in[1]
+ sb_6__4_/chany_top_in[2] sb_6__4_/chany_top_in[3] sb_6__4_/chany_top_in[4] sb_6__4_/chany_top_in[5]
+ sb_6__4_/chany_top_in[6] sb_6__4_/chany_top_in[7] sb_6__4_/chany_top_in[8] sb_6__4_/chany_top_in[9]
+ sb_6__4_/chany_top_out[0] sb_6__4_/chany_top_out[10] sb_6__4_/chany_top_out[11]
+ sb_6__4_/chany_top_out[12] sb_6__4_/chany_top_out[13] sb_6__4_/chany_top_out[14]
+ sb_6__4_/chany_top_out[15] sb_6__4_/chany_top_out[16] sb_6__4_/chany_top_out[17]
+ sb_6__4_/chany_top_out[18] sb_6__4_/chany_top_out[19] sb_6__4_/chany_top_out[1]
+ sb_6__4_/chany_top_out[2] sb_6__4_/chany_top_out[3] sb_6__4_/chany_top_out[4] sb_6__4_/chany_top_out[5]
+ sb_6__4_/chany_top_out[6] sb_6__4_/chany_top_out[7] sb_6__4_/chany_top_out[8] sb_6__4_/chany_top_out[9]
+ sb_6__4_/clk_1_E_out sb_6__4_/clk_1_N_in sb_6__4_/clk_1_W_out sb_6__4_/clk_2_E_out
+ sb_6__4_/clk_2_N_in sb_6__4_/clk_2_N_out sb_6__4_/clk_2_S_out sb_6__4_/clk_2_W_out
+ sb_6__4_/clk_3_E_out sb_6__4_/clk_3_N_in sb_6__4_/clk_3_N_out sb_6__4_/clk_3_S_out
+ sb_6__4_/clk_3_W_out sb_6__4_/left_bottom_grid_pin_34_ sb_6__4_/left_bottom_grid_pin_35_
+ sb_6__4_/left_bottom_grid_pin_36_ sb_6__4_/left_bottom_grid_pin_37_ sb_6__4_/left_bottom_grid_pin_38_
+ sb_6__4_/left_bottom_grid_pin_39_ sb_6__4_/left_bottom_grid_pin_40_ sb_6__4_/left_bottom_grid_pin_41_
+ sb_6__4_/prog_clk_0_N_in sb_6__4_/prog_clk_1_E_out sb_6__4_/prog_clk_1_N_in sb_6__4_/prog_clk_1_W_out
+ sb_6__4_/prog_clk_2_E_out sb_6__4_/prog_clk_2_N_in sb_6__4_/prog_clk_2_N_out sb_6__4_/prog_clk_2_S_out
+ sb_6__4_/prog_clk_2_W_out sb_6__4_/prog_clk_3_E_out sb_6__4_/prog_clk_3_N_in sb_6__4_/prog_clk_3_N_out
+ sb_6__4_/prog_clk_3_S_out sb_6__4_/prog_clk_3_W_out sb_6__4_/right_bottom_grid_pin_34_
+ sb_6__4_/right_bottom_grid_pin_35_ sb_6__4_/right_bottom_grid_pin_36_ sb_6__4_/right_bottom_grid_pin_37_
+ sb_6__4_/right_bottom_grid_pin_38_ sb_6__4_/right_bottom_grid_pin_39_ sb_6__4_/right_bottom_grid_pin_40_
+ sb_6__4_/right_bottom_grid_pin_41_ sb_6__4_/top_left_grid_pin_42_ sb_6__4_/top_left_grid_pin_43_
+ sb_6__4_/top_left_grid_pin_44_ sb_6__4_/top_left_grid_pin_45_ sb_6__4_/top_left_grid_pin_46_
+ sb_6__4_/top_left_grid_pin_47_ sb_6__4_/top_left_grid_pin_48_ sb_6__4_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_8__2_ cbx_8__1_/SC_OUT_TOP grid_clb_8__2_/SC_OUT_BOT cbx_8__2_/SC_IN_BOT
+ cby_7__2_/Test_en_E_out grid_clb_8__2_/Test_en_E_out cby_7__2_/Test_en_E_out grid_clb_8__2_/Test_en_W_out
+ VGND VPWR cbx_8__1_/REGIN_FEEDTHROUGH grid_clb_8__2_/bottom_width_0_height_0__pin_51_
+ cby_7__2_/ccff_tail cby_8__2_/ccff_head cbx_8__1_/clk_1_N_out cbx_8__1_/clk_1_N_out
+ cby_8__2_/prog_clk_0_W_in cbx_8__1_/prog_clk_1_N_out grid_clb_8__2_/prog_clk_0_N_out
+ cbx_8__1_/prog_clk_1_N_out cbx_8__1_/prog_clk_0_N_in grid_clb_8__2_/prog_clk_0_W_out
+ cby_8__2_/left_grid_pin_16_ cby_8__2_/left_grid_pin_17_ cby_8__2_/left_grid_pin_18_
+ cby_8__2_/left_grid_pin_19_ cby_8__2_/left_grid_pin_20_ cby_8__2_/left_grid_pin_21_
+ cby_8__2_/left_grid_pin_22_ cby_8__2_/left_grid_pin_23_ cby_8__2_/left_grid_pin_24_
+ cby_8__2_/left_grid_pin_25_ cby_8__2_/left_grid_pin_26_ cby_8__2_/left_grid_pin_27_
+ cby_8__2_/left_grid_pin_28_ cby_8__2_/left_grid_pin_29_ cby_8__2_/left_grid_pin_30_
+ cby_8__2_/left_grid_pin_31_ sb_8__1_/top_left_grid_pin_42_ sb_8__2_/bottom_left_grid_pin_42_
+ sb_8__1_/top_left_grid_pin_43_ sb_8__2_/bottom_left_grid_pin_43_ sb_8__1_/top_left_grid_pin_44_
+ sb_8__2_/bottom_left_grid_pin_44_ sb_8__1_/top_left_grid_pin_45_ sb_8__2_/bottom_left_grid_pin_45_
+ sb_8__1_/top_left_grid_pin_46_ sb_8__2_/bottom_left_grid_pin_46_ sb_8__1_/top_left_grid_pin_47_
+ sb_8__2_/bottom_left_grid_pin_47_ sb_8__1_/top_left_grid_pin_48_ sb_8__2_/bottom_left_grid_pin_48_
+ sb_8__1_/top_left_grid_pin_49_ sb_8__2_/bottom_left_grid_pin_49_ cbx_8__2_/bottom_grid_pin_0_
+ cbx_8__2_/bottom_grid_pin_10_ cbx_8__2_/bottom_grid_pin_11_ cbx_8__2_/bottom_grid_pin_12_
+ cbx_8__2_/bottom_grid_pin_13_ cbx_8__2_/bottom_grid_pin_14_ cbx_8__2_/bottom_grid_pin_15_
+ cbx_8__2_/bottom_grid_pin_1_ cbx_8__2_/bottom_grid_pin_2_ cbx_8__2_/REGOUT_FEEDTHROUGH
+ grid_clb_8__2_/top_width_0_height_0__pin_33_ sb_8__2_/left_bottom_grid_pin_34_ sb_7__2_/right_bottom_grid_pin_34_
+ sb_8__2_/left_bottom_grid_pin_35_ sb_7__2_/right_bottom_grid_pin_35_ sb_8__2_/left_bottom_grid_pin_36_
+ sb_7__2_/right_bottom_grid_pin_36_ sb_8__2_/left_bottom_grid_pin_37_ sb_7__2_/right_bottom_grid_pin_37_
+ sb_8__2_/left_bottom_grid_pin_38_ sb_7__2_/right_bottom_grid_pin_38_ sb_8__2_/left_bottom_grid_pin_39_
+ sb_7__2_/right_bottom_grid_pin_39_ cbx_8__2_/bottom_grid_pin_3_ sb_8__2_/left_bottom_grid_pin_40_
+ sb_7__2_/right_bottom_grid_pin_40_ sb_8__2_/left_bottom_grid_pin_41_ sb_7__2_/right_bottom_grid_pin_41_
+ cbx_8__2_/bottom_grid_pin_4_ cbx_8__2_/bottom_grid_pin_5_ cbx_8__2_/bottom_grid_pin_6_
+ cbx_8__2_/bottom_grid_pin_7_ cbx_8__2_/bottom_grid_pin_8_ cbx_8__2_/bottom_grid_pin_9_
+ grid_clb
Xgrid_clb_1__7_ cbx_1__7_/SC_OUT_BOT cbx_1__6_/SC_IN_TOP grid_clb_1__7_/SC_OUT_TOP
+ cby_1__7_/Test_en_W_out grid_clb_1__7_/Test_en_E_out cby_1__7_/Test_en_W_out grid_clb_1__7_/Test_en_W_out
+ VGND VPWR cbx_1__6_/REGIN_FEEDTHROUGH grid_clb_1__7_/bottom_width_0_height_0__pin_51_
+ cby_0__7_/ccff_tail cby_1__7_/ccff_head cbx_1__7_/clk_1_S_out cbx_1__7_/clk_1_S_out
+ cby_1__7_/prog_clk_0_W_in cbx_1__7_/prog_clk_1_S_out grid_clb_1__7_/prog_clk_0_N_out
+ cbx_1__7_/prog_clk_1_S_out cbx_1__6_/prog_clk_0_N_in cby_0__7_/prog_clk_0_E_in cby_1__7_/left_grid_pin_16_
+ cby_1__7_/left_grid_pin_17_ cby_1__7_/left_grid_pin_18_ cby_1__7_/left_grid_pin_19_
+ cby_1__7_/left_grid_pin_20_ cby_1__7_/left_grid_pin_21_ cby_1__7_/left_grid_pin_22_
+ cby_1__7_/left_grid_pin_23_ cby_1__7_/left_grid_pin_24_ cby_1__7_/left_grid_pin_25_
+ cby_1__7_/left_grid_pin_26_ cby_1__7_/left_grid_pin_27_ cby_1__7_/left_grid_pin_28_
+ cby_1__7_/left_grid_pin_29_ cby_1__7_/left_grid_pin_30_ cby_1__7_/left_grid_pin_31_
+ sb_1__6_/top_left_grid_pin_42_ sb_1__7_/bottom_left_grid_pin_42_ sb_1__6_/top_left_grid_pin_43_
+ sb_1__7_/bottom_left_grid_pin_43_ sb_1__6_/top_left_grid_pin_44_ sb_1__7_/bottom_left_grid_pin_44_
+ sb_1__6_/top_left_grid_pin_45_ sb_1__7_/bottom_left_grid_pin_45_ sb_1__6_/top_left_grid_pin_46_
+ sb_1__7_/bottom_left_grid_pin_46_ sb_1__6_/top_left_grid_pin_47_ sb_1__7_/bottom_left_grid_pin_47_
+ sb_1__6_/top_left_grid_pin_48_ sb_1__7_/bottom_left_grid_pin_48_ sb_1__6_/top_left_grid_pin_49_
+ sb_1__7_/bottom_left_grid_pin_49_ cbx_1__7_/bottom_grid_pin_0_ cbx_1__7_/bottom_grid_pin_10_
+ cbx_1__7_/bottom_grid_pin_11_ cbx_1__7_/bottom_grid_pin_12_ cbx_1__7_/bottom_grid_pin_13_
+ cbx_1__7_/bottom_grid_pin_14_ cbx_1__7_/bottom_grid_pin_15_ cbx_1__7_/bottom_grid_pin_1_
+ cbx_1__7_/bottom_grid_pin_2_ cbx_1__7_/REGOUT_FEEDTHROUGH grid_clb_1__7_/top_width_0_height_0__pin_33_
+ sb_1__7_/left_bottom_grid_pin_34_ sb_0__7_/right_bottom_grid_pin_34_ sb_1__7_/left_bottom_grid_pin_35_
+ sb_0__7_/right_bottom_grid_pin_35_ sb_1__7_/left_bottom_grid_pin_36_ sb_0__7_/right_bottom_grid_pin_36_
+ sb_1__7_/left_bottom_grid_pin_37_ sb_0__7_/right_bottom_grid_pin_37_ sb_1__7_/left_bottom_grid_pin_38_
+ sb_0__7_/right_bottom_grid_pin_38_ sb_1__7_/left_bottom_grid_pin_39_ sb_0__7_/right_bottom_grid_pin_39_
+ cbx_1__7_/bottom_grid_pin_3_ sb_1__7_/left_bottom_grid_pin_40_ sb_0__7_/right_bottom_grid_pin_40_
+ sb_1__7_/left_bottom_grid_pin_41_ sb_0__7_/right_bottom_grid_pin_41_ cbx_1__7_/bottom_grid_pin_4_
+ cbx_1__7_/bottom_grid_pin_5_ cbx_1__7_/bottom_grid_pin_6_ cbx_1__7_/bottom_grid_pin_7_
+ cbx_1__7_/bottom_grid_pin_8_ cbx_1__7_/bottom_grid_pin_9_ grid_clb
Xsb_3__1_ sb_3__1_/Test_en_N_out sb_3__1_/Test_en_S_in VGND VPWR sb_3__1_/bottom_left_grid_pin_42_
+ sb_3__1_/bottom_left_grid_pin_43_ sb_3__1_/bottom_left_grid_pin_44_ sb_3__1_/bottom_left_grid_pin_45_
+ sb_3__1_/bottom_left_grid_pin_46_ sb_3__1_/bottom_left_grid_pin_47_ sb_3__1_/bottom_left_grid_pin_48_
+ sb_3__1_/bottom_left_grid_pin_49_ sb_3__1_/ccff_head sb_3__1_/ccff_tail sb_3__1_/chanx_left_in[0]
+ sb_3__1_/chanx_left_in[10] sb_3__1_/chanx_left_in[11] sb_3__1_/chanx_left_in[12]
+ sb_3__1_/chanx_left_in[13] sb_3__1_/chanx_left_in[14] sb_3__1_/chanx_left_in[15]
+ sb_3__1_/chanx_left_in[16] sb_3__1_/chanx_left_in[17] sb_3__1_/chanx_left_in[18]
+ sb_3__1_/chanx_left_in[19] sb_3__1_/chanx_left_in[1] sb_3__1_/chanx_left_in[2] sb_3__1_/chanx_left_in[3]
+ sb_3__1_/chanx_left_in[4] sb_3__1_/chanx_left_in[5] sb_3__1_/chanx_left_in[6] sb_3__1_/chanx_left_in[7]
+ sb_3__1_/chanx_left_in[8] sb_3__1_/chanx_left_in[9] sb_3__1_/chanx_left_out[0] sb_3__1_/chanx_left_out[10]
+ sb_3__1_/chanx_left_out[11] sb_3__1_/chanx_left_out[12] sb_3__1_/chanx_left_out[13]
+ sb_3__1_/chanx_left_out[14] sb_3__1_/chanx_left_out[15] sb_3__1_/chanx_left_out[16]
+ sb_3__1_/chanx_left_out[17] sb_3__1_/chanx_left_out[18] sb_3__1_/chanx_left_out[19]
+ sb_3__1_/chanx_left_out[1] sb_3__1_/chanx_left_out[2] sb_3__1_/chanx_left_out[3]
+ sb_3__1_/chanx_left_out[4] sb_3__1_/chanx_left_out[5] sb_3__1_/chanx_left_out[6]
+ sb_3__1_/chanx_left_out[7] sb_3__1_/chanx_left_out[8] sb_3__1_/chanx_left_out[9]
+ sb_3__1_/chanx_right_in[0] sb_3__1_/chanx_right_in[10] sb_3__1_/chanx_right_in[11]
+ sb_3__1_/chanx_right_in[12] sb_3__1_/chanx_right_in[13] sb_3__1_/chanx_right_in[14]
+ sb_3__1_/chanx_right_in[15] sb_3__1_/chanx_right_in[16] sb_3__1_/chanx_right_in[17]
+ sb_3__1_/chanx_right_in[18] sb_3__1_/chanx_right_in[19] sb_3__1_/chanx_right_in[1]
+ sb_3__1_/chanx_right_in[2] sb_3__1_/chanx_right_in[3] sb_3__1_/chanx_right_in[4]
+ sb_3__1_/chanx_right_in[5] sb_3__1_/chanx_right_in[6] sb_3__1_/chanx_right_in[7]
+ sb_3__1_/chanx_right_in[8] sb_3__1_/chanx_right_in[9] cbx_4__1_/chanx_left_in[0]
+ cbx_4__1_/chanx_left_in[10] cbx_4__1_/chanx_left_in[11] cbx_4__1_/chanx_left_in[12]
+ cbx_4__1_/chanx_left_in[13] cbx_4__1_/chanx_left_in[14] cbx_4__1_/chanx_left_in[15]
+ cbx_4__1_/chanx_left_in[16] cbx_4__1_/chanx_left_in[17] cbx_4__1_/chanx_left_in[18]
+ cbx_4__1_/chanx_left_in[19] cbx_4__1_/chanx_left_in[1] cbx_4__1_/chanx_left_in[2]
+ cbx_4__1_/chanx_left_in[3] cbx_4__1_/chanx_left_in[4] cbx_4__1_/chanx_left_in[5]
+ cbx_4__1_/chanx_left_in[6] cbx_4__1_/chanx_left_in[7] cbx_4__1_/chanx_left_in[8]
+ cbx_4__1_/chanx_left_in[9] cby_3__1_/chany_top_out[0] cby_3__1_/chany_top_out[10]
+ cby_3__1_/chany_top_out[11] cby_3__1_/chany_top_out[12] cby_3__1_/chany_top_out[13]
+ cby_3__1_/chany_top_out[14] cby_3__1_/chany_top_out[15] cby_3__1_/chany_top_out[16]
+ cby_3__1_/chany_top_out[17] cby_3__1_/chany_top_out[18] cby_3__1_/chany_top_out[19]
+ cby_3__1_/chany_top_out[1] cby_3__1_/chany_top_out[2] cby_3__1_/chany_top_out[3]
+ cby_3__1_/chany_top_out[4] cby_3__1_/chany_top_out[5] cby_3__1_/chany_top_out[6]
+ cby_3__1_/chany_top_out[7] cby_3__1_/chany_top_out[8] cby_3__1_/chany_top_out[9]
+ cby_3__1_/chany_top_in[0] cby_3__1_/chany_top_in[10] cby_3__1_/chany_top_in[11]
+ cby_3__1_/chany_top_in[12] cby_3__1_/chany_top_in[13] cby_3__1_/chany_top_in[14]
+ cby_3__1_/chany_top_in[15] cby_3__1_/chany_top_in[16] cby_3__1_/chany_top_in[17]
+ cby_3__1_/chany_top_in[18] cby_3__1_/chany_top_in[19] cby_3__1_/chany_top_in[1]
+ cby_3__1_/chany_top_in[2] cby_3__1_/chany_top_in[3] cby_3__1_/chany_top_in[4] cby_3__1_/chany_top_in[5]
+ cby_3__1_/chany_top_in[6] cby_3__1_/chany_top_in[7] cby_3__1_/chany_top_in[8] cby_3__1_/chany_top_in[9]
+ sb_3__1_/chany_top_in[0] sb_3__1_/chany_top_in[10] sb_3__1_/chany_top_in[11] sb_3__1_/chany_top_in[12]
+ sb_3__1_/chany_top_in[13] sb_3__1_/chany_top_in[14] sb_3__1_/chany_top_in[15] sb_3__1_/chany_top_in[16]
+ sb_3__1_/chany_top_in[17] sb_3__1_/chany_top_in[18] sb_3__1_/chany_top_in[19] sb_3__1_/chany_top_in[1]
+ sb_3__1_/chany_top_in[2] sb_3__1_/chany_top_in[3] sb_3__1_/chany_top_in[4] sb_3__1_/chany_top_in[5]
+ sb_3__1_/chany_top_in[6] sb_3__1_/chany_top_in[7] sb_3__1_/chany_top_in[8] sb_3__1_/chany_top_in[9]
+ sb_3__1_/chany_top_out[0] sb_3__1_/chany_top_out[10] sb_3__1_/chany_top_out[11]
+ sb_3__1_/chany_top_out[12] sb_3__1_/chany_top_out[13] sb_3__1_/chany_top_out[14]
+ sb_3__1_/chany_top_out[15] sb_3__1_/chany_top_out[16] sb_3__1_/chany_top_out[17]
+ sb_3__1_/chany_top_out[18] sb_3__1_/chany_top_out[19] sb_3__1_/chany_top_out[1]
+ sb_3__1_/chany_top_out[2] sb_3__1_/chany_top_out[3] sb_3__1_/chany_top_out[4] sb_3__1_/chany_top_out[5]
+ sb_3__1_/chany_top_out[6] sb_3__1_/chany_top_out[7] sb_3__1_/chany_top_out[8] sb_3__1_/chany_top_out[9]
+ sb_3__1_/clk_1_E_out sb_3__1_/clk_1_N_in sb_3__1_/clk_1_W_out sb_3__1_/clk_2_E_out
+ sb_3__1_/clk_2_N_in sb_3__1_/clk_2_N_out sb_3__1_/clk_2_S_out sb_3__1_/clk_2_W_out
+ sb_3__1_/clk_3_E_out sb_3__1_/clk_3_N_in sb_3__1_/clk_3_N_out sb_3__1_/clk_3_S_out
+ sb_3__1_/clk_3_W_out sb_3__1_/left_bottom_grid_pin_34_ sb_3__1_/left_bottom_grid_pin_35_
+ sb_3__1_/left_bottom_grid_pin_36_ sb_3__1_/left_bottom_grid_pin_37_ sb_3__1_/left_bottom_grid_pin_38_
+ sb_3__1_/left_bottom_grid_pin_39_ sb_3__1_/left_bottom_grid_pin_40_ sb_3__1_/left_bottom_grid_pin_41_
+ sb_3__1_/prog_clk_0_N_in sb_3__1_/prog_clk_1_E_out sb_3__1_/prog_clk_1_N_in sb_3__1_/prog_clk_1_W_out
+ sb_3__1_/prog_clk_2_E_out sb_3__1_/prog_clk_2_N_in sb_3__1_/prog_clk_2_N_out sb_3__1_/prog_clk_2_S_out
+ sb_3__1_/prog_clk_2_W_out sb_3__1_/prog_clk_3_E_out sb_3__1_/prog_clk_3_N_in sb_3__1_/prog_clk_3_N_out
+ sb_3__1_/prog_clk_3_S_out sb_3__1_/prog_clk_3_W_out sb_3__1_/right_bottom_grid_pin_34_
+ sb_3__1_/right_bottom_grid_pin_35_ sb_3__1_/right_bottom_grid_pin_36_ sb_3__1_/right_bottom_grid_pin_37_
+ sb_3__1_/right_bottom_grid_pin_38_ sb_3__1_/right_bottom_grid_pin_39_ sb_3__1_/right_bottom_grid_pin_40_
+ sb_3__1_/right_bottom_grid_pin_41_ sb_3__1_/top_left_grid_pin_42_ sb_3__1_/top_left_grid_pin_43_
+ sb_3__1_/top_left_grid_pin_44_ sb_3__1_/top_left_grid_pin_45_ sb_3__1_/top_left_grid_pin_46_
+ sb_3__1_/top_left_grid_pin_47_ sb_3__1_/top_left_grid_pin_48_ sb_3__1_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_5__8_ cby_5__8_/Test_en_W_in cby_5__8_/Test_en_E_out cby_5__8_/Test_en_N_out
+ cby_5__8_/Test_en_W_in cby_5__8_/Test_en_W_in cby_5__8_/Test_en_W_out VGND VPWR
+ cby_5__8_/ccff_head cby_5__8_/ccff_tail sb_5__7_/chany_top_out[0] sb_5__7_/chany_top_out[10]
+ sb_5__7_/chany_top_out[11] sb_5__7_/chany_top_out[12] sb_5__7_/chany_top_out[13]
+ sb_5__7_/chany_top_out[14] sb_5__7_/chany_top_out[15] sb_5__7_/chany_top_out[16]
+ sb_5__7_/chany_top_out[17] sb_5__7_/chany_top_out[18] sb_5__7_/chany_top_out[19]
+ sb_5__7_/chany_top_out[1] sb_5__7_/chany_top_out[2] sb_5__7_/chany_top_out[3] sb_5__7_/chany_top_out[4]
+ sb_5__7_/chany_top_out[5] sb_5__7_/chany_top_out[6] sb_5__7_/chany_top_out[7] sb_5__7_/chany_top_out[8]
+ sb_5__7_/chany_top_out[9] sb_5__7_/chany_top_in[0] sb_5__7_/chany_top_in[10] sb_5__7_/chany_top_in[11]
+ sb_5__7_/chany_top_in[12] sb_5__7_/chany_top_in[13] sb_5__7_/chany_top_in[14] sb_5__7_/chany_top_in[15]
+ sb_5__7_/chany_top_in[16] sb_5__7_/chany_top_in[17] sb_5__7_/chany_top_in[18] sb_5__7_/chany_top_in[19]
+ sb_5__7_/chany_top_in[1] sb_5__7_/chany_top_in[2] sb_5__7_/chany_top_in[3] sb_5__7_/chany_top_in[4]
+ sb_5__7_/chany_top_in[5] sb_5__7_/chany_top_in[6] sb_5__7_/chany_top_in[7] sb_5__7_/chany_top_in[8]
+ sb_5__7_/chany_top_in[9] cby_5__8_/chany_top_in[0] cby_5__8_/chany_top_in[10] cby_5__8_/chany_top_in[11]
+ cby_5__8_/chany_top_in[12] cby_5__8_/chany_top_in[13] cby_5__8_/chany_top_in[14]
+ cby_5__8_/chany_top_in[15] cby_5__8_/chany_top_in[16] cby_5__8_/chany_top_in[17]
+ cby_5__8_/chany_top_in[18] cby_5__8_/chany_top_in[19] cby_5__8_/chany_top_in[1]
+ cby_5__8_/chany_top_in[2] cby_5__8_/chany_top_in[3] cby_5__8_/chany_top_in[4] cby_5__8_/chany_top_in[5]
+ cby_5__8_/chany_top_in[6] cby_5__8_/chany_top_in[7] cby_5__8_/chany_top_in[8] cby_5__8_/chany_top_in[9]
+ cby_5__8_/chany_top_out[0] cby_5__8_/chany_top_out[10] cby_5__8_/chany_top_out[11]
+ cby_5__8_/chany_top_out[12] cby_5__8_/chany_top_out[13] cby_5__8_/chany_top_out[14]
+ cby_5__8_/chany_top_out[15] cby_5__8_/chany_top_out[16] cby_5__8_/chany_top_out[17]
+ cby_5__8_/chany_top_out[18] cby_5__8_/chany_top_out[19] cby_5__8_/chany_top_out[1]
+ cby_5__8_/chany_top_out[2] cby_5__8_/chany_top_out[3] cby_5__8_/chany_top_out[4]
+ cby_5__8_/chany_top_out[5] cby_5__8_/chany_top_out[6] cby_5__8_/chany_top_out[7]
+ cby_5__8_/chany_top_out[8] cby_5__8_/chany_top_out[9] cby_5__8_/clk_2_N_out cby_5__8_/clk_2_S_in
+ cby_5__8_/clk_2_S_out cby_5__8_/clk_3_N_out cby_5__8_/clk_3_S_in cby_5__8_/clk_3_S_out
+ cby_5__8_/left_grid_pin_16_ cby_5__8_/left_grid_pin_17_ cby_5__8_/left_grid_pin_18_
+ cby_5__8_/left_grid_pin_19_ cby_5__8_/left_grid_pin_20_ cby_5__8_/left_grid_pin_21_
+ cby_5__8_/left_grid_pin_22_ cby_5__8_/left_grid_pin_23_ cby_5__8_/left_grid_pin_24_
+ cby_5__8_/left_grid_pin_25_ cby_5__8_/left_grid_pin_26_ cby_5__8_/left_grid_pin_27_
+ cby_5__8_/left_grid_pin_28_ cby_5__8_/left_grid_pin_29_ cby_5__8_/left_grid_pin_30_
+ cby_5__8_/left_grid_pin_31_ sb_5__8_/prog_clk_0_S_in sb_5__7_/prog_clk_0_N_in cby_5__8_/prog_clk_0_W_in
+ cby_5__8_/prog_clk_2_N_out cby_5__8_/prog_clk_2_S_in cby_5__8_/prog_clk_2_S_out
+ cby_5__8_/prog_clk_3_N_out cby_5__8_/prog_clk_3_S_in cby_5__8_/prog_clk_3_S_out
+ cby_1__1_
Xcby_2__5_ cby_2__5_/Test_en_W_in cby_2__5_/Test_en_E_out cby_2__5_/Test_en_N_out
+ cby_2__5_/Test_en_W_in cby_2__5_/Test_en_W_in cby_2__5_/Test_en_W_out VGND VPWR
+ cby_2__5_/ccff_head cby_2__5_/ccff_tail sb_2__4_/chany_top_out[0] sb_2__4_/chany_top_out[10]
+ sb_2__4_/chany_top_out[11] sb_2__4_/chany_top_out[12] sb_2__4_/chany_top_out[13]
+ sb_2__4_/chany_top_out[14] sb_2__4_/chany_top_out[15] sb_2__4_/chany_top_out[16]
+ sb_2__4_/chany_top_out[17] sb_2__4_/chany_top_out[18] sb_2__4_/chany_top_out[19]
+ sb_2__4_/chany_top_out[1] sb_2__4_/chany_top_out[2] sb_2__4_/chany_top_out[3] sb_2__4_/chany_top_out[4]
+ sb_2__4_/chany_top_out[5] sb_2__4_/chany_top_out[6] sb_2__4_/chany_top_out[7] sb_2__4_/chany_top_out[8]
+ sb_2__4_/chany_top_out[9] sb_2__4_/chany_top_in[0] sb_2__4_/chany_top_in[10] sb_2__4_/chany_top_in[11]
+ sb_2__4_/chany_top_in[12] sb_2__4_/chany_top_in[13] sb_2__4_/chany_top_in[14] sb_2__4_/chany_top_in[15]
+ sb_2__4_/chany_top_in[16] sb_2__4_/chany_top_in[17] sb_2__4_/chany_top_in[18] sb_2__4_/chany_top_in[19]
+ sb_2__4_/chany_top_in[1] sb_2__4_/chany_top_in[2] sb_2__4_/chany_top_in[3] sb_2__4_/chany_top_in[4]
+ sb_2__4_/chany_top_in[5] sb_2__4_/chany_top_in[6] sb_2__4_/chany_top_in[7] sb_2__4_/chany_top_in[8]
+ sb_2__4_/chany_top_in[9] cby_2__5_/chany_top_in[0] cby_2__5_/chany_top_in[10] cby_2__5_/chany_top_in[11]
+ cby_2__5_/chany_top_in[12] cby_2__5_/chany_top_in[13] cby_2__5_/chany_top_in[14]
+ cby_2__5_/chany_top_in[15] cby_2__5_/chany_top_in[16] cby_2__5_/chany_top_in[17]
+ cby_2__5_/chany_top_in[18] cby_2__5_/chany_top_in[19] cby_2__5_/chany_top_in[1]
+ cby_2__5_/chany_top_in[2] cby_2__5_/chany_top_in[3] cby_2__5_/chany_top_in[4] cby_2__5_/chany_top_in[5]
+ cby_2__5_/chany_top_in[6] cby_2__5_/chany_top_in[7] cby_2__5_/chany_top_in[8] cby_2__5_/chany_top_in[9]
+ cby_2__5_/chany_top_out[0] cby_2__5_/chany_top_out[10] cby_2__5_/chany_top_out[11]
+ cby_2__5_/chany_top_out[12] cby_2__5_/chany_top_out[13] cby_2__5_/chany_top_out[14]
+ cby_2__5_/chany_top_out[15] cby_2__5_/chany_top_out[16] cby_2__5_/chany_top_out[17]
+ cby_2__5_/chany_top_out[18] cby_2__5_/chany_top_out[19] cby_2__5_/chany_top_out[1]
+ cby_2__5_/chany_top_out[2] cby_2__5_/chany_top_out[3] cby_2__5_/chany_top_out[4]
+ cby_2__5_/chany_top_out[5] cby_2__5_/chany_top_out[6] cby_2__5_/chany_top_out[7]
+ cby_2__5_/chany_top_out[8] cby_2__5_/chany_top_out[9] cby_2__5_/clk_2_N_out cby_2__5_/clk_2_S_in
+ cby_2__5_/clk_2_S_out sb_2__5_/clk_3_N_in sb_2__4_/clk_3_N_out cby_2__5_/clk_3_S_out
+ cby_2__5_/left_grid_pin_16_ cby_2__5_/left_grid_pin_17_ cby_2__5_/left_grid_pin_18_
+ cby_2__5_/left_grid_pin_19_ cby_2__5_/left_grid_pin_20_ cby_2__5_/left_grid_pin_21_
+ cby_2__5_/left_grid_pin_22_ cby_2__5_/left_grid_pin_23_ cby_2__5_/left_grid_pin_24_
+ cby_2__5_/left_grid_pin_25_ cby_2__5_/left_grid_pin_26_ cby_2__5_/left_grid_pin_27_
+ cby_2__5_/left_grid_pin_28_ cby_2__5_/left_grid_pin_29_ cby_2__5_/left_grid_pin_30_
+ cby_2__5_/left_grid_pin_31_ cby_2__5_/prog_clk_0_N_out sb_2__4_/prog_clk_0_N_in
+ cby_2__5_/prog_clk_0_W_in cby_2__5_/prog_clk_2_N_out cby_2__5_/prog_clk_2_S_in cby_2__5_/prog_clk_2_S_out
+ sb_2__5_/prog_clk_3_N_in sb_2__4_/prog_clk_3_N_out cby_2__5_/prog_clk_3_S_out cby_1__1_
Xgrid_clb_8__1_ cbx_8__0_/SC_OUT_TOP grid_clb_8__1_/SC_OUT_BOT cbx_8__1_/SC_IN_BOT
+ cby_7__1_/Test_en_E_out grid_clb_8__1_/Test_en_E_out cby_7__1_/Test_en_E_out grid_clb_8__1_/Test_en_W_out
+ VGND VPWR grid_clb_8__1_/bottom_width_0_height_0__pin_50_ grid_clb_8__1_/bottom_width_0_height_0__pin_51_
+ cby_7__1_/ccff_tail cby_8__1_/ccff_head cbx_8__1_/clk_1_S_out cbx_8__1_/clk_1_S_out
+ cby_8__1_/prog_clk_0_W_in cbx_8__1_/prog_clk_1_S_out grid_clb_8__1_/prog_clk_0_N_out
+ cbx_8__1_/prog_clk_1_S_out cbx_8__0_/prog_clk_0_N_in grid_clb_8__1_/prog_clk_0_W_out
+ cby_8__1_/left_grid_pin_16_ cby_8__1_/left_grid_pin_17_ cby_8__1_/left_grid_pin_18_
+ cby_8__1_/left_grid_pin_19_ cby_8__1_/left_grid_pin_20_ cby_8__1_/left_grid_pin_21_
+ cby_8__1_/left_grid_pin_22_ cby_8__1_/left_grid_pin_23_ cby_8__1_/left_grid_pin_24_
+ cby_8__1_/left_grid_pin_25_ cby_8__1_/left_grid_pin_26_ cby_8__1_/left_grid_pin_27_
+ cby_8__1_/left_grid_pin_28_ cby_8__1_/left_grid_pin_29_ cby_8__1_/left_grid_pin_30_
+ cby_8__1_/left_grid_pin_31_ sb_8__0_/top_left_grid_pin_42_ sb_8__1_/bottom_left_grid_pin_42_
+ sb_8__0_/top_left_grid_pin_43_ sb_8__1_/bottom_left_grid_pin_43_ sb_8__0_/top_left_grid_pin_44_
+ sb_8__1_/bottom_left_grid_pin_44_ sb_8__0_/top_left_grid_pin_45_ sb_8__1_/bottom_left_grid_pin_45_
+ sb_8__0_/top_left_grid_pin_46_ sb_8__1_/bottom_left_grid_pin_46_ sb_8__0_/top_left_grid_pin_47_
+ sb_8__1_/bottom_left_grid_pin_47_ sb_8__0_/top_left_grid_pin_48_ sb_8__1_/bottom_left_grid_pin_48_
+ sb_8__0_/top_left_grid_pin_49_ sb_8__1_/bottom_left_grid_pin_49_ cbx_8__1_/bottom_grid_pin_0_
+ cbx_8__1_/bottom_grid_pin_10_ cbx_8__1_/bottom_grid_pin_11_ cbx_8__1_/bottom_grid_pin_12_
+ cbx_8__1_/bottom_grid_pin_13_ cbx_8__1_/bottom_grid_pin_14_ cbx_8__1_/bottom_grid_pin_15_
+ cbx_8__1_/bottom_grid_pin_1_ cbx_8__1_/bottom_grid_pin_2_ cbx_8__1_/REGOUT_FEEDTHROUGH
+ grid_clb_8__1_/top_width_0_height_0__pin_33_ sb_8__1_/left_bottom_grid_pin_34_ sb_7__1_/right_bottom_grid_pin_34_
+ sb_8__1_/left_bottom_grid_pin_35_ sb_7__1_/right_bottom_grid_pin_35_ sb_8__1_/left_bottom_grid_pin_36_
+ sb_7__1_/right_bottom_grid_pin_36_ sb_8__1_/left_bottom_grid_pin_37_ sb_7__1_/right_bottom_grid_pin_37_
+ sb_8__1_/left_bottom_grid_pin_38_ sb_7__1_/right_bottom_grid_pin_38_ sb_8__1_/left_bottom_grid_pin_39_
+ sb_7__1_/right_bottom_grid_pin_39_ cbx_8__1_/bottom_grid_pin_3_ sb_8__1_/left_bottom_grid_pin_40_
+ sb_7__1_/right_bottom_grid_pin_40_ sb_8__1_/left_bottom_grid_pin_41_ sb_7__1_/right_bottom_grid_pin_41_
+ cbx_8__1_/bottom_grid_pin_4_ cbx_8__1_/bottom_grid_pin_5_ cbx_8__1_/bottom_grid_pin_6_
+ cbx_8__1_/bottom_grid_pin_7_ cbx_8__1_/bottom_grid_pin_8_ cbx_8__1_/bottom_grid_pin_9_
+ grid_clb
Xcbx_2__6_ cbx_2__6_/REGIN_FEEDTHROUGH cbx_2__6_/REGOUT_FEEDTHROUGH cbx_2__6_/SC_IN_BOT
+ cbx_2__6_/SC_IN_TOP cbx_2__6_/SC_OUT_BOT cbx_2__6_/SC_OUT_TOP VGND VPWR cbx_2__6_/bottom_grid_pin_0_
+ cbx_2__6_/bottom_grid_pin_10_ cbx_2__6_/bottom_grid_pin_11_ cbx_2__6_/bottom_grid_pin_12_
+ cbx_2__6_/bottom_grid_pin_13_ cbx_2__6_/bottom_grid_pin_14_ cbx_2__6_/bottom_grid_pin_15_
+ cbx_2__6_/bottom_grid_pin_1_ cbx_2__6_/bottom_grid_pin_2_ cbx_2__6_/bottom_grid_pin_3_
+ cbx_2__6_/bottom_grid_pin_4_ cbx_2__6_/bottom_grid_pin_5_ cbx_2__6_/bottom_grid_pin_6_
+ cbx_2__6_/bottom_grid_pin_7_ cbx_2__6_/bottom_grid_pin_8_ cbx_2__6_/bottom_grid_pin_9_
+ sb_2__6_/ccff_tail sb_1__6_/ccff_head cbx_2__6_/chanx_left_in[0] cbx_2__6_/chanx_left_in[10]
+ cbx_2__6_/chanx_left_in[11] cbx_2__6_/chanx_left_in[12] cbx_2__6_/chanx_left_in[13]
+ cbx_2__6_/chanx_left_in[14] cbx_2__6_/chanx_left_in[15] cbx_2__6_/chanx_left_in[16]
+ cbx_2__6_/chanx_left_in[17] cbx_2__6_/chanx_left_in[18] cbx_2__6_/chanx_left_in[19]
+ cbx_2__6_/chanx_left_in[1] cbx_2__6_/chanx_left_in[2] cbx_2__6_/chanx_left_in[3]
+ cbx_2__6_/chanx_left_in[4] cbx_2__6_/chanx_left_in[5] cbx_2__6_/chanx_left_in[6]
+ cbx_2__6_/chanx_left_in[7] cbx_2__6_/chanx_left_in[8] cbx_2__6_/chanx_left_in[9]
+ sb_1__6_/chanx_right_in[0] sb_1__6_/chanx_right_in[10] sb_1__6_/chanx_right_in[11]
+ sb_1__6_/chanx_right_in[12] sb_1__6_/chanx_right_in[13] sb_1__6_/chanx_right_in[14]
+ sb_1__6_/chanx_right_in[15] sb_1__6_/chanx_right_in[16] sb_1__6_/chanx_right_in[17]
+ sb_1__6_/chanx_right_in[18] sb_1__6_/chanx_right_in[19] sb_1__6_/chanx_right_in[1]
+ sb_1__6_/chanx_right_in[2] sb_1__6_/chanx_right_in[3] sb_1__6_/chanx_right_in[4]
+ sb_1__6_/chanx_right_in[5] sb_1__6_/chanx_right_in[6] sb_1__6_/chanx_right_in[7]
+ sb_1__6_/chanx_right_in[8] sb_1__6_/chanx_right_in[9] sb_2__6_/chanx_left_out[0]
+ sb_2__6_/chanx_left_out[10] sb_2__6_/chanx_left_out[11] sb_2__6_/chanx_left_out[12]
+ sb_2__6_/chanx_left_out[13] sb_2__6_/chanx_left_out[14] sb_2__6_/chanx_left_out[15]
+ sb_2__6_/chanx_left_out[16] sb_2__6_/chanx_left_out[17] sb_2__6_/chanx_left_out[18]
+ sb_2__6_/chanx_left_out[19] sb_2__6_/chanx_left_out[1] sb_2__6_/chanx_left_out[2]
+ sb_2__6_/chanx_left_out[3] sb_2__6_/chanx_left_out[4] sb_2__6_/chanx_left_out[5]
+ sb_2__6_/chanx_left_out[6] sb_2__6_/chanx_left_out[7] sb_2__6_/chanx_left_out[8]
+ sb_2__6_/chanx_left_out[9] sb_2__6_/chanx_left_in[0] sb_2__6_/chanx_left_in[10]
+ sb_2__6_/chanx_left_in[11] sb_2__6_/chanx_left_in[12] sb_2__6_/chanx_left_in[13]
+ sb_2__6_/chanx_left_in[14] sb_2__6_/chanx_left_in[15] sb_2__6_/chanx_left_in[16]
+ sb_2__6_/chanx_left_in[17] sb_2__6_/chanx_left_in[18] sb_2__6_/chanx_left_in[19]
+ sb_2__6_/chanx_left_in[1] sb_2__6_/chanx_left_in[2] sb_2__6_/chanx_left_in[3] sb_2__6_/chanx_left_in[4]
+ sb_2__6_/chanx_left_in[5] sb_2__6_/chanx_left_in[6] sb_2__6_/chanx_left_in[7] sb_2__6_/chanx_left_in[8]
+ sb_2__6_/chanx_left_in[9] cbx_2__6_/clk_1_N_out cbx_2__6_/clk_1_S_out cbx_2__6_/clk_1_W_in
+ cbx_2__6_/clk_2_E_out sb_2__6_/clk_2_W_out sb_1__6_/clk_2_N_in cbx_2__6_/clk_3_E_out
+ cbx_2__6_/clk_3_W_in cbx_2__6_/clk_3_W_out cbx_2__6_/prog_clk_0_N_in cbx_2__6_/prog_clk_0_W_out
+ cbx_2__6_/prog_clk_1_N_out cbx_2__6_/prog_clk_1_S_out cbx_2__6_/prog_clk_1_W_in
+ cbx_2__6_/prog_clk_2_E_out sb_2__6_/prog_clk_2_W_out sb_1__6_/prog_clk_2_N_in cbx_2__6_/prog_clk_3_E_out
+ cbx_2__6_/prog_clk_3_W_in cbx_2__6_/prog_clk_3_W_out cbx_1__1_
Xgrid_clb_1__6_ cbx_1__6_/SC_OUT_BOT cbx_1__5_/SC_IN_TOP grid_clb_1__6_/SC_OUT_TOP
+ cby_1__6_/Test_en_W_out grid_clb_1__6_/Test_en_E_out cby_1__6_/Test_en_W_out grid_clb_1__6_/Test_en_W_out
+ VGND VPWR cbx_1__5_/REGIN_FEEDTHROUGH grid_clb_1__6_/bottom_width_0_height_0__pin_51_
+ cby_0__6_/ccff_tail cby_1__6_/ccff_head cbx_1__5_/clk_1_N_out cbx_1__5_/clk_1_N_out
+ cby_1__6_/prog_clk_0_W_in cbx_1__5_/prog_clk_1_N_out grid_clb_1__6_/prog_clk_0_N_out
+ cbx_1__5_/prog_clk_1_N_out cbx_1__5_/prog_clk_0_N_in cby_0__6_/prog_clk_0_E_in cby_1__6_/left_grid_pin_16_
+ cby_1__6_/left_grid_pin_17_ cby_1__6_/left_grid_pin_18_ cby_1__6_/left_grid_pin_19_
+ cby_1__6_/left_grid_pin_20_ cby_1__6_/left_grid_pin_21_ cby_1__6_/left_grid_pin_22_
+ cby_1__6_/left_grid_pin_23_ cby_1__6_/left_grid_pin_24_ cby_1__6_/left_grid_pin_25_
+ cby_1__6_/left_grid_pin_26_ cby_1__6_/left_grid_pin_27_ cby_1__6_/left_grid_pin_28_
+ cby_1__6_/left_grid_pin_29_ cby_1__6_/left_grid_pin_30_ cby_1__6_/left_grid_pin_31_
+ sb_1__5_/top_left_grid_pin_42_ sb_1__6_/bottom_left_grid_pin_42_ sb_1__5_/top_left_grid_pin_43_
+ sb_1__6_/bottom_left_grid_pin_43_ sb_1__5_/top_left_grid_pin_44_ sb_1__6_/bottom_left_grid_pin_44_
+ sb_1__5_/top_left_grid_pin_45_ sb_1__6_/bottom_left_grid_pin_45_ sb_1__5_/top_left_grid_pin_46_
+ sb_1__6_/bottom_left_grid_pin_46_ sb_1__5_/top_left_grid_pin_47_ sb_1__6_/bottom_left_grid_pin_47_
+ sb_1__5_/top_left_grid_pin_48_ sb_1__6_/bottom_left_grid_pin_48_ sb_1__5_/top_left_grid_pin_49_
+ sb_1__6_/bottom_left_grid_pin_49_ cbx_1__6_/bottom_grid_pin_0_ cbx_1__6_/bottom_grid_pin_10_
+ cbx_1__6_/bottom_grid_pin_11_ cbx_1__6_/bottom_grid_pin_12_ cbx_1__6_/bottom_grid_pin_13_
+ cbx_1__6_/bottom_grid_pin_14_ cbx_1__6_/bottom_grid_pin_15_ cbx_1__6_/bottom_grid_pin_1_
+ cbx_1__6_/bottom_grid_pin_2_ cbx_1__6_/REGOUT_FEEDTHROUGH grid_clb_1__6_/top_width_0_height_0__pin_33_
+ sb_1__6_/left_bottom_grid_pin_34_ sb_0__6_/right_bottom_grid_pin_34_ sb_1__6_/left_bottom_grid_pin_35_
+ sb_0__6_/right_bottom_grid_pin_35_ sb_1__6_/left_bottom_grid_pin_36_ sb_0__6_/right_bottom_grid_pin_36_
+ sb_1__6_/left_bottom_grid_pin_37_ sb_0__6_/right_bottom_grid_pin_37_ sb_1__6_/left_bottom_grid_pin_38_
+ sb_0__6_/right_bottom_grid_pin_38_ sb_1__6_/left_bottom_grid_pin_39_ sb_0__6_/right_bottom_grid_pin_39_
+ cbx_1__6_/bottom_grid_pin_3_ sb_1__6_/left_bottom_grid_pin_40_ sb_0__6_/right_bottom_grid_pin_40_
+ sb_1__6_/left_bottom_grid_pin_41_ sb_0__6_/right_bottom_grid_pin_41_ cbx_1__6_/bottom_grid_pin_4_
+ cbx_1__6_/bottom_grid_pin_5_ cbx_1__6_/bottom_grid_pin_6_ cbx_1__6_/bottom_grid_pin_7_
+ cbx_1__6_/bottom_grid_pin_8_ cbx_1__6_/bottom_grid_pin_9_ grid_clb
Xsb_6__3_ sb_6__3_/Test_en_N_out sb_6__3_/Test_en_S_in VGND VPWR sb_6__3_/bottom_left_grid_pin_42_
+ sb_6__3_/bottom_left_grid_pin_43_ sb_6__3_/bottom_left_grid_pin_44_ sb_6__3_/bottom_left_grid_pin_45_
+ sb_6__3_/bottom_left_grid_pin_46_ sb_6__3_/bottom_left_grid_pin_47_ sb_6__3_/bottom_left_grid_pin_48_
+ sb_6__3_/bottom_left_grid_pin_49_ sb_6__3_/ccff_head sb_6__3_/ccff_tail sb_6__3_/chanx_left_in[0]
+ sb_6__3_/chanx_left_in[10] sb_6__3_/chanx_left_in[11] sb_6__3_/chanx_left_in[12]
+ sb_6__3_/chanx_left_in[13] sb_6__3_/chanx_left_in[14] sb_6__3_/chanx_left_in[15]
+ sb_6__3_/chanx_left_in[16] sb_6__3_/chanx_left_in[17] sb_6__3_/chanx_left_in[18]
+ sb_6__3_/chanx_left_in[19] sb_6__3_/chanx_left_in[1] sb_6__3_/chanx_left_in[2] sb_6__3_/chanx_left_in[3]
+ sb_6__3_/chanx_left_in[4] sb_6__3_/chanx_left_in[5] sb_6__3_/chanx_left_in[6] sb_6__3_/chanx_left_in[7]
+ sb_6__3_/chanx_left_in[8] sb_6__3_/chanx_left_in[9] sb_6__3_/chanx_left_out[0] sb_6__3_/chanx_left_out[10]
+ sb_6__3_/chanx_left_out[11] sb_6__3_/chanx_left_out[12] sb_6__3_/chanx_left_out[13]
+ sb_6__3_/chanx_left_out[14] sb_6__3_/chanx_left_out[15] sb_6__3_/chanx_left_out[16]
+ sb_6__3_/chanx_left_out[17] sb_6__3_/chanx_left_out[18] sb_6__3_/chanx_left_out[19]
+ sb_6__3_/chanx_left_out[1] sb_6__3_/chanx_left_out[2] sb_6__3_/chanx_left_out[3]
+ sb_6__3_/chanx_left_out[4] sb_6__3_/chanx_left_out[5] sb_6__3_/chanx_left_out[6]
+ sb_6__3_/chanx_left_out[7] sb_6__3_/chanx_left_out[8] sb_6__3_/chanx_left_out[9]
+ sb_6__3_/chanx_right_in[0] sb_6__3_/chanx_right_in[10] sb_6__3_/chanx_right_in[11]
+ sb_6__3_/chanx_right_in[12] sb_6__3_/chanx_right_in[13] sb_6__3_/chanx_right_in[14]
+ sb_6__3_/chanx_right_in[15] sb_6__3_/chanx_right_in[16] sb_6__3_/chanx_right_in[17]
+ sb_6__3_/chanx_right_in[18] sb_6__3_/chanx_right_in[19] sb_6__3_/chanx_right_in[1]
+ sb_6__3_/chanx_right_in[2] sb_6__3_/chanx_right_in[3] sb_6__3_/chanx_right_in[4]
+ sb_6__3_/chanx_right_in[5] sb_6__3_/chanx_right_in[6] sb_6__3_/chanx_right_in[7]
+ sb_6__3_/chanx_right_in[8] sb_6__3_/chanx_right_in[9] cbx_7__3_/chanx_left_in[0]
+ cbx_7__3_/chanx_left_in[10] cbx_7__3_/chanx_left_in[11] cbx_7__3_/chanx_left_in[12]
+ cbx_7__3_/chanx_left_in[13] cbx_7__3_/chanx_left_in[14] cbx_7__3_/chanx_left_in[15]
+ cbx_7__3_/chanx_left_in[16] cbx_7__3_/chanx_left_in[17] cbx_7__3_/chanx_left_in[18]
+ cbx_7__3_/chanx_left_in[19] cbx_7__3_/chanx_left_in[1] cbx_7__3_/chanx_left_in[2]
+ cbx_7__3_/chanx_left_in[3] cbx_7__3_/chanx_left_in[4] cbx_7__3_/chanx_left_in[5]
+ cbx_7__3_/chanx_left_in[6] cbx_7__3_/chanx_left_in[7] cbx_7__3_/chanx_left_in[8]
+ cbx_7__3_/chanx_left_in[9] cby_6__3_/chany_top_out[0] cby_6__3_/chany_top_out[10]
+ cby_6__3_/chany_top_out[11] cby_6__3_/chany_top_out[12] cby_6__3_/chany_top_out[13]
+ cby_6__3_/chany_top_out[14] cby_6__3_/chany_top_out[15] cby_6__3_/chany_top_out[16]
+ cby_6__3_/chany_top_out[17] cby_6__3_/chany_top_out[18] cby_6__3_/chany_top_out[19]
+ cby_6__3_/chany_top_out[1] cby_6__3_/chany_top_out[2] cby_6__3_/chany_top_out[3]
+ cby_6__3_/chany_top_out[4] cby_6__3_/chany_top_out[5] cby_6__3_/chany_top_out[6]
+ cby_6__3_/chany_top_out[7] cby_6__3_/chany_top_out[8] cby_6__3_/chany_top_out[9]
+ cby_6__3_/chany_top_in[0] cby_6__3_/chany_top_in[10] cby_6__3_/chany_top_in[11]
+ cby_6__3_/chany_top_in[12] cby_6__3_/chany_top_in[13] cby_6__3_/chany_top_in[14]
+ cby_6__3_/chany_top_in[15] cby_6__3_/chany_top_in[16] cby_6__3_/chany_top_in[17]
+ cby_6__3_/chany_top_in[18] cby_6__3_/chany_top_in[19] cby_6__3_/chany_top_in[1]
+ cby_6__3_/chany_top_in[2] cby_6__3_/chany_top_in[3] cby_6__3_/chany_top_in[4] cby_6__3_/chany_top_in[5]
+ cby_6__3_/chany_top_in[6] cby_6__3_/chany_top_in[7] cby_6__3_/chany_top_in[8] cby_6__3_/chany_top_in[9]
+ sb_6__3_/chany_top_in[0] sb_6__3_/chany_top_in[10] sb_6__3_/chany_top_in[11] sb_6__3_/chany_top_in[12]
+ sb_6__3_/chany_top_in[13] sb_6__3_/chany_top_in[14] sb_6__3_/chany_top_in[15] sb_6__3_/chany_top_in[16]
+ sb_6__3_/chany_top_in[17] sb_6__3_/chany_top_in[18] sb_6__3_/chany_top_in[19] sb_6__3_/chany_top_in[1]
+ sb_6__3_/chany_top_in[2] sb_6__3_/chany_top_in[3] sb_6__3_/chany_top_in[4] sb_6__3_/chany_top_in[5]
+ sb_6__3_/chany_top_in[6] sb_6__3_/chany_top_in[7] sb_6__3_/chany_top_in[8] sb_6__3_/chany_top_in[9]
+ sb_6__3_/chany_top_out[0] sb_6__3_/chany_top_out[10] sb_6__3_/chany_top_out[11]
+ sb_6__3_/chany_top_out[12] sb_6__3_/chany_top_out[13] sb_6__3_/chany_top_out[14]
+ sb_6__3_/chany_top_out[15] sb_6__3_/chany_top_out[16] sb_6__3_/chany_top_out[17]
+ sb_6__3_/chany_top_out[18] sb_6__3_/chany_top_out[19] sb_6__3_/chany_top_out[1]
+ sb_6__3_/chany_top_out[2] sb_6__3_/chany_top_out[3] sb_6__3_/chany_top_out[4] sb_6__3_/chany_top_out[5]
+ sb_6__3_/chany_top_out[6] sb_6__3_/chany_top_out[7] sb_6__3_/chany_top_out[8] sb_6__3_/chany_top_out[9]
+ sb_6__3_/clk_1_E_out sb_6__3_/clk_1_N_in sb_6__3_/clk_1_W_out sb_6__3_/clk_2_E_out
+ sb_6__3_/clk_2_N_in sb_6__3_/clk_2_N_out sb_6__3_/clk_2_S_out sb_6__3_/clk_2_W_out
+ sb_6__3_/clk_3_E_out sb_6__3_/clk_3_N_in sb_6__3_/clk_3_N_out sb_6__3_/clk_3_S_out
+ sb_6__3_/clk_3_W_out sb_6__3_/left_bottom_grid_pin_34_ sb_6__3_/left_bottom_grid_pin_35_
+ sb_6__3_/left_bottom_grid_pin_36_ sb_6__3_/left_bottom_grid_pin_37_ sb_6__3_/left_bottom_grid_pin_38_
+ sb_6__3_/left_bottom_grid_pin_39_ sb_6__3_/left_bottom_grid_pin_40_ sb_6__3_/left_bottom_grid_pin_41_
+ sb_6__3_/prog_clk_0_N_in sb_6__3_/prog_clk_1_E_out sb_6__3_/prog_clk_1_N_in sb_6__3_/prog_clk_1_W_out
+ sb_6__3_/prog_clk_2_E_out sb_6__3_/prog_clk_2_N_in sb_6__3_/prog_clk_2_N_out sb_6__3_/prog_clk_2_S_out
+ sb_6__3_/prog_clk_2_W_out sb_6__3_/prog_clk_3_E_out sb_6__3_/prog_clk_3_N_in sb_6__3_/prog_clk_3_N_out
+ sb_6__3_/prog_clk_3_S_out sb_6__3_/prog_clk_3_W_out sb_6__3_/right_bottom_grid_pin_34_
+ sb_6__3_/right_bottom_grid_pin_35_ sb_6__3_/right_bottom_grid_pin_36_ sb_6__3_/right_bottom_grid_pin_37_
+ sb_6__3_/right_bottom_grid_pin_38_ sb_6__3_/right_bottom_grid_pin_39_ sb_6__3_/right_bottom_grid_pin_40_
+ sb_6__3_/right_bottom_grid_pin_41_ sb_6__3_/top_left_grid_pin_42_ sb_6__3_/top_left_grid_pin_43_
+ sb_6__3_/top_left_grid_pin_44_ sb_6__3_/top_left_grid_pin_45_ sb_6__3_/top_left_grid_pin_46_
+ sb_6__3_/top_left_grid_pin_47_ sb_6__3_/top_left_grid_pin_48_ sb_6__3_/top_left_grid_pin_49_
+ sb_1__1_
Xsb_3__0_ sb_3__0_/SC_IN_TOP sb_3__0_/SC_OUT_TOP sb_3__0_/Test_en_N_out sb_3__0_/Test_en_S_in
+ VGND VPWR sb_3__0_/ccff_head sb_3__0_/ccff_tail sb_3__0_/chanx_left_in[0] sb_3__0_/chanx_left_in[10]
+ sb_3__0_/chanx_left_in[11] sb_3__0_/chanx_left_in[12] sb_3__0_/chanx_left_in[13]
+ sb_3__0_/chanx_left_in[14] sb_3__0_/chanx_left_in[15] sb_3__0_/chanx_left_in[16]
+ sb_3__0_/chanx_left_in[17] sb_3__0_/chanx_left_in[18] sb_3__0_/chanx_left_in[19]
+ sb_3__0_/chanx_left_in[1] sb_3__0_/chanx_left_in[2] sb_3__0_/chanx_left_in[3] sb_3__0_/chanx_left_in[4]
+ sb_3__0_/chanx_left_in[5] sb_3__0_/chanx_left_in[6] sb_3__0_/chanx_left_in[7] sb_3__0_/chanx_left_in[8]
+ sb_3__0_/chanx_left_in[9] sb_3__0_/chanx_left_out[0] sb_3__0_/chanx_left_out[10]
+ sb_3__0_/chanx_left_out[11] sb_3__0_/chanx_left_out[12] sb_3__0_/chanx_left_out[13]
+ sb_3__0_/chanx_left_out[14] sb_3__0_/chanx_left_out[15] sb_3__0_/chanx_left_out[16]
+ sb_3__0_/chanx_left_out[17] sb_3__0_/chanx_left_out[18] sb_3__0_/chanx_left_out[19]
+ sb_3__0_/chanx_left_out[1] sb_3__0_/chanx_left_out[2] sb_3__0_/chanx_left_out[3]
+ sb_3__0_/chanx_left_out[4] sb_3__0_/chanx_left_out[5] sb_3__0_/chanx_left_out[6]
+ sb_3__0_/chanx_left_out[7] sb_3__0_/chanx_left_out[8] sb_3__0_/chanx_left_out[9]
+ sb_3__0_/chanx_right_in[0] sb_3__0_/chanx_right_in[10] sb_3__0_/chanx_right_in[11]
+ sb_3__0_/chanx_right_in[12] sb_3__0_/chanx_right_in[13] sb_3__0_/chanx_right_in[14]
+ sb_3__0_/chanx_right_in[15] sb_3__0_/chanx_right_in[16] sb_3__0_/chanx_right_in[17]
+ sb_3__0_/chanx_right_in[18] sb_3__0_/chanx_right_in[19] sb_3__0_/chanx_right_in[1]
+ sb_3__0_/chanx_right_in[2] sb_3__0_/chanx_right_in[3] sb_3__0_/chanx_right_in[4]
+ sb_3__0_/chanx_right_in[5] sb_3__0_/chanx_right_in[6] sb_3__0_/chanx_right_in[7]
+ sb_3__0_/chanx_right_in[8] sb_3__0_/chanx_right_in[9] cbx_4__0_/chanx_left_in[0]
+ cbx_4__0_/chanx_left_in[10] cbx_4__0_/chanx_left_in[11] cbx_4__0_/chanx_left_in[12]
+ cbx_4__0_/chanx_left_in[13] cbx_4__0_/chanx_left_in[14] cbx_4__0_/chanx_left_in[15]
+ cbx_4__0_/chanx_left_in[16] cbx_4__0_/chanx_left_in[17] cbx_4__0_/chanx_left_in[18]
+ cbx_4__0_/chanx_left_in[19] cbx_4__0_/chanx_left_in[1] cbx_4__0_/chanx_left_in[2]
+ cbx_4__0_/chanx_left_in[3] cbx_4__0_/chanx_left_in[4] cbx_4__0_/chanx_left_in[5]
+ cbx_4__0_/chanx_left_in[6] cbx_4__0_/chanx_left_in[7] cbx_4__0_/chanx_left_in[8]
+ cbx_4__0_/chanx_left_in[9] sb_3__0_/chany_top_in[0] sb_3__0_/chany_top_in[10] sb_3__0_/chany_top_in[11]
+ sb_3__0_/chany_top_in[12] sb_3__0_/chany_top_in[13] sb_3__0_/chany_top_in[14] sb_3__0_/chany_top_in[15]
+ sb_3__0_/chany_top_in[16] sb_3__0_/chany_top_in[17] sb_3__0_/chany_top_in[18] sb_3__0_/chany_top_in[19]
+ sb_3__0_/chany_top_in[1] sb_3__0_/chany_top_in[2] sb_3__0_/chany_top_in[3] sb_3__0_/chany_top_in[4]
+ sb_3__0_/chany_top_in[5] sb_3__0_/chany_top_in[6] sb_3__0_/chany_top_in[7] sb_3__0_/chany_top_in[8]
+ sb_3__0_/chany_top_in[9] sb_3__0_/chany_top_out[0] sb_3__0_/chany_top_out[10] sb_3__0_/chany_top_out[11]
+ sb_3__0_/chany_top_out[12] sb_3__0_/chany_top_out[13] sb_3__0_/chany_top_out[14]
+ sb_3__0_/chany_top_out[15] sb_3__0_/chany_top_out[16] sb_3__0_/chany_top_out[17]
+ sb_3__0_/chany_top_out[18] sb_3__0_/chany_top_out[19] sb_3__0_/chany_top_out[1]
+ sb_3__0_/chany_top_out[2] sb_3__0_/chany_top_out[3] sb_3__0_/chany_top_out[4] sb_3__0_/chany_top_out[5]
+ sb_3__0_/chany_top_out[6] sb_3__0_/chany_top_out[7] sb_3__0_/chany_top_out[8] sb_3__0_/chany_top_out[9]
+ sb_3__0_/clk_3_N_out sb_3__0_/clk_3_S_in sb_3__0_/left_bottom_grid_pin_11_ sb_3__0_/left_bottom_grid_pin_13_
+ sb_3__0_/left_bottom_grid_pin_15_ sb_3__0_/left_bottom_grid_pin_17_ sb_3__0_/left_bottom_grid_pin_1_
+ sb_3__0_/left_bottom_grid_pin_3_ sb_3__0_/left_bottom_grid_pin_5_ sb_3__0_/left_bottom_grid_pin_7_
+ sb_3__0_/left_bottom_grid_pin_9_ sb_3__0_/prog_clk_0_N_in sb_3__0_/prog_clk_3_N_out
+ sb_3__0_/prog_clk_3_S_in sb_3__0_/right_bottom_grid_pin_11_ sb_3__0_/right_bottom_grid_pin_13_
+ sb_3__0_/right_bottom_grid_pin_15_ sb_3__0_/right_bottom_grid_pin_17_ sb_3__0_/right_bottom_grid_pin_1_
+ sb_3__0_/right_bottom_grid_pin_3_ sb_3__0_/right_bottom_grid_pin_5_ sb_3__0_/right_bottom_grid_pin_7_
+ sb_3__0_/right_bottom_grid_pin_9_ sb_3__0_/top_left_grid_pin_42_ sb_3__0_/top_left_grid_pin_43_
+ sb_3__0_/top_left_grid_pin_44_ sb_3__0_/top_left_grid_pin_45_ sb_3__0_/top_left_grid_pin_46_
+ sb_3__0_/top_left_grid_pin_47_ sb_3__0_/top_left_grid_pin_48_ sb_3__0_/top_left_grid_pin_49_
+ sb_1__0_
Xcby_5__7_ cby_5__7_/Test_en_W_in cby_5__7_/Test_en_E_out cby_5__7_/Test_en_N_out
+ cby_5__7_/Test_en_W_in cby_5__7_/Test_en_W_in cby_5__7_/Test_en_W_out VGND VPWR
+ cby_5__7_/ccff_head cby_5__7_/ccff_tail sb_5__6_/chany_top_out[0] sb_5__6_/chany_top_out[10]
+ sb_5__6_/chany_top_out[11] sb_5__6_/chany_top_out[12] sb_5__6_/chany_top_out[13]
+ sb_5__6_/chany_top_out[14] sb_5__6_/chany_top_out[15] sb_5__6_/chany_top_out[16]
+ sb_5__6_/chany_top_out[17] sb_5__6_/chany_top_out[18] sb_5__6_/chany_top_out[19]
+ sb_5__6_/chany_top_out[1] sb_5__6_/chany_top_out[2] sb_5__6_/chany_top_out[3] sb_5__6_/chany_top_out[4]
+ sb_5__6_/chany_top_out[5] sb_5__6_/chany_top_out[6] sb_5__6_/chany_top_out[7] sb_5__6_/chany_top_out[8]
+ sb_5__6_/chany_top_out[9] sb_5__6_/chany_top_in[0] sb_5__6_/chany_top_in[10] sb_5__6_/chany_top_in[11]
+ sb_5__6_/chany_top_in[12] sb_5__6_/chany_top_in[13] sb_5__6_/chany_top_in[14] sb_5__6_/chany_top_in[15]
+ sb_5__6_/chany_top_in[16] sb_5__6_/chany_top_in[17] sb_5__6_/chany_top_in[18] sb_5__6_/chany_top_in[19]
+ sb_5__6_/chany_top_in[1] sb_5__6_/chany_top_in[2] sb_5__6_/chany_top_in[3] sb_5__6_/chany_top_in[4]
+ sb_5__6_/chany_top_in[5] sb_5__6_/chany_top_in[6] sb_5__6_/chany_top_in[7] sb_5__6_/chany_top_in[8]
+ sb_5__6_/chany_top_in[9] cby_5__7_/chany_top_in[0] cby_5__7_/chany_top_in[10] cby_5__7_/chany_top_in[11]
+ cby_5__7_/chany_top_in[12] cby_5__7_/chany_top_in[13] cby_5__7_/chany_top_in[14]
+ cby_5__7_/chany_top_in[15] cby_5__7_/chany_top_in[16] cby_5__7_/chany_top_in[17]
+ cby_5__7_/chany_top_in[18] cby_5__7_/chany_top_in[19] cby_5__7_/chany_top_in[1]
+ cby_5__7_/chany_top_in[2] cby_5__7_/chany_top_in[3] cby_5__7_/chany_top_in[4] cby_5__7_/chany_top_in[5]
+ cby_5__7_/chany_top_in[6] cby_5__7_/chany_top_in[7] cby_5__7_/chany_top_in[8] cby_5__7_/chany_top_in[9]
+ cby_5__7_/chany_top_out[0] cby_5__7_/chany_top_out[10] cby_5__7_/chany_top_out[11]
+ cby_5__7_/chany_top_out[12] cby_5__7_/chany_top_out[13] cby_5__7_/chany_top_out[14]
+ cby_5__7_/chany_top_out[15] cby_5__7_/chany_top_out[16] cby_5__7_/chany_top_out[17]
+ cby_5__7_/chany_top_out[18] cby_5__7_/chany_top_out[19] cby_5__7_/chany_top_out[1]
+ cby_5__7_/chany_top_out[2] cby_5__7_/chany_top_out[3] cby_5__7_/chany_top_out[4]
+ cby_5__7_/chany_top_out[5] cby_5__7_/chany_top_out[6] cby_5__7_/chany_top_out[7]
+ cby_5__7_/chany_top_out[8] cby_5__7_/chany_top_out[9] sb_5__7_/clk_1_N_in sb_5__6_/clk_2_N_out
+ cby_5__7_/clk_2_S_out cby_5__7_/clk_3_N_out cby_5__7_/clk_3_S_in cby_5__7_/clk_3_S_out
+ cby_5__7_/left_grid_pin_16_ cby_5__7_/left_grid_pin_17_ cby_5__7_/left_grid_pin_18_
+ cby_5__7_/left_grid_pin_19_ cby_5__7_/left_grid_pin_20_ cby_5__7_/left_grid_pin_21_
+ cby_5__7_/left_grid_pin_22_ cby_5__7_/left_grid_pin_23_ cby_5__7_/left_grid_pin_24_
+ cby_5__7_/left_grid_pin_25_ cby_5__7_/left_grid_pin_26_ cby_5__7_/left_grid_pin_27_
+ cby_5__7_/left_grid_pin_28_ cby_5__7_/left_grid_pin_29_ cby_5__7_/left_grid_pin_30_
+ cby_5__7_/left_grid_pin_31_ cby_5__7_/prog_clk_0_N_out sb_5__6_/prog_clk_0_N_in
+ cby_5__7_/prog_clk_0_W_in sb_5__7_/prog_clk_1_N_in sb_5__6_/prog_clk_2_N_out cby_5__7_/prog_clk_2_S_out
+ cby_5__7_/prog_clk_3_N_out cby_5__7_/prog_clk_3_S_in cby_5__7_/prog_clk_3_S_out
+ cby_1__1_
Xcby_2__4_ cby_2__4_/Test_en_W_in cby_2__4_/Test_en_E_out cby_2__4_/Test_en_N_out
+ cby_2__4_/Test_en_W_in cby_2__4_/Test_en_W_in cby_2__4_/Test_en_W_out VGND VPWR
+ cby_2__4_/ccff_head cby_2__4_/ccff_tail sb_2__3_/chany_top_out[0] sb_2__3_/chany_top_out[10]
+ sb_2__3_/chany_top_out[11] sb_2__3_/chany_top_out[12] sb_2__3_/chany_top_out[13]
+ sb_2__3_/chany_top_out[14] sb_2__3_/chany_top_out[15] sb_2__3_/chany_top_out[16]
+ sb_2__3_/chany_top_out[17] sb_2__3_/chany_top_out[18] sb_2__3_/chany_top_out[19]
+ sb_2__3_/chany_top_out[1] sb_2__3_/chany_top_out[2] sb_2__3_/chany_top_out[3] sb_2__3_/chany_top_out[4]
+ sb_2__3_/chany_top_out[5] sb_2__3_/chany_top_out[6] sb_2__3_/chany_top_out[7] sb_2__3_/chany_top_out[8]
+ sb_2__3_/chany_top_out[9] sb_2__3_/chany_top_in[0] sb_2__3_/chany_top_in[10] sb_2__3_/chany_top_in[11]
+ sb_2__3_/chany_top_in[12] sb_2__3_/chany_top_in[13] sb_2__3_/chany_top_in[14] sb_2__3_/chany_top_in[15]
+ sb_2__3_/chany_top_in[16] sb_2__3_/chany_top_in[17] sb_2__3_/chany_top_in[18] sb_2__3_/chany_top_in[19]
+ sb_2__3_/chany_top_in[1] sb_2__3_/chany_top_in[2] sb_2__3_/chany_top_in[3] sb_2__3_/chany_top_in[4]
+ sb_2__3_/chany_top_in[5] sb_2__3_/chany_top_in[6] sb_2__3_/chany_top_in[7] sb_2__3_/chany_top_in[8]
+ sb_2__3_/chany_top_in[9] cby_2__4_/chany_top_in[0] cby_2__4_/chany_top_in[10] cby_2__4_/chany_top_in[11]
+ cby_2__4_/chany_top_in[12] cby_2__4_/chany_top_in[13] cby_2__4_/chany_top_in[14]
+ cby_2__4_/chany_top_in[15] cby_2__4_/chany_top_in[16] cby_2__4_/chany_top_in[17]
+ cby_2__4_/chany_top_in[18] cby_2__4_/chany_top_in[19] cby_2__4_/chany_top_in[1]
+ cby_2__4_/chany_top_in[2] cby_2__4_/chany_top_in[3] cby_2__4_/chany_top_in[4] cby_2__4_/chany_top_in[5]
+ cby_2__4_/chany_top_in[6] cby_2__4_/chany_top_in[7] cby_2__4_/chany_top_in[8] cby_2__4_/chany_top_in[9]
+ cby_2__4_/chany_top_out[0] cby_2__4_/chany_top_out[10] cby_2__4_/chany_top_out[11]
+ cby_2__4_/chany_top_out[12] cby_2__4_/chany_top_out[13] cby_2__4_/chany_top_out[14]
+ cby_2__4_/chany_top_out[15] cby_2__4_/chany_top_out[16] cby_2__4_/chany_top_out[17]
+ cby_2__4_/chany_top_out[18] cby_2__4_/chany_top_out[19] cby_2__4_/chany_top_out[1]
+ cby_2__4_/chany_top_out[2] cby_2__4_/chany_top_out[3] cby_2__4_/chany_top_out[4]
+ cby_2__4_/chany_top_out[5] cby_2__4_/chany_top_out[6] cby_2__4_/chany_top_out[7]
+ cby_2__4_/chany_top_out[8] cby_2__4_/chany_top_out[9] cby_2__4_/clk_2_N_out cby_2__4_/clk_2_S_in
+ cby_2__4_/clk_2_S_out cby_2__4_/clk_3_N_out sb_2__4_/clk_3_S_out sb_2__3_/clk_3_N_in
+ cby_2__4_/left_grid_pin_16_ cby_2__4_/left_grid_pin_17_ cby_2__4_/left_grid_pin_18_
+ cby_2__4_/left_grid_pin_19_ cby_2__4_/left_grid_pin_20_ cby_2__4_/left_grid_pin_21_
+ cby_2__4_/left_grid_pin_22_ cby_2__4_/left_grid_pin_23_ cby_2__4_/left_grid_pin_24_
+ cby_2__4_/left_grid_pin_25_ cby_2__4_/left_grid_pin_26_ cby_2__4_/left_grid_pin_27_
+ cby_2__4_/left_grid_pin_28_ cby_2__4_/left_grid_pin_29_ cby_2__4_/left_grid_pin_30_
+ cby_2__4_/left_grid_pin_31_ cby_2__4_/prog_clk_0_N_out sb_2__3_/prog_clk_0_N_in
+ cby_2__4_/prog_clk_0_W_in cby_2__4_/prog_clk_2_N_out cby_2__4_/prog_clk_2_S_in cby_2__4_/prog_clk_2_S_out
+ cby_2__4_/prog_clk_3_N_out sb_2__4_/prog_clk_3_S_out sb_2__3_/prog_clk_3_N_in cby_1__1_
Xcbx_5__8_ IO_ISOL_N cbx_5__8_/SC_IN_BOT sb_4__8_/SC_OUT_BOT cbx_5__8_/SC_OUT_BOT
+ cbx_5__8_/SC_OUT_TOP VGND VPWR cbx_5__8_/bottom_grid_pin_0_ cbx_5__8_/bottom_grid_pin_10_
+ cbx_5__8_/bottom_grid_pin_11_ cbx_5__8_/bottom_grid_pin_12_ cbx_5__8_/bottom_grid_pin_13_
+ cbx_5__8_/bottom_grid_pin_14_ cbx_5__8_/bottom_grid_pin_15_ cbx_5__8_/bottom_grid_pin_1_
+ cbx_5__8_/bottom_grid_pin_2_ cbx_5__8_/bottom_grid_pin_3_ cbx_5__8_/bottom_grid_pin_4_
+ cbx_5__8_/bottom_grid_pin_5_ cbx_5__8_/bottom_grid_pin_6_ cbx_5__8_/bottom_grid_pin_7_
+ cbx_5__8_/bottom_grid_pin_8_ cbx_5__8_/bottom_grid_pin_9_ cbx_5__8_/top_grid_pin_0_
+ sb_5__8_/left_top_grid_pin_1_ sb_4__8_/right_top_grid_pin_1_ sb_5__8_/ccff_tail
+ sb_4__8_/ccff_head cbx_5__8_/chanx_left_in[0] cbx_5__8_/chanx_left_in[10] cbx_5__8_/chanx_left_in[11]
+ cbx_5__8_/chanx_left_in[12] cbx_5__8_/chanx_left_in[13] cbx_5__8_/chanx_left_in[14]
+ cbx_5__8_/chanx_left_in[15] cbx_5__8_/chanx_left_in[16] cbx_5__8_/chanx_left_in[17]
+ cbx_5__8_/chanx_left_in[18] cbx_5__8_/chanx_left_in[19] cbx_5__8_/chanx_left_in[1]
+ cbx_5__8_/chanx_left_in[2] cbx_5__8_/chanx_left_in[3] cbx_5__8_/chanx_left_in[4]
+ cbx_5__8_/chanx_left_in[5] cbx_5__8_/chanx_left_in[6] cbx_5__8_/chanx_left_in[7]
+ cbx_5__8_/chanx_left_in[8] cbx_5__8_/chanx_left_in[9] sb_4__8_/chanx_right_in[0]
+ sb_4__8_/chanx_right_in[10] sb_4__8_/chanx_right_in[11] sb_4__8_/chanx_right_in[12]
+ sb_4__8_/chanx_right_in[13] sb_4__8_/chanx_right_in[14] sb_4__8_/chanx_right_in[15]
+ sb_4__8_/chanx_right_in[16] sb_4__8_/chanx_right_in[17] sb_4__8_/chanx_right_in[18]
+ sb_4__8_/chanx_right_in[19] sb_4__8_/chanx_right_in[1] sb_4__8_/chanx_right_in[2]
+ sb_4__8_/chanx_right_in[3] sb_4__8_/chanx_right_in[4] sb_4__8_/chanx_right_in[5]
+ sb_4__8_/chanx_right_in[6] sb_4__8_/chanx_right_in[7] sb_4__8_/chanx_right_in[8]
+ sb_4__8_/chanx_right_in[9] sb_5__8_/chanx_left_out[0] sb_5__8_/chanx_left_out[10]
+ sb_5__8_/chanx_left_out[11] sb_5__8_/chanx_left_out[12] sb_5__8_/chanx_left_out[13]
+ sb_5__8_/chanx_left_out[14] sb_5__8_/chanx_left_out[15] sb_5__8_/chanx_left_out[16]
+ sb_5__8_/chanx_left_out[17] sb_5__8_/chanx_left_out[18] sb_5__8_/chanx_left_out[19]
+ sb_5__8_/chanx_left_out[1] sb_5__8_/chanx_left_out[2] sb_5__8_/chanx_left_out[3]
+ sb_5__8_/chanx_left_out[4] sb_5__8_/chanx_left_out[5] sb_5__8_/chanx_left_out[6]
+ sb_5__8_/chanx_left_out[7] sb_5__8_/chanx_left_out[8] sb_5__8_/chanx_left_out[9]
+ sb_5__8_/chanx_left_in[0] sb_5__8_/chanx_left_in[10] sb_5__8_/chanx_left_in[11]
+ sb_5__8_/chanx_left_in[12] sb_5__8_/chanx_left_in[13] sb_5__8_/chanx_left_in[14]
+ sb_5__8_/chanx_left_in[15] sb_5__8_/chanx_left_in[16] sb_5__8_/chanx_left_in[17]
+ sb_5__8_/chanx_left_in[18] sb_5__8_/chanx_left_in[19] sb_5__8_/chanx_left_in[1]
+ sb_5__8_/chanx_left_in[2] sb_5__8_/chanx_left_in[3] sb_5__8_/chanx_left_in[4] sb_5__8_/chanx_left_in[5]
+ sb_5__8_/chanx_left_in[6] sb_5__8_/chanx_left_in[7] sb_5__8_/chanx_left_in[8] sb_5__8_/chanx_left_in[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
+ cbx_5__8_/prog_clk_0_S_in cbx_5__8_/prog_clk_0_W_out cbx_5__8_/top_grid_pin_0_ cbx_1__2_
Xcbx_2__5_ cbx_2__5_/REGIN_FEEDTHROUGH cbx_2__5_/REGOUT_FEEDTHROUGH cbx_2__5_/SC_IN_BOT
+ cbx_2__5_/SC_IN_TOP cbx_2__5_/SC_OUT_BOT cbx_2__5_/SC_OUT_TOP VGND VPWR cbx_2__5_/bottom_grid_pin_0_
+ cbx_2__5_/bottom_grid_pin_10_ cbx_2__5_/bottom_grid_pin_11_ cbx_2__5_/bottom_grid_pin_12_
+ cbx_2__5_/bottom_grid_pin_13_ cbx_2__5_/bottom_grid_pin_14_ cbx_2__5_/bottom_grid_pin_15_
+ cbx_2__5_/bottom_grid_pin_1_ cbx_2__5_/bottom_grid_pin_2_ cbx_2__5_/bottom_grid_pin_3_
+ cbx_2__5_/bottom_grid_pin_4_ cbx_2__5_/bottom_grid_pin_5_ cbx_2__5_/bottom_grid_pin_6_
+ cbx_2__5_/bottom_grid_pin_7_ cbx_2__5_/bottom_grid_pin_8_ cbx_2__5_/bottom_grid_pin_9_
+ sb_2__5_/ccff_tail sb_1__5_/ccff_head cbx_2__5_/chanx_left_in[0] cbx_2__5_/chanx_left_in[10]
+ cbx_2__5_/chanx_left_in[11] cbx_2__5_/chanx_left_in[12] cbx_2__5_/chanx_left_in[13]
+ cbx_2__5_/chanx_left_in[14] cbx_2__5_/chanx_left_in[15] cbx_2__5_/chanx_left_in[16]
+ cbx_2__5_/chanx_left_in[17] cbx_2__5_/chanx_left_in[18] cbx_2__5_/chanx_left_in[19]
+ cbx_2__5_/chanx_left_in[1] cbx_2__5_/chanx_left_in[2] cbx_2__5_/chanx_left_in[3]
+ cbx_2__5_/chanx_left_in[4] cbx_2__5_/chanx_left_in[5] cbx_2__5_/chanx_left_in[6]
+ cbx_2__5_/chanx_left_in[7] cbx_2__5_/chanx_left_in[8] cbx_2__5_/chanx_left_in[9]
+ sb_1__5_/chanx_right_in[0] sb_1__5_/chanx_right_in[10] sb_1__5_/chanx_right_in[11]
+ sb_1__5_/chanx_right_in[12] sb_1__5_/chanx_right_in[13] sb_1__5_/chanx_right_in[14]
+ sb_1__5_/chanx_right_in[15] sb_1__5_/chanx_right_in[16] sb_1__5_/chanx_right_in[17]
+ sb_1__5_/chanx_right_in[18] sb_1__5_/chanx_right_in[19] sb_1__5_/chanx_right_in[1]
+ sb_1__5_/chanx_right_in[2] sb_1__5_/chanx_right_in[3] sb_1__5_/chanx_right_in[4]
+ sb_1__5_/chanx_right_in[5] sb_1__5_/chanx_right_in[6] sb_1__5_/chanx_right_in[7]
+ sb_1__5_/chanx_right_in[8] sb_1__5_/chanx_right_in[9] sb_2__5_/chanx_left_out[0]
+ sb_2__5_/chanx_left_out[10] sb_2__5_/chanx_left_out[11] sb_2__5_/chanx_left_out[12]
+ sb_2__5_/chanx_left_out[13] sb_2__5_/chanx_left_out[14] sb_2__5_/chanx_left_out[15]
+ sb_2__5_/chanx_left_out[16] sb_2__5_/chanx_left_out[17] sb_2__5_/chanx_left_out[18]
+ sb_2__5_/chanx_left_out[19] sb_2__5_/chanx_left_out[1] sb_2__5_/chanx_left_out[2]
+ sb_2__5_/chanx_left_out[3] sb_2__5_/chanx_left_out[4] sb_2__5_/chanx_left_out[5]
+ sb_2__5_/chanx_left_out[6] sb_2__5_/chanx_left_out[7] sb_2__5_/chanx_left_out[8]
+ sb_2__5_/chanx_left_out[9] sb_2__5_/chanx_left_in[0] sb_2__5_/chanx_left_in[10]
+ sb_2__5_/chanx_left_in[11] sb_2__5_/chanx_left_in[12] sb_2__5_/chanx_left_in[13]
+ sb_2__5_/chanx_left_in[14] sb_2__5_/chanx_left_in[15] sb_2__5_/chanx_left_in[16]
+ sb_2__5_/chanx_left_in[17] sb_2__5_/chanx_left_in[18] sb_2__5_/chanx_left_in[19]
+ sb_2__5_/chanx_left_in[1] sb_2__5_/chanx_left_in[2] sb_2__5_/chanx_left_in[3] sb_2__5_/chanx_left_in[4]
+ sb_2__5_/chanx_left_in[5] sb_2__5_/chanx_left_in[6] sb_2__5_/chanx_left_in[7] sb_2__5_/chanx_left_in[8]
+ sb_2__5_/chanx_left_in[9] cbx_2__5_/clk_1_N_out cbx_2__5_/clk_1_S_out sb_1__5_/clk_1_E_out
+ cbx_2__5_/clk_2_E_out cbx_2__5_/clk_2_W_in cbx_2__5_/clk_2_W_out cbx_2__5_/clk_3_E_out
+ cbx_2__5_/clk_3_W_in cbx_2__5_/clk_3_W_out cbx_2__5_/prog_clk_0_N_in cbx_2__5_/prog_clk_0_W_out
+ cbx_2__5_/prog_clk_1_N_out cbx_2__5_/prog_clk_1_S_out sb_1__5_/prog_clk_1_E_out
+ cbx_2__5_/prog_clk_2_E_out cbx_2__5_/prog_clk_2_W_in cbx_2__5_/prog_clk_2_W_out
+ cbx_2__5_/prog_clk_3_E_out cbx_2__5_/prog_clk_3_W_in cbx_2__5_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_4__8_ cbx_4__7_/SC_OUT_TOP grid_clb_4__8_/SC_OUT_BOT cbx_4__8_/SC_IN_BOT
+ cby_4__8_/Test_en_W_out grid_clb_4__8_/Test_en_E_out cby_4__8_/Test_en_W_out cby_3__8_/Test_en_W_in
+ VGND VPWR cbx_4__7_/REGIN_FEEDTHROUGH grid_clb_4__8_/bottom_width_0_height_0__pin_51_
+ cby_3__8_/ccff_tail cby_4__8_/ccff_head cbx_4__7_/clk_1_N_out cbx_4__7_/clk_1_N_out
+ cby_4__8_/prog_clk_0_W_in cbx_4__7_/prog_clk_1_N_out cbx_4__8_/prog_clk_0_S_in cbx_4__7_/prog_clk_1_N_out
+ cbx_4__7_/prog_clk_0_N_in grid_clb_4__8_/prog_clk_0_W_out cby_4__8_/left_grid_pin_16_
+ cby_4__8_/left_grid_pin_17_ cby_4__8_/left_grid_pin_18_ cby_4__8_/left_grid_pin_19_
+ cby_4__8_/left_grid_pin_20_ cby_4__8_/left_grid_pin_21_ cby_4__8_/left_grid_pin_22_
+ cby_4__8_/left_grid_pin_23_ cby_4__8_/left_grid_pin_24_ cby_4__8_/left_grid_pin_25_
+ cby_4__8_/left_grid_pin_26_ cby_4__8_/left_grid_pin_27_ cby_4__8_/left_grid_pin_28_
+ cby_4__8_/left_grid_pin_29_ cby_4__8_/left_grid_pin_30_ cby_4__8_/left_grid_pin_31_
+ sb_4__7_/top_left_grid_pin_42_ sb_4__8_/bottom_left_grid_pin_42_ sb_4__7_/top_left_grid_pin_43_
+ sb_4__8_/bottom_left_grid_pin_43_ sb_4__7_/top_left_grid_pin_44_ sb_4__8_/bottom_left_grid_pin_44_
+ sb_4__7_/top_left_grid_pin_45_ sb_4__8_/bottom_left_grid_pin_45_ sb_4__7_/top_left_grid_pin_46_
+ sb_4__8_/bottom_left_grid_pin_46_ sb_4__7_/top_left_grid_pin_47_ sb_4__8_/bottom_left_grid_pin_47_
+ sb_4__7_/top_left_grid_pin_48_ sb_4__8_/bottom_left_grid_pin_48_ sb_4__7_/top_left_grid_pin_49_
+ sb_4__8_/bottom_left_grid_pin_49_ cbx_4__8_/bottom_grid_pin_0_ cbx_4__8_/bottom_grid_pin_10_
+ cbx_4__8_/bottom_grid_pin_11_ cbx_4__8_/bottom_grid_pin_12_ cbx_4__8_/bottom_grid_pin_13_
+ cbx_4__8_/bottom_grid_pin_14_ cbx_4__8_/bottom_grid_pin_15_ cbx_4__8_/bottom_grid_pin_1_
+ cbx_4__8_/bottom_grid_pin_2_ tie_array/x[3] grid_clb_4__8_/top_width_0_height_0__pin_33_
+ sb_4__8_/left_bottom_grid_pin_34_ sb_3__8_/right_bottom_grid_pin_34_ sb_4__8_/left_bottom_grid_pin_35_
+ sb_3__8_/right_bottom_grid_pin_35_ sb_4__8_/left_bottom_grid_pin_36_ sb_3__8_/right_bottom_grid_pin_36_
+ sb_4__8_/left_bottom_grid_pin_37_ sb_3__8_/right_bottom_grid_pin_37_ sb_4__8_/left_bottom_grid_pin_38_
+ sb_3__8_/right_bottom_grid_pin_38_ sb_4__8_/left_bottom_grid_pin_39_ sb_3__8_/right_bottom_grid_pin_39_
+ cbx_4__8_/bottom_grid_pin_3_ sb_4__8_/left_bottom_grid_pin_40_ sb_3__8_/right_bottom_grid_pin_40_
+ sb_4__8_/left_bottom_grid_pin_41_ sb_3__8_/right_bottom_grid_pin_41_ cbx_4__8_/bottom_grid_pin_4_
+ cbx_4__8_/bottom_grid_pin_5_ cbx_4__8_/bottom_grid_pin_6_ cbx_4__8_/bottom_grid_pin_7_
+ cbx_4__8_/bottom_grid_pin_8_ cbx_4__8_/bottom_grid_pin_9_ grid_clb
Xgrid_clb_1__5_ cbx_1__5_/SC_OUT_BOT cbx_1__4_/SC_IN_TOP grid_clb_1__5_/SC_OUT_TOP
+ cby_1__5_/Test_en_W_out grid_clb_1__5_/Test_en_E_out cby_1__5_/Test_en_W_out grid_clb_1__5_/Test_en_W_out
+ VGND VPWR cbx_1__4_/REGIN_FEEDTHROUGH grid_clb_1__5_/bottom_width_0_height_0__pin_51_
+ cby_0__5_/ccff_tail cby_1__5_/ccff_head cbx_1__5_/clk_1_S_out cbx_1__5_/clk_1_S_out
+ cby_1__5_/prog_clk_0_W_in cbx_1__5_/prog_clk_1_S_out grid_clb_1__5_/prog_clk_0_N_out
+ cbx_1__5_/prog_clk_1_S_out cbx_1__4_/prog_clk_0_N_in cby_0__5_/prog_clk_0_E_in cby_1__5_/left_grid_pin_16_
+ cby_1__5_/left_grid_pin_17_ cby_1__5_/left_grid_pin_18_ cby_1__5_/left_grid_pin_19_
+ cby_1__5_/left_grid_pin_20_ cby_1__5_/left_grid_pin_21_ cby_1__5_/left_grid_pin_22_
+ cby_1__5_/left_grid_pin_23_ cby_1__5_/left_grid_pin_24_ cby_1__5_/left_grid_pin_25_
+ cby_1__5_/left_grid_pin_26_ cby_1__5_/left_grid_pin_27_ cby_1__5_/left_grid_pin_28_
+ cby_1__5_/left_grid_pin_29_ cby_1__5_/left_grid_pin_30_ cby_1__5_/left_grid_pin_31_
+ sb_1__4_/top_left_grid_pin_42_ sb_1__5_/bottom_left_grid_pin_42_ sb_1__4_/top_left_grid_pin_43_
+ sb_1__5_/bottom_left_grid_pin_43_ sb_1__4_/top_left_grid_pin_44_ sb_1__5_/bottom_left_grid_pin_44_
+ sb_1__4_/top_left_grid_pin_45_ sb_1__5_/bottom_left_grid_pin_45_ sb_1__4_/top_left_grid_pin_46_
+ sb_1__5_/bottom_left_grid_pin_46_ sb_1__4_/top_left_grid_pin_47_ sb_1__5_/bottom_left_grid_pin_47_
+ sb_1__4_/top_left_grid_pin_48_ sb_1__5_/bottom_left_grid_pin_48_ sb_1__4_/top_left_grid_pin_49_
+ sb_1__5_/bottom_left_grid_pin_49_ cbx_1__5_/bottom_grid_pin_0_ cbx_1__5_/bottom_grid_pin_10_
+ cbx_1__5_/bottom_grid_pin_11_ cbx_1__5_/bottom_grid_pin_12_ cbx_1__5_/bottom_grid_pin_13_
+ cbx_1__5_/bottom_grid_pin_14_ cbx_1__5_/bottom_grid_pin_15_ cbx_1__5_/bottom_grid_pin_1_
+ cbx_1__5_/bottom_grid_pin_2_ cbx_1__5_/REGOUT_FEEDTHROUGH grid_clb_1__5_/top_width_0_height_0__pin_33_
+ sb_1__5_/left_bottom_grid_pin_34_ sb_0__5_/right_bottom_grid_pin_34_ sb_1__5_/left_bottom_grid_pin_35_
+ sb_0__5_/right_bottom_grid_pin_35_ sb_1__5_/left_bottom_grid_pin_36_ sb_0__5_/right_bottom_grid_pin_36_
+ sb_1__5_/left_bottom_grid_pin_37_ sb_0__5_/right_bottom_grid_pin_37_ sb_1__5_/left_bottom_grid_pin_38_
+ sb_0__5_/right_bottom_grid_pin_38_ sb_1__5_/left_bottom_grid_pin_39_ sb_0__5_/right_bottom_grid_pin_39_
+ cbx_1__5_/bottom_grid_pin_3_ sb_1__5_/left_bottom_grid_pin_40_ sb_0__5_/right_bottom_grid_pin_40_
+ sb_1__5_/left_bottom_grid_pin_41_ sb_0__5_/right_bottom_grid_pin_41_ cbx_1__5_/bottom_grid_pin_4_
+ cbx_1__5_/bottom_grid_pin_5_ cbx_1__5_/bottom_grid_pin_6_ cbx_1__5_/bottom_grid_pin_7_
+ cbx_1__5_/bottom_grid_pin_8_ cbx_1__5_/bottom_grid_pin_9_ grid_clb
Xsb_6__2_ sb_6__2_/Test_en_N_out sb_6__2_/Test_en_S_in VGND VPWR sb_6__2_/bottom_left_grid_pin_42_
+ sb_6__2_/bottom_left_grid_pin_43_ sb_6__2_/bottom_left_grid_pin_44_ sb_6__2_/bottom_left_grid_pin_45_
+ sb_6__2_/bottom_left_grid_pin_46_ sb_6__2_/bottom_left_grid_pin_47_ sb_6__2_/bottom_left_grid_pin_48_
+ sb_6__2_/bottom_left_grid_pin_49_ sb_6__2_/ccff_head sb_6__2_/ccff_tail sb_6__2_/chanx_left_in[0]
+ sb_6__2_/chanx_left_in[10] sb_6__2_/chanx_left_in[11] sb_6__2_/chanx_left_in[12]
+ sb_6__2_/chanx_left_in[13] sb_6__2_/chanx_left_in[14] sb_6__2_/chanx_left_in[15]
+ sb_6__2_/chanx_left_in[16] sb_6__2_/chanx_left_in[17] sb_6__2_/chanx_left_in[18]
+ sb_6__2_/chanx_left_in[19] sb_6__2_/chanx_left_in[1] sb_6__2_/chanx_left_in[2] sb_6__2_/chanx_left_in[3]
+ sb_6__2_/chanx_left_in[4] sb_6__2_/chanx_left_in[5] sb_6__2_/chanx_left_in[6] sb_6__2_/chanx_left_in[7]
+ sb_6__2_/chanx_left_in[8] sb_6__2_/chanx_left_in[9] sb_6__2_/chanx_left_out[0] sb_6__2_/chanx_left_out[10]
+ sb_6__2_/chanx_left_out[11] sb_6__2_/chanx_left_out[12] sb_6__2_/chanx_left_out[13]
+ sb_6__2_/chanx_left_out[14] sb_6__2_/chanx_left_out[15] sb_6__2_/chanx_left_out[16]
+ sb_6__2_/chanx_left_out[17] sb_6__2_/chanx_left_out[18] sb_6__2_/chanx_left_out[19]
+ sb_6__2_/chanx_left_out[1] sb_6__2_/chanx_left_out[2] sb_6__2_/chanx_left_out[3]
+ sb_6__2_/chanx_left_out[4] sb_6__2_/chanx_left_out[5] sb_6__2_/chanx_left_out[6]
+ sb_6__2_/chanx_left_out[7] sb_6__2_/chanx_left_out[8] sb_6__2_/chanx_left_out[9]
+ sb_6__2_/chanx_right_in[0] sb_6__2_/chanx_right_in[10] sb_6__2_/chanx_right_in[11]
+ sb_6__2_/chanx_right_in[12] sb_6__2_/chanx_right_in[13] sb_6__2_/chanx_right_in[14]
+ sb_6__2_/chanx_right_in[15] sb_6__2_/chanx_right_in[16] sb_6__2_/chanx_right_in[17]
+ sb_6__2_/chanx_right_in[18] sb_6__2_/chanx_right_in[19] sb_6__2_/chanx_right_in[1]
+ sb_6__2_/chanx_right_in[2] sb_6__2_/chanx_right_in[3] sb_6__2_/chanx_right_in[4]
+ sb_6__2_/chanx_right_in[5] sb_6__2_/chanx_right_in[6] sb_6__2_/chanx_right_in[7]
+ sb_6__2_/chanx_right_in[8] sb_6__2_/chanx_right_in[9] cbx_7__2_/chanx_left_in[0]
+ cbx_7__2_/chanx_left_in[10] cbx_7__2_/chanx_left_in[11] cbx_7__2_/chanx_left_in[12]
+ cbx_7__2_/chanx_left_in[13] cbx_7__2_/chanx_left_in[14] cbx_7__2_/chanx_left_in[15]
+ cbx_7__2_/chanx_left_in[16] cbx_7__2_/chanx_left_in[17] cbx_7__2_/chanx_left_in[18]
+ cbx_7__2_/chanx_left_in[19] cbx_7__2_/chanx_left_in[1] cbx_7__2_/chanx_left_in[2]
+ cbx_7__2_/chanx_left_in[3] cbx_7__2_/chanx_left_in[4] cbx_7__2_/chanx_left_in[5]
+ cbx_7__2_/chanx_left_in[6] cbx_7__2_/chanx_left_in[7] cbx_7__2_/chanx_left_in[8]
+ cbx_7__2_/chanx_left_in[9] cby_6__2_/chany_top_out[0] cby_6__2_/chany_top_out[10]
+ cby_6__2_/chany_top_out[11] cby_6__2_/chany_top_out[12] cby_6__2_/chany_top_out[13]
+ cby_6__2_/chany_top_out[14] cby_6__2_/chany_top_out[15] cby_6__2_/chany_top_out[16]
+ cby_6__2_/chany_top_out[17] cby_6__2_/chany_top_out[18] cby_6__2_/chany_top_out[19]
+ cby_6__2_/chany_top_out[1] cby_6__2_/chany_top_out[2] cby_6__2_/chany_top_out[3]
+ cby_6__2_/chany_top_out[4] cby_6__2_/chany_top_out[5] cby_6__2_/chany_top_out[6]
+ cby_6__2_/chany_top_out[7] cby_6__2_/chany_top_out[8] cby_6__2_/chany_top_out[9]
+ cby_6__2_/chany_top_in[0] cby_6__2_/chany_top_in[10] cby_6__2_/chany_top_in[11]
+ cby_6__2_/chany_top_in[12] cby_6__2_/chany_top_in[13] cby_6__2_/chany_top_in[14]
+ cby_6__2_/chany_top_in[15] cby_6__2_/chany_top_in[16] cby_6__2_/chany_top_in[17]
+ cby_6__2_/chany_top_in[18] cby_6__2_/chany_top_in[19] cby_6__2_/chany_top_in[1]
+ cby_6__2_/chany_top_in[2] cby_6__2_/chany_top_in[3] cby_6__2_/chany_top_in[4] cby_6__2_/chany_top_in[5]
+ cby_6__2_/chany_top_in[6] cby_6__2_/chany_top_in[7] cby_6__2_/chany_top_in[8] cby_6__2_/chany_top_in[9]
+ sb_6__2_/chany_top_in[0] sb_6__2_/chany_top_in[10] sb_6__2_/chany_top_in[11] sb_6__2_/chany_top_in[12]
+ sb_6__2_/chany_top_in[13] sb_6__2_/chany_top_in[14] sb_6__2_/chany_top_in[15] sb_6__2_/chany_top_in[16]
+ sb_6__2_/chany_top_in[17] sb_6__2_/chany_top_in[18] sb_6__2_/chany_top_in[19] sb_6__2_/chany_top_in[1]
+ sb_6__2_/chany_top_in[2] sb_6__2_/chany_top_in[3] sb_6__2_/chany_top_in[4] sb_6__2_/chany_top_in[5]
+ sb_6__2_/chany_top_in[6] sb_6__2_/chany_top_in[7] sb_6__2_/chany_top_in[8] sb_6__2_/chany_top_in[9]
+ sb_6__2_/chany_top_out[0] sb_6__2_/chany_top_out[10] sb_6__2_/chany_top_out[11]
+ sb_6__2_/chany_top_out[12] sb_6__2_/chany_top_out[13] sb_6__2_/chany_top_out[14]
+ sb_6__2_/chany_top_out[15] sb_6__2_/chany_top_out[16] sb_6__2_/chany_top_out[17]
+ sb_6__2_/chany_top_out[18] sb_6__2_/chany_top_out[19] sb_6__2_/chany_top_out[1]
+ sb_6__2_/chany_top_out[2] sb_6__2_/chany_top_out[3] sb_6__2_/chany_top_out[4] sb_6__2_/chany_top_out[5]
+ sb_6__2_/chany_top_out[6] sb_6__2_/chany_top_out[7] sb_6__2_/chany_top_out[8] sb_6__2_/chany_top_out[9]
+ sb_6__2_/clk_1_E_out sb_6__2_/clk_1_N_in sb_6__2_/clk_1_W_out sb_6__2_/clk_2_E_out
+ sb_6__2_/clk_2_N_in sb_6__2_/clk_2_N_out sb_6__2_/clk_2_S_out sb_6__2_/clk_2_W_out
+ sb_6__2_/clk_3_E_out sb_6__2_/clk_3_N_in sb_6__2_/clk_3_N_out sb_6__2_/clk_3_S_out
+ sb_6__2_/clk_3_W_out sb_6__2_/left_bottom_grid_pin_34_ sb_6__2_/left_bottom_grid_pin_35_
+ sb_6__2_/left_bottom_grid_pin_36_ sb_6__2_/left_bottom_grid_pin_37_ sb_6__2_/left_bottom_grid_pin_38_
+ sb_6__2_/left_bottom_grid_pin_39_ sb_6__2_/left_bottom_grid_pin_40_ sb_6__2_/left_bottom_grid_pin_41_
+ sb_6__2_/prog_clk_0_N_in sb_6__2_/prog_clk_1_E_out sb_6__2_/prog_clk_1_N_in sb_6__2_/prog_clk_1_W_out
+ sb_6__2_/prog_clk_2_E_out sb_6__2_/prog_clk_2_N_in sb_6__2_/prog_clk_2_N_out sb_6__2_/prog_clk_2_S_out
+ sb_6__2_/prog_clk_2_W_out sb_6__2_/prog_clk_3_E_out sb_6__2_/prog_clk_3_N_in sb_6__2_/prog_clk_3_N_out
+ sb_6__2_/prog_clk_3_S_out sb_6__2_/prog_clk_3_W_out sb_6__2_/right_bottom_grid_pin_34_
+ sb_6__2_/right_bottom_grid_pin_35_ sb_6__2_/right_bottom_grid_pin_36_ sb_6__2_/right_bottom_grid_pin_37_
+ sb_6__2_/right_bottom_grid_pin_38_ sb_6__2_/right_bottom_grid_pin_39_ sb_6__2_/right_bottom_grid_pin_40_
+ sb_6__2_/right_bottom_grid_pin_41_ sb_6__2_/top_left_grid_pin_42_ sb_6__2_/top_left_grid_pin_43_
+ sb_6__2_/top_left_grid_pin_44_ sb_6__2_/top_left_grid_pin_45_ sb_6__2_/top_left_grid_pin_46_
+ sb_6__2_/top_left_grid_pin_47_ sb_6__2_/top_left_grid_pin_48_ sb_6__2_/top_left_grid_pin_49_
+ sb_1__1_
Xcby_5__6_ cby_5__6_/Test_en_W_in cby_5__6_/Test_en_E_out cby_5__6_/Test_en_N_out
+ cby_5__6_/Test_en_W_in cby_5__6_/Test_en_W_in cby_5__6_/Test_en_W_out VGND VPWR
+ cby_5__6_/ccff_head cby_5__6_/ccff_tail sb_5__5_/chany_top_out[0] sb_5__5_/chany_top_out[10]
+ sb_5__5_/chany_top_out[11] sb_5__5_/chany_top_out[12] sb_5__5_/chany_top_out[13]
+ sb_5__5_/chany_top_out[14] sb_5__5_/chany_top_out[15] sb_5__5_/chany_top_out[16]
+ sb_5__5_/chany_top_out[17] sb_5__5_/chany_top_out[18] sb_5__5_/chany_top_out[19]
+ sb_5__5_/chany_top_out[1] sb_5__5_/chany_top_out[2] sb_5__5_/chany_top_out[3] sb_5__5_/chany_top_out[4]
+ sb_5__5_/chany_top_out[5] sb_5__5_/chany_top_out[6] sb_5__5_/chany_top_out[7] sb_5__5_/chany_top_out[8]
+ sb_5__5_/chany_top_out[9] sb_5__5_/chany_top_in[0] sb_5__5_/chany_top_in[10] sb_5__5_/chany_top_in[11]
+ sb_5__5_/chany_top_in[12] sb_5__5_/chany_top_in[13] sb_5__5_/chany_top_in[14] sb_5__5_/chany_top_in[15]
+ sb_5__5_/chany_top_in[16] sb_5__5_/chany_top_in[17] sb_5__5_/chany_top_in[18] sb_5__5_/chany_top_in[19]
+ sb_5__5_/chany_top_in[1] sb_5__5_/chany_top_in[2] sb_5__5_/chany_top_in[3] sb_5__5_/chany_top_in[4]
+ sb_5__5_/chany_top_in[5] sb_5__5_/chany_top_in[6] sb_5__5_/chany_top_in[7] sb_5__5_/chany_top_in[8]
+ sb_5__5_/chany_top_in[9] cby_5__6_/chany_top_in[0] cby_5__6_/chany_top_in[10] cby_5__6_/chany_top_in[11]
+ cby_5__6_/chany_top_in[12] cby_5__6_/chany_top_in[13] cby_5__6_/chany_top_in[14]
+ cby_5__6_/chany_top_in[15] cby_5__6_/chany_top_in[16] cby_5__6_/chany_top_in[17]
+ cby_5__6_/chany_top_in[18] cby_5__6_/chany_top_in[19] cby_5__6_/chany_top_in[1]
+ cby_5__6_/chany_top_in[2] cby_5__6_/chany_top_in[3] cby_5__6_/chany_top_in[4] cby_5__6_/chany_top_in[5]
+ cby_5__6_/chany_top_in[6] cby_5__6_/chany_top_in[7] cby_5__6_/chany_top_in[8] cby_5__6_/chany_top_in[9]
+ cby_5__6_/chany_top_out[0] cby_5__6_/chany_top_out[10] cby_5__6_/chany_top_out[11]
+ cby_5__6_/chany_top_out[12] cby_5__6_/chany_top_out[13] cby_5__6_/chany_top_out[14]
+ cby_5__6_/chany_top_out[15] cby_5__6_/chany_top_out[16] cby_5__6_/chany_top_out[17]
+ cby_5__6_/chany_top_out[18] cby_5__6_/chany_top_out[19] cby_5__6_/chany_top_out[1]
+ cby_5__6_/chany_top_out[2] cby_5__6_/chany_top_out[3] cby_5__6_/chany_top_out[4]
+ cby_5__6_/chany_top_out[5] cby_5__6_/chany_top_out[6] cby_5__6_/chany_top_out[7]
+ cby_5__6_/chany_top_out[8] cby_5__6_/chany_top_out[9] cby_5__6_/clk_2_N_out sb_5__6_/clk_2_S_out
+ sb_5__5_/clk_1_N_in cby_5__6_/clk_3_N_out cby_5__6_/clk_3_S_in cby_5__6_/clk_3_S_out
+ cby_5__6_/left_grid_pin_16_ cby_5__6_/left_grid_pin_17_ cby_5__6_/left_grid_pin_18_
+ cby_5__6_/left_grid_pin_19_ cby_5__6_/left_grid_pin_20_ cby_5__6_/left_grid_pin_21_
+ cby_5__6_/left_grid_pin_22_ cby_5__6_/left_grid_pin_23_ cby_5__6_/left_grid_pin_24_
+ cby_5__6_/left_grid_pin_25_ cby_5__6_/left_grid_pin_26_ cby_5__6_/left_grid_pin_27_
+ cby_5__6_/left_grid_pin_28_ cby_5__6_/left_grid_pin_29_ cby_5__6_/left_grid_pin_30_
+ cby_5__6_/left_grid_pin_31_ cby_5__6_/prog_clk_0_N_out sb_5__5_/prog_clk_0_N_in
+ cby_5__6_/prog_clk_0_W_in cby_5__6_/prog_clk_2_N_out sb_5__6_/prog_clk_2_S_out sb_5__5_/prog_clk_1_N_in
+ cby_5__6_/prog_clk_3_N_out cby_5__6_/prog_clk_3_S_in cby_5__6_/prog_clk_3_S_out
+ cby_1__1_
Xcby_2__3_ cby_2__3_/Test_en_W_in cby_2__3_/Test_en_E_out cby_2__3_/Test_en_N_out
+ cby_2__3_/Test_en_W_in cby_2__3_/Test_en_W_in cby_2__3_/Test_en_W_out VGND VPWR
+ cby_2__3_/ccff_head cby_2__3_/ccff_tail sb_2__2_/chany_top_out[0] sb_2__2_/chany_top_out[10]
+ sb_2__2_/chany_top_out[11] sb_2__2_/chany_top_out[12] sb_2__2_/chany_top_out[13]
+ sb_2__2_/chany_top_out[14] sb_2__2_/chany_top_out[15] sb_2__2_/chany_top_out[16]
+ sb_2__2_/chany_top_out[17] sb_2__2_/chany_top_out[18] sb_2__2_/chany_top_out[19]
+ sb_2__2_/chany_top_out[1] sb_2__2_/chany_top_out[2] sb_2__2_/chany_top_out[3] sb_2__2_/chany_top_out[4]
+ sb_2__2_/chany_top_out[5] sb_2__2_/chany_top_out[6] sb_2__2_/chany_top_out[7] sb_2__2_/chany_top_out[8]
+ sb_2__2_/chany_top_out[9] sb_2__2_/chany_top_in[0] sb_2__2_/chany_top_in[10] sb_2__2_/chany_top_in[11]
+ sb_2__2_/chany_top_in[12] sb_2__2_/chany_top_in[13] sb_2__2_/chany_top_in[14] sb_2__2_/chany_top_in[15]
+ sb_2__2_/chany_top_in[16] sb_2__2_/chany_top_in[17] sb_2__2_/chany_top_in[18] sb_2__2_/chany_top_in[19]
+ sb_2__2_/chany_top_in[1] sb_2__2_/chany_top_in[2] sb_2__2_/chany_top_in[3] sb_2__2_/chany_top_in[4]
+ sb_2__2_/chany_top_in[5] sb_2__2_/chany_top_in[6] sb_2__2_/chany_top_in[7] sb_2__2_/chany_top_in[8]
+ sb_2__2_/chany_top_in[9] cby_2__3_/chany_top_in[0] cby_2__3_/chany_top_in[10] cby_2__3_/chany_top_in[11]
+ cby_2__3_/chany_top_in[12] cby_2__3_/chany_top_in[13] cby_2__3_/chany_top_in[14]
+ cby_2__3_/chany_top_in[15] cby_2__3_/chany_top_in[16] cby_2__3_/chany_top_in[17]
+ cby_2__3_/chany_top_in[18] cby_2__3_/chany_top_in[19] cby_2__3_/chany_top_in[1]
+ cby_2__3_/chany_top_in[2] cby_2__3_/chany_top_in[3] cby_2__3_/chany_top_in[4] cby_2__3_/chany_top_in[5]
+ cby_2__3_/chany_top_in[6] cby_2__3_/chany_top_in[7] cby_2__3_/chany_top_in[8] cby_2__3_/chany_top_in[9]
+ cby_2__3_/chany_top_out[0] cby_2__3_/chany_top_out[10] cby_2__3_/chany_top_out[11]
+ cby_2__3_/chany_top_out[12] cby_2__3_/chany_top_out[13] cby_2__3_/chany_top_out[14]
+ cby_2__3_/chany_top_out[15] cby_2__3_/chany_top_out[16] cby_2__3_/chany_top_out[17]
+ cby_2__3_/chany_top_out[18] cby_2__3_/chany_top_out[19] cby_2__3_/chany_top_out[1]
+ cby_2__3_/chany_top_out[2] cby_2__3_/chany_top_out[3] cby_2__3_/chany_top_out[4]
+ cby_2__3_/chany_top_out[5] cby_2__3_/chany_top_out[6] cby_2__3_/chany_top_out[7]
+ cby_2__3_/chany_top_out[8] cby_2__3_/chany_top_out[9] cby_2__3_/clk_2_N_out cby_2__3_/clk_2_S_in
+ cby_2__3_/clk_2_S_out cby_2__3_/clk_3_N_out sb_2__3_/clk_3_S_out sb_2__2_/clk_2_N_in
+ cby_2__3_/left_grid_pin_16_ cby_2__3_/left_grid_pin_17_ cby_2__3_/left_grid_pin_18_
+ cby_2__3_/left_grid_pin_19_ cby_2__3_/left_grid_pin_20_ cby_2__3_/left_grid_pin_21_
+ cby_2__3_/left_grid_pin_22_ cby_2__3_/left_grid_pin_23_ cby_2__3_/left_grid_pin_24_
+ cby_2__3_/left_grid_pin_25_ cby_2__3_/left_grid_pin_26_ cby_2__3_/left_grid_pin_27_
+ cby_2__3_/left_grid_pin_28_ cby_2__3_/left_grid_pin_29_ cby_2__3_/left_grid_pin_30_
+ cby_2__3_/left_grid_pin_31_ cby_2__3_/prog_clk_0_N_out sb_2__2_/prog_clk_0_N_in
+ cby_2__3_/prog_clk_0_W_in cby_2__3_/prog_clk_2_N_out cby_2__3_/prog_clk_2_S_in cby_2__3_/prog_clk_2_S_out
+ cby_2__3_/prog_clk_3_N_out sb_2__3_/prog_clk_3_S_out sb_2__2_/prog_clk_2_N_in cby_1__1_
Xcbx_5__7_ cbx_5__7_/REGIN_FEEDTHROUGH cbx_5__7_/REGOUT_FEEDTHROUGH cbx_5__7_/SC_IN_BOT
+ cbx_5__7_/SC_IN_TOP cbx_5__7_/SC_OUT_BOT cbx_5__7_/SC_OUT_TOP VGND VPWR cbx_5__7_/bottom_grid_pin_0_
+ cbx_5__7_/bottom_grid_pin_10_ cbx_5__7_/bottom_grid_pin_11_ cbx_5__7_/bottom_grid_pin_12_
+ cbx_5__7_/bottom_grid_pin_13_ cbx_5__7_/bottom_grid_pin_14_ cbx_5__7_/bottom_grid_pin_15_
+ cbx_5__7_/bottom_grid_pin_1_ cbx_5__7_/bottom_grid_pin_2_ cbx_5__7_/bottom_grid_pin_3_
+ cbx_5__7_/bottom_grid_pin_4_ cbx_5__7_/bottom_grid_pin_5_ cbx_5__7_/bottom_grid_pin_6_
+ cbx_5__7_/bottom_grid_pin_7_ cbx_5__7_/bottom_grid_pin_8_ cbx_5__7_/bottom_grid_pin_9_
+ sb_5__7_/ccff_tail sb_4__7_/ccff_head cbx_5__7_/chanx_left_in[0] cbx_5__7_/chanx_left_in[10]
+ cbx_5__7_/chanx_left_in[11] cbx_5__7_/chanx_left_in[12] cbx_5__7_/chanx_left_in[13]
+ cbx_5__7_/chanx_left_in[14] cbx_5__7_/chanx_left_in[15] cbx_5__7_/chanx_left_in[16]
+ cbx_5__7_/chanx_left_in[17] cbx_5__7_/chanx_left_in[18] cbx_5__7_/chanx_left_in[19]
+ cbx_5__7_/chanx_left_in[1] cbx_5__7_/chanx_left_in[2] cbx_5__7_/chanx_left_in[3]
+ cbx_5__7_/chanx_left_in[4] cbx_5__7_/chanx_left_in[5] cbx_5__7_/chanx_left_in[6]
+ cbx_5__7_/chanx_left_in[7] cbx_5__7_/chanx_left_in[8] cbx_5__7_/chanx_left_in[9]
+ sb_4__7_/chanx_right_in[0] sb_4__7_/chanx_right_in[10] sb_4__7_/chanx_right_in[11]
+ sb_4__7_/chanx_right_in[12] sb_4__7_/chanx_right_in[13] sb_4__7_/chanx_right_in[14]
+ sb_4__7_/chanx_right_in[15] sb_4__7_/chanx_right_in[16] sb_4__7_/chanx_right_in[17]
+ sb_4__7_/chanx_right_in[18] sb_4__7_/chanx_right_in[19] sb_4__7_/chanx_right_in[1]
+ sb_4__7_/chanx_right_in[2] sb_4__7_/chanx_right_in[3] sb_4__7_/chanx_right_in[4]
+ sb_4__7_/chanx_right_in[5] sb_4__7_/chanx_right_in[6] sb_4__7_/chanx_right_in[7]
+ sb_4__7_/chanx_right_in[8] sb_4__7_/chanx_right_in[9] sb_5__7_/chanx_left_out[0]
+ sb_5__7_/chanx_left_out[10] sb_5__7_/chanx_left_out[11] sb_5__7_/chanx_left_out[12]
+ sb_5__7_/chanx_left_out[13] sb_5__7_/chanx_left_out[14] sb_5__7_/chanx_left_out[15]
+ sb_5__7_/chanx_left_out[16] sb_5__7_/chanx_left_out[17] sb_5__7_/chanx_left_out[18]
+ sb_5__7_/chanx_left_out[19] sb_5__7_/chanx_left_out[1] sb_5__7_/chanx_left_out[2]
+ sb_5__7_/chanx_left_out[3] sb_5__7_/chanx_left_out[4] sb_5__7_/chanx_left_out[5]
+ sb_5__7_/chanx_left_out[6] sb_5__7_/chanx_left_out[7] sb_5__7_/chanx_left_out[8]
+ sb_5__7_/chanx_left_out[9] sb_5__7_/chanx_left_in[0] sb_5__7_/chanx_left_in[10]
+ sb_5__7_/chanx_left_in[11] sb_5__7_/chanx_left_in[12] sb_5__7_/chanx_left_in[13]
+ sb_5__7_/chanx_left_in[14] sb_5__7_/chanx_left_in[15] sb_5__7_/chanx_left_in[16]
+ sb_5__7_/chanx_left_in[17] sb_5__7_/chanx_left_in[18] sb_5__7_/chanx_left_in[19]
+ sb_5__7_/chanx_left_in[1] sb_5__7_/chanx_left_in[2] sb_5__7_/chanx_left_in[3] sb_5__7_/chanx_left_in[4]
+ sb_5__7_/chanx_left_in[5] sb_5__7_/chanx_left_in[6] sb_5__7_/chanx_left_in[7] sb_5__7_/chanx_left_in[8]
+ sb_5__7_/chanx_left_in[9] cbx_5__7_/clk_1_N_out cbx_5__7_/clk_1_S_out sb_5__7_/clk_1_W_out
+ cbx_5__7_/clk_2_E_out cbx_5__7_/clk_2_W_in cbx_5__7_/clk_2_W_out cbx_5__7_/clk_3_E_out
+ cbx_5__7_/clk_3_W_in cbx_5__7_/clk_3_W_out cbx_5__7_/prog_clk_0_N_in cbx_5__7_/prog_clk_0_W_out
+ cbx_5__7_/prog_clk_1_N_out cbx_5__7_/prog_clk_1_S_out sb_5__7_/prog_clk_1_W_out
+ cbx_5__7_/prog_clk_2_E_out cbx_5__7_/prog_clk_2_W_in cbx_5__7_/prog_clk_2_W_out
+ cbx_5__7_/prog_clk_3_E_out cbx_5__7_/prog_clk_3_W_in cbx_5__7_/prog_clk_3_W_out
+ cbx_1__1_
Xgrid_clb_4__7_ cbx_4__6_/SC_OUT_TOP grid_clb_4__7_/SC_OUT_BOT cbx_4__7_/SC_IN_BOT
+ cby_4__7_/Test_en_W_out grid_clb_4__7_/Test_en_E_out cby_4__7_/Test_en_W_out cby_3__7_/Test_en_W_in
+ VGND VPWR cbx_4__6_/REGIN_FEEDTHROUGH grid_clb_4__7_/bottom_width_0_height_0__pin_51_
+ cby_3__7_/ccff_tail cby_4__7_/ccff_head cbx_4__7_/clk_1_S_out cbx_4__7_/clk_1_S_out
+ cby_4__7_/prog_clk_0_W_in cbx_4__7_/prog_clk_1_S_out grid_clb_4__7_/prog_clk_0_N_out
+ cbx_4__7_/prog_clk_1_S_out cbx_4__6_/prog_clk_0_N_in grid_clb_4__7_/prog_clk_0_W_out
+ cby_4__7_/left_grid_pin_16_ cby_4__7_/left_grid_pin_17_ cby_4__7_/left_grid_pin_18_
+ cby_4__7_/left_grid_pin_19_ cby_4__7_/left_grid_pin_20_ cby_4__7_/left_grid_pin_21_
+ cby_4__7_/left_grid_pin_22_ cby_4__7_/left_grid_pin_23_ cby_4__7_/left_grid_pin_24_
+ cby_4__7_/left_grid_pin_25_ cby_4__7_/left_grid_pin_26_ cby_4__7_/left_grid_pin_27_
+ cby_4__7_/left_grid_pin_28_ cby_4__7_/left_grid_pin_29_ cby_4__7_/left_grid_pin_30_
+ cby_4__7_/left_grid_pin_31_ sb_4__6_/top_left_grid_pin_42_ sb_4__7_/bottom_left_grid_pin_42_
+ sb_4__6_/top_left_grid_pin_43_ sb_4__7_/bottom_left_grid_pin_43_ sb_4__6_/top_left_grid_pin_44_
+ sb_4__7_/bottom_left_grid_pin_44_ sb_4__6_/top_left_grid_pin_45_ sb_4__7_/bottom_left_grid_pin_45_
+ sb_4__6_/top_left_grid_pin_46_ sb_4__7_/bottom_left_grid_pin_46_ sb_4__6_/top_left_grid_pin_47_
+ sb_4__7_/bottom_left_grid_pin_47_ sb_4__6_/top_left_grid_pin_48_ sb_4__7_/bottom_left_grid_pin_48_
+ sb_4__6_/top_left_grid_pin_49_ sb_4__7_/bottom_left_grid_pin_49_ cbx_4__7_/bottom_grid_pin_0_
+ cbx_4__7_/bottom_grid_pin_10_ cbx_4__7_/bottom_grid_pin_11_ cbx_4__7_/bottom_grid_pin_12_
+ cbx_4__7_/bottom_grid_pin_13_ cbx_4__7_/bottom_grid_pin_14_ cbx_4__7_/bottom_grid_pin_15_
+ cbx_4__7_/bottom_grid_pin_1_ cbx_4__7_/bottom_grid_pin_2_ cbx_4__7_/REGOUT_FEEDTHROUGH
+ grid_clb_4__7_/top_width_0_height_0__pin_33_ sb_4__7_/left_bottom_grid_pin_34_ sb_3__7_/right_bottom_grid_pin_34_
+ sb_4__7_/left_bottom_grid_pin_35_ sb_3__7_/right_bottom_grid_pin_35_ sb_4__7_/left_bottom_grid_pin_36_
+ sb_3__7_/right_bottom_grid_pin_36_ sb_4__7_/left_bottom_grid_pin_37_ sb_3__7_/right_bottom_grid_pin_37_
+ sb_4__7_/left_bottom_grid_pin_38_ sb_3__7_/right_bottom_grid_pin_38_ sb_4__7_/left_bottom_grid_pin_39_
+ sb_3__7_/right_bottom_grid_pin_39_ cbx_4__7_/bottom_grid_pin_3_ sb_4__7_/left_bottom_grid_pin_40_
+ sb_3__7_/right_bottom_grid_pin_40_ sb_4__7_/left_bottom_grid_pin_41_ sb_3__7_/right_bottom_grid_pin_41_
+ cbx_4__7_/bottom_grid_pin_4_ cbx_4__7_/bottom_grid_pin_5_ cbx_4__7_/bottom_grid_pin_6_
+ cbx_4__7_/bottom_grid_pin_7_ cbx_4__7_/bottom_grid_pin_8_ cbx_4__7_/bottom_grid_pin_9_
+ grid_clb
Xcbx_2__4_ cbx_2__4_/REGIN_FEEDTHROUGH cbx_2__4_/REGOUT_FEEDTHROUGH cbx_2__4_/SC_IN_BOT
+ cbx_2__4_/SC_IN_TOP cbx_2__4_/SC_OUT_BOT cbx_2__4_/SC_OUT_TOP VGND VPWR cbx_2__4_/bottom_grid_pin_0_
+ cbx_2__4_/bottom_grid_pin_10_ cbx_2__4_/bottom_grid_pin_11_ cbx_2__4_/bottom_grid_pin_12_
+ cbx_2__4_/bottom_grid_pin_13_ cbx_2__4_/bottom_grid_pin_14_ cbx_2__4_/bottom_grid_pin_15_
+ cbx_2__4_/bottom_grid_pin_1_ cbx_2__4_/bottom_grid_pin_2_ cbx_2__4_/bottom_grid_pin_3_
+ cbx_2__4_/bottom_grid_pin_4_ cbx_2__4_/bottom_grid_pin_5_ cbx_2__4_/bottom_grid_pin_6_
+ cbx_2__4_/bottom_grid_pin_7_ cbx_2__4_/bottom_grid_pin_8_ cbx_2__4_/bottom_grid_pin_9_
+ sb_2__4_/ccff_tail sb_1__4_/ccff_head cbx_2__4_/chanx_left_in[0] cbx_2__4_/chanx_left_in[10]
+ cbx_2__4_/chanx_left_in[11] cbx_2__4_/chanx_left_in[12] cbx_2__4_/chanx_left_in[13]
+ cbx_2__4_/chanx_left_in[14] cbx_2__4_/chanx_left_in[15] cbx_2__4_/chanx_left_in[16]
+ cbx_2__4_/chanx_left_in[17] cbx_2__4_/chanx_left_in[18] cbx_2__4_/chanx_left_in[19]
+ cbx_2__4_/chanx_left_in[1] cbx_2__4_/chanx_left_in[2] cbx_2__4_/chanx_left_in[3]
+ cbx_2__4_/chanx_left_in[4] cbx_2__4_/chanx_left_in[5] cbx_2__4_/chanx_left_in[6]
+ cbx_2__4_/chanx_left_in[7] cbx_2__4_/chanx_left_in[8] cbx_2__4_/chanx_left_in[9]
+ sb_1__4_/chanx_right_in[0] sb_1__4_/chanx_right_in[10] sb_1__4_/chanx_right_in[11]
+ sb_1__4_/chanx_right_in[12] sb_1__4_/chanx_right_in[13] sb_1__4_/chanx_right_in[14]
+ sb_1__4_/chanx_right_in[15] sb_1__4_/chanx_right_in[16] sb_1__4_/chanx_right_in[17]
+ sb_1__4_/chanx_right_in[18] sb_1__4_/chanx_right_in[19] sb_1__4_/chanx_right_in[1]
+ sb_1__4_/chanx_right_in[2] sb_1__4_/chanx_right_in[3] sb_1__4_/chanx_right_in[4]
+ sb_1__4_/chanx_right_in[5] sb_1__4_/chanx_right_in[6] sb_1__4_/chanx_right_in[7]
+ sb_1__4_/chanx_right_in[8] sb_1__4_/chanx_right_in[9] sb_2__4_/chanx_left_out[0]
+ sb_2__4_/chanx_left_out[10] sb_2__4_/chanx_left_out[11] sb_2__4_/chanx_left_out[12]
+ sb_2__4_/chanx_left_out[13] sb_2__4_/chanx_left_out[14] sb_2__4_/chanx_left_out[15]
+ sb_2__4_/chanx_left_out[16] sb_2__4_/chanx_left_out[17] sb_2__4_/chanx_left_out[18]
+ sb_2__4_/chanx_left_out[19] sb_2__4_/chanx_left_out[1] sb_2__4_/chanx_left_out[2]
+ sb_2__4_/chanx_left_out[3] sb_2__4_/chanx_left_out[4] sb_2__4_/chanx_left_out[5]
+ sb_2__4_/chanx_left_out[6] sb_2__4_/chanx_left_out[7] sb_2__4_/chanx_left_out[8]
+ sb_2__4_/chanx_left_out[9] sb_2__4_/chanx_left_in[0] sb_2__4_/chanx_left_in[10]
+ sb_2__4_/chanx_left_in[11] sb_2__4_/chanx_left_in[12] sb_2__4_/chanx_left_in[13]
+ sb_2__4_/chanx_left_in[14] sb_2__4_/chanx_left_in[15] sb_2__4_/chanx_left_in[16]
+ sb_2__4_/chanx_left_in[17] sb_2__4_/chanx_left_in[18] sb_2__4_/chanx_left_in[19]
+ sb_2__4_/chanx_left_in[1] sb_2__4_/chanx_left_in[2] sb_2__4_/chanx_left_in[3] sb_2__4_/chanx_left_in[4]
+ sb_2__4_/chanx_left_in[5] sb_2__4_/chanx_left_in[6] sb_2__4_/chanx_left_in[7] sb_2__4_/chanx_left_in[8]
+ sb_2__4_/chanx_left_in[9] cbx_2__4_/clk_1_N_out cbx_2__4_/clk_1_S_out cbx_2__4_/clk_1_W_in
+ cbx_2__4_/clk_2_E_out cbx_2__4_/clk_2_W_in cbx_2__4_/clk_2_W_out cbx_2__4_/clk_3_E_out
+ cbx_2__4_/clk_3_W_in cbx_2__4_/clk_3_W_out cbx_2__4_/prog_clk_0_N_in cbx_2__4_/prog_clk_0_W_out
+ cbx_2__4_/prog_clk_1_N_out cbx_2__4_/prog_clk_1_S_out cbx_2__4_/prog_clk_1_W_in
+ cbx_2__4_/prog_clk_2_E_out cbx_2__4_/prog_clk_2_W_in cbx_2__4_/prog_clk_2_W_out
+ cbx_2__4_/prog_clk_3_E_out cbx_2__4_/prog_clk_3_W_in cbx_2__4_/prog_clk_3_W_out
+ cbx_1__1_
Xsb_6__1_ sb_6__1_/Test_en_N_out sb_6__1_/Test_en_S_in VGND VPWR sb_6__1_/bottom_left_grid_pin_42_
+ sb_6__1_/bottom_left_grid_pin_43_ sb_6__1_/bottom_left_grid_pin_44_ sb_6__1_/bottom_left_grid_pin_45_
+ sb_6__1_/bottom_left_grid_pin_46_ sb_6__1_/bottom_left_grid_pin_47_ sb_6__1_/bottom_left_grid_pin_48_
+ sb_6__1_/bottom_left_grid_pin_49_ sb_6__1_/ccff_head sb_6__1_/ccff_tail sb_6__1_/chanx_left_in[0]
+ sb_6__1_/chanx_left_in[10] sb_6__1_/chanx_left_in[11] sb_6__1_/chanx_left_in[12]
+ sb_6__1_/chanx_left_in[13] sb_6__1_/chanx_left_in[14] sb_6__1_/chanx_left_in[15]
+ sb_6__1_/chanx_left_in[16] sb_6__1_/chanx_left_in[17] sb_6__1_/chanx_left_in[18]
+ sb_6__1_/chanx_left_in[19] sb_6__1_/chanx_left_in[1] sb_6__1_/chanx_left_in[2] sb_6__1_/chanx_left_in[3]
+ sb_6__1_/chanx_left_in[4] sb_6__1_/chanx_left_in[5] sb_6__1_/chanx_left_in[6] sb_6__1_/chanx_left_in[7]
+ sb_6__1_/chanx_left_in[8] sb_6__1_/chanx_left_in[9] sb_6__1_/chanx_left_out[0] sb_6__1_/chanx_left_out[10]
+ sb_6__1_/chanx_left_out[11] sb_6__1_/chanx_left_out[12] sb_6__1_/chanx_left_out[13]
+ sb_6__1_/chanx_left_out[14] sb_6__1_/chanx_left_out[15] sb_6__1_/chanx_left_out[16]
+ sb_6__1_/chanx_left_out[17] sb_6__1_/chanx_left_out[18] sb_6__1_/chanx_left_out[19]
+ sb_6__1_/chanx_left_out[1] sb_6__1_/chanx_left_out[2] sb_6__1_/chanx_left_out[3]
+ sb_6__1_/chanx_left_out[4] sb_6__1_/chanx_left_out[5] sb_6__1_/chanx_left_out[6]
+ sb_6__1_/chanx_left_out[7] sb_6__1_/chanx_left_out[8] sb_6__1_/chanx_left_out[9]
+ sb_6__1_/chanx_right_in[0] sb_6__1_/chanx_right_in[10] sb_6__1_/chanx_right_in[11]
+ sb_6__1_/chanx_right_in[12] sb_6__1_/chanx_right_in[13] sb_6__1_/chanx_right_in[14]
+ sb_6__1_/chanx_right_in[15] sb_6__1_/chanx_right_in[16] sb_6__1_/chanx_right_in[17]
+ sb_6__1_/chanx_right_in[18] sb_6__1_/chanx_right_in[19] sb_6__1_/chanx_right_in[1]
+ sb_6__1_/chanx_right_in[2] sb_6__1_/chanx_right_in[3] sb_6__1_/chanx_right_in[4]
+ sb_6__1_/chanx_right_in[5] sb_6__1_/chanx_right_in[6] sb_6__1_/chanx_right_in[7]
+ sb_6__1_/chanx_right_in[8] sb_6__1_/chanx_right_in[9] cbx_7__1_/chanx_left_in[0]
+ cbx_7__1_/chanx_left_in[10] cbx_7__1_/chanx_left_in[11] cbx_7__1_/chanx_left_in[12]
+ cbx_7__1_/chanx_left_in[13] cbx_7__1_/chanx_left_in[14] cbx_7__1_/chanx_left_in[15]
+ cbx_7__1_/chanx_left_in[16] cbx_7__1_/chanx_left_in[17] cbx_7__1_/chanx_left_in[18]
+ cbx_7__1_/chanx_left_in[19] cbx_7__1_/chanx_left_in[1] cbx_7__1_/chanx_left_in[2]
+ cbx_7__1_/chanx_left_in[3] cbx_7__1_/chanx_left_in[4] cbx_7__1_/chanx_left_in[5]
+ cbx_7__1_/chanx_left_in[6] cbx_7__1_/chanx_left_in[7] cbx_7__1_/chanx_left_in[8]
+ cbx_7__1_/chanx_left_in[9] cby_6__1_/chany_top_out[0] cby_6__1_/chany_top_out[10]
+ cby_6__1_/chany_top_out[11] cby_6__1_/chany_top_out[12] cby_6__1_/chany_top_out[13]
+ cby_6__1_/chany_top_out[14] cby_6__1_/chany_top_out[15] cby_6__1_/chany_top_out[16]
+ cby_6__1_/chany_top_out[17] cby_6__1_/chany_top_out[18] cby_6__1_/chany_top_out[19]
+ cby_6__1_/chany_top_out[1] cby_6__1_/chany_top_out[2] cby_6__1_/chany_top_out[3]
+ cby_6__1_/chany_top_out[4] cby_6__1_/chany_top_out[5] cby_6__1_/chany_top_out[6]
+ cby_6__1_/chany_top_out[7] cby_6__1_/chany_top_out[8] cby_6__1_/chany_top_out[9]
+ cby_6__1_/chany_top_in[0] cby_6__1_/chany_top_in[10] cby_6__1_/chany_top_in[11]
+ cby_6__1_/chany_top_in[12] cby_6__1_/chany_top_in[13] cby_6__1_/chany_top_in[14]
+ cby_6__1_/chany_top_in[15] cby_6__1_/chany_top_in[16] cby_6__1_/chany_top_in[17]
+ cby_6__1_/chany_top_in[18] cby_6__1_/chany_top_in[19] cby_6__1_/chany_top_in[1]
+ cby_6__1_/chany_top_in[2] cby_6__1_/chany_top_in[3] cby_6__1_/chany_top_in[4] cby_6__1_/chany_top_in[5]
+ cby_6__1_/chany_top_in[6] cby_6__1_/chany_top_in[7] cby_6__1_/chany_top_in[8] cby_6__1_/chany_top_in[9]
+ sb_6__1_/chany_top_in[0] sb_6__1_/chany_top_in[10] sb_6__1_/chany_top_in[11] sb_6__1_/chany_top_in[12]
+ sb_6__1_/chany_top_in[13] sb_6__1_/chany_top_in[14] sb_6__1_/chany_top_in[15] sb_6__1_/chany_top_in[16]
+ sb_6__1_/chany_top_in[17] sb_6__1_/chany_top_in[18] sb_6__1_/chany_top_in[19] sb_6__1_/chany_top_in[1]
+ sb_6__1_/chany_top_in[2] sb_6__1_/chany_top_in[3] sb_6__1_/chany_top_in[4] sb_6__1_/chany_top_in[5]
+ sb_6__1_/chany_top_in[6] sb_6__1_/chany_top_in[7] sb_6__1_/chany_top_in[8] sb_6__1_/chany_top_in[9]
+ sb_6__1_/chany_top_out[0] sb_6__1_/chany_top_out[10] sb_6__1_/chany_top_out[11]
+ sb_6__1_/chany_top_out[12] sb_6__1_/chany_top_out[13] sb_6__1_/chany_top_out[14]
+ sb_6__1_/chany_top_out[15] sb_6__1_/chany_top_out[16] sb_6__1_/chany_top_out[17]
+ sb_6__1_/chany_top_out[18] sb_6__1_/chany_top_out[19] sb_6__1_/chany_top_out[1]
+ sb_6__1_/chany_top_out[2] sb_6__1_/chany_top_out[3] sb_6__1_/chany_top_out[4] sb_6__1_/chany_top_out[5]
+ sb_6__1_/chany_top_out[6] sb_6__1_/chany_top_out[7] sb_6__1_/chany_top_out[8] sb_6__1_/chany_top_out[9]
+ sb_6__1_/clk_1_E_out sb_6__1_/clk_1_N_in sb_6__1_/clk_1_W_out sb_6__1_/clk_2_E_out
+ sb_6__1_/clk_2_N_in sb_6__1_/clk_2_N_out sb_6__1_/clk_2_S_out sb_6__1_/clk_2_W_out
+ sb_6__1_/clk_3_E_out sb_6__1_/clk_3_N_in sb_6__1_/clk_3_N_out sb_6__1_/clk_3_S_out
+ sb_6__1_/clk_3_W_out sb_6__1_/left_bottom_grid_pin_34_ sb_6__1_/left_bottom_grid_pin_35_
+ sb_6__1_/left_bottom_grid_pin_36_ sb_6__1_/left_bottom_grid_pin_37_ sb_6__1_/left_bottom_grid_pin_38_
+ sb_6__1_/left_bottom_grid_pin_39_ sb_6__1_/left_bottom_grid_pin_40_ sb_6__1_/left_bottom_grid_pin_41_
+ sb_6__1_/prog_clk_0_N_in sb_6__1_/prog_clk_1_E_out sb_6__1_/prog_clk_1_N_in sb_6__1_/prog_clk_1_W_out
+ sb_6__1_/prog_clk_2_E_out sb_6__1_/prog_clk_2_N_in sb_6__1_/prog_clk_2_N_out sb_6__1_/prog_clk_2_S_out
+ sb_6__1_/prog_clk_2_W_out sb_6__1_/prog_clk_3_E_out sb_6__1_/prog_clk_3_N_in sb_6__1_/prog_clk_3_N_out
+ sb_6__1_/prog_clk_3_S_out sb_6__1_/prog_clk_3_W_out sb_6__1_/right_bottom_grid_pin_34_
+ sb_6__1_/right_bottom_grid_pin_35_ sb_6__1_/right_bottom_grid_pin_36_ sb_6__1_/right_bottom_grid_pin_37_
+ sb_6__1_/right_bottom_grid_pin_38_ sb_6__1_/right_bottom_grid_pin_39_ sb_6__1_/right_bottom_grid_pin_40_
+ sb_6__1_/right_bottom_grid_pin_41_ sb_6__1_/top_left_grid_pin_42_ sb_6__1_/top_left_grid_pin_43_
+ sb_6__1_/top_left_grid_pin_44_ sb_6__1_/top_left_grid_pin_45_ sb_6__1_/top_left_grid_pin_46_
+ sb_6__1_/top_left_grid_pin_47_ sb_6__1_/top_left_grid_pin_48_ sb_6__1_/top_left_grid_pin_49_
+ sb_1__1_
Xgrid_clb_1__4_ cbx_1__4_/SC_OUT_BOT cbx_1__3_/SC_IN_TOP grid_clb_1__4_/SC_OUT_TOP
+ cby_1__4_/Test_en_W_out grid_clb_1__4_/Test_en_E_out cby_1__4_/Test_en_W_out grid_clb_1__4_/Test_en_W_out
+ VGND VPWR cbx_1__3_/REGIN_FEEDTHROUGH grid_clb_1__4_/bottom_width_0_height_0__pin_51_
+ cby_0__4_/ccff_tail cby_1__4_/ccff_head cbx_1__3_/clk_1_N_out cbx_1__3_/clk_1_N_out
+ cby_1__4_/prog_clk_0_W_in cbx_1__3_/prog_clk_1_N_out grid_clb_1__4_/prog_clk_0_N_out
+ cbx_1__3_/prog_clk_1_N_out cbx_1__3_/prog_clk_0_N_in cby_0__4_/prog_clk_0_E_in cby_1__4_/left_grid_pin_16_
+ cby_1__4_/left_grid_pin_17_ cby_1__4_/left_grid_pin_18_ cby_1__4_/left_grid_pin_19_
+ cby_1__4_/left_grid_pin_20_ cby_1__4_/left_grid_pin_21_ cby_1__4_/left_grid_pin_22_
+ cby_1__4_/left_grid_pin_23_ cby_1__4_/left_grid_pin_24_ cby_1__4_/left_grid_pin_25_
+ cby_1__4_/left_grid_pin_26_ cby_1__4_/left_grid_pin_27_ cby_1__4_/left_grid_pin_28_
+ cby_1__4_/left_grid_pin_29_ cby_1__4_/left_grid_pin_30_ cby_1__4_/left_grid_pin_31_
+ sb_1__3_/top_left_grid_pin_42_ sb_1__4_/bottom_left_grid_pin_42_ sb_1__3_/top_left_grid_pin_43_
+ sb_1__4_/bottom_left_grid_pin_43_ sb_1__3_/top_left_grid_pin_44_ sb_1__4_/bottom_left_grid_pin_44_
+ sb_1__3_/top_left_grid_pin_45_ sb_1__4_/bottom_left_grid_pin_45_ sb_1__3_/top_left_grid_pin_46_
+ sb_1__4_/bottom_left_grid_pin_46_ sb_1__3_/top_left_grid_pin_47_ sb_1__4_/bottom_left_grid_pin_47_
+ sb_1__3_/top_left_grid_pin_48_ sb_1__4_/bottom_left_grid_pin_48_ sb_1__3_/top_left_grid_pin_49_
+ sb_1__4_/bottom_left_grid_pin_49_ cbx_1__4_/bottom_grid_pin_0_ cbx_1__4_/bottom_grid_pin_10_
+ cbx_1__4_/bottom_grid_pin_11_ cbx_1__4_/bottom_grid_pin_12_ cbx_1__4_/bottom_grid_pin_13_
+ cbx_1__4_/bottom_grid_pin_14_ cbx_1__4_/bottom_grid_pin_15_ cbx_1__4_/bottom_grid_pin_1_
+ cbx_1__4_/bottom_grid_pin_2_ cbx_1__4_/REGOUT_FEEDTHROUGH grid_clb_1__4_/top_width_0_height_0__pin_33_
+ sb_1__4_/left_bottom_grid_pin_34_ sb_0__4_/right_bottom_grid_pin_34_ sb_1__4_/left_bottom_grid_pin_35_
+ sb_0__4_/right_bottom_grid_pin_35_ sb_1__4_/left_bottom_grid_pin_36_ sb_0__4_/right_bottom_grid_pin_36_
+ sb_1__4_/left_bottom_grid_pin_37_ sb_0__4_/right_bottom_grid_pin_37_ sb_1__4_/left_bottom_grid_pin_38_
+ sb_0__4_/right_bottom_grid_pin_38_ sb_1__4_/left_bottom_grid_pin_39_ sb_0__4_/right_bottom_grid_pin_39_
+ cbx_1__4_/bottom_grid_pin_3_ sb_1__4_/left_bottom_grid_pin_40_ sb_0__4_/right_bottom_grid_pin_40_
+ sb_1__4_/left_bottom_grid_pin_41_ sb_0__4_/right_bottom_grid_pin_41_ cbx_1__4_/bottom_grid_pin_4_
+ cbx_1__4_/bottom_grid_pin_5_ cbx_1__4_/bottom_grid_pin_6_ cbx_1__4_/bottom_grid_pin_7_
+ cbx_1__4_/bottom_grid_pin_8_ cbx_1__4_/bottom_grid_pin_9_ grid_clb
Xcby_8__8_ IO_ISOL_N VGND VPWR cby_8__8_/ccff_head sb_8__7_/ccff_head sb_8__7_/chany_top_out[0]
+ sb_8__7_/chany_top_out[10] sb_8__7_/chany_top_out[11] sb_8__7_/chany_top_out[12]
+ sb_8__7_/chany_top_out[13] sb_8__7_/chany_top_out[14] sb_8__7_/chany_top_out[15]
+ sb_8__7_/chany_top_out[16] sb_8__7_/chany_top_out[17] sb_8__7_/chany_top_out[18]
+ sb_8__7_/chany_top_out[19] sb_8__7_/chany_top_out[1] sb_8__7_/chany_top_out[2] sb_8__7_/chany_top_out[3]
+ sb_8__7_/chany_top_out[4] sb_8__7_/chany_top_out[5] sb_8__7_/chany_top_out[6] sb_8__7_/chany_top_out[7]
+ sb_8__7_/chany_top_out[8] sb_8__7_/chany_top_out[9] sb_8__7_/chany_top_in[0] sb_8__7_/chany_top_in[10]
+ sb_8__7_/chany_top_in[11] sb_8__7_/chany_top_in[12] sb_8__7_/chany_top_in[13] sb_8__7_/chany_top_in[14]
+ sb_8__7_/chany_top_in[15] sb_8__7_/chany_top_in[16] sb_8__7_/chany_top_in[17] sb_8__7_/chany_top_in[18]
+ sb_8__7_/chany_top_in[19] sb_8__7_/chany_top_in[1] sb_8__7_/chany_top_in[2] sb_8__7_/chany_top_in[3]
+ sb_8__7_/chany_top_in[4] sb_8__7_/chany_top_in[5] sb_8__7_/chany_top_in[6] sb_8__7_/chany_top_in[7]
+ sb_8__7_/chany_top_in[8] sb_8__7_/chany_top_in[9] cby_8__8_/chany_top_in[0] cby_8__8_/chany_top_in[10]
+ cby_8__8_/chany_top_in[11] cby_8__8_/chany_top_in[12] cby_8__8_/chany_top_in[13]
+ cby_8__8_/chany_top_in[14] cby_8__8_/chany_top_in[15] cby_8__8_/chany_top_in[16]
+ cby_8__8_/chany_top_in[17] cby_8__8_/chany_top_in[18] cby_8__8_/chany_top_in[19]
+ cby_8__8_/chany_top_in[1] cby_8__8_/chany_top_in[2] cby_8__8_/chany_top_in[3] cby_8__8_/chany_top_in[4]
+ cby_8__8_/chany_top_in[5] cby_8__8_/chany_top_in[6] cby_8__8_/chany_top_in[7] cby_8__8_/chany_top_in[8]
+ cby_8__8_/chany_top_in[9] cby_8__8_/chany_top_out[0] cby_8__8_/chany_top_out[10]
+ cby_8__8_/chany_top_out[11] cby_8__8_/chany_top_out[12] cby_8__8_/chany_top_out[13]
+ cby_8__8_/chany_top_out[14] cby_8__8_/chany_top_out[15] cby_8__8_/chany_top_out[16]
+ cby_8__8_/chany_top_out[17] cby_8__8_/chany_top_out[18] cby_8__8_/chany_top_out[19]
+ cby_8__8_/chany_top_out[1] cby_8__8_/chany_top_out[2] cby_8__8_/chany_top_out[3]
+ cby_8__8_/chany_top_out[4] cby_8__8_/chany_top_out[5] cby_8__8_/chany_top_out[6]
+ cby_8__8_/chany_top_out[7] cby_8__8_/chany_top_out[8] cby_8__8_/chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
+ cby_8__8_/left_grid_pin_16_ cby_8__8_/left_grid_pin_17_ cby_8__8_/left_grid_pin_18_
+ cby_8__8_/left_grid_pin_19_ cby_8__8_/left_grid_pin_20_ cby_8__8_/left_grid_pin_21_
+ cby_8__8_/left_grid_pin_22_ cby_8__8_/left_grid_pin_23_ cby_8__8_/left_grid_pin_24_
+ cby_8__8_/left_grid_pin_25_ cby_8__8_/left_grid_pin_26_ cby_8__8_/left_grid_pin_27_
+ cby_8__8_/left_grid_pin_28_ cby_8__8_/left_grid_pin_29_ cby_8__8_/left_grid_pin_30_
+ cby_8__8_/left_grid_pin_31_ cby_8__8_/right_grid_pin_0_ sb_8__7_/top_right_grid_pin_1_
+ sb_8__8_/bottom_right_grid_pin_1_ sb_8__8_/prog_clk_0_S_in sb_8__7_/prog_clk_0_N_in
+ cby_8__8_/prog_clk_0_W_in cby_8__8_/right_grid_pin_0_ cby_2__1_
Xcby_5__5_ cby_5__5_/Test_en_W_in cby_5__5_/Test_en_E_out cby_5__5_/Test_en_N_out
+ cby_5__5_/Test_en_W_in cby_5__5_/Test_en_W_in cby_5__5_/Test_en_W_out VGND VPWR
+ cby_5__5_/ccff_head cby_5__5_/ccff_tail sb_5__4_/chany_top_out[0] sb_5__4_/chany_top_out[10]
+ sb_5__4_/chany_top_out[11] sb_5__4_/chany_top_out[12] sb_5__4_/chany_top_out[13]
+ sb_5__4_/chany_top_out[14] sb_5__4_/chany_top_out[15] sb_5__4_/chany_top_out[16]
+ sb_5__4_/chany_top_out[17] sb_5__4_/chany_top_out[18] sb_5__4_/chany_top_out[19]
+ sb_5__4_/chany_top_out[1] sb_5__4_/chany_top_out[2] sb_5__4_/chany_top_out[3] sb_5__4_/chany_top_out[4]
+ sb_5__4_/chany_top_out[5] sb_5__4_/chany_top_out[6] sb_5__4_/chany_top_out[7] sb_5__4_/chany_top_out[8]
+ sb_5__4_/chany_top_out[9] sb_5__4_/chany_top_in[0] sb_5__4_/chany_top_in[10] sb_5__4_/chany_top_in[11]
+ sb_5__4_/chany_top_in[12] sb_5__4_/chany_top_in[13] sb_5__4_/chany_top_in[14] sb_5__4_/chany_top_in[15]
+ sb_5__4_/chany_top_in[16] sb_5__4_/chany_top_in[17] sb_5__4_/chany_top_in[18] sb_5__4_/chany_top_in[19]
+ sb_5__4_/chany_top_in[1] sb_5__4_/chany_top_in[2] sb_5__4_/chany_top_in[3] sb_5__4_/chany_top_in[4]
+ sb_5__4_/chany_top_in[5] sb_5__4_/chany_top_in[6] sb_5__4_/chany_top_in[7] sb_5__4_/chany_top_in[8]
+ sb_5__4_/chany_top_in[9] cby_5__5_/chany_top_in[0] cby_5__5_/chany_top_in[10] cby_5__5_/chany_top_in[11]
+ cby_5__5_/chany_top_in[12] cby_5__5_/chany_top_in[13] cby_5__5_/chany_top_in[14]
+ cby_5__5_/chany_top_in[15] cby_5__5_/chany_top_in[16] cby_5__5_/chany_top_in[17]
+ cby_5__5_/chany_top_in[18] cby_5__5_/chany_top_in[19] cby_5__5_/chany_top_in[1]
+ cby_5__5_/chany_top_in[2] cby_5__5_/chany_top_in[3] cby_5__5_/chany_top_in[4] cby_5__5_/chany_top_in[5]
+ cby_5__5_/chany_top_in[6] cby_5__5_/chany_top_in[7] cby_5__5_/chany_top_in[8] cby_5__5_/chany_top_in[9]
+ cby_5__5_/chany_top_out[0] cby_5__5_/chany_top_out[10] cby_5__5_/chany_top_out[11]
+ cby_5__5_/chany_top_out[12] cby_5__5_/chany_top_out[13] cby_5__5_/chany_top_out[14]
+ cby_5__5_/chany_top_out[15] cby_5__5_/chany_top_out[16] cby_5__5_/chany_top_out[17]
+ cby_5__5_/chany_top_out[18] cby_5__5_/chany_top_out[19] cby_5__5_/chany_top_out[1]
+ cby_5__5_/chany_top_out[2] cby_5__5_/chany_top_out[3] cby_5__5_/chany_top_out[4]
+ cby_5__5_/chany_top_out[5] cby_5__5_/chany_top_out[6] cby_5__5_/chany_top_out[7]
+ cby_5__5_/chany_top_out[8] cby_5__5_/chany_top_out[9] cby_5__5_/clk_2_N_out cby_5__5_/clk_2_S_in
+ cby_5__5_/clk_2_S_out cby_5__5_/clk_3_N_out cby_5__5_/clk_3_S_in cby_5__5_/clk_3_S_out
+ cby_5__5_/left_grid_pin_16_ cby_5__5_/left_grid_pin_17_ cby_5__5_/left_grid_pin_18_
+ cby_5__5_/left_grid_pin_19_ cby_5__5_/left_grid_pin_20_ cby_5__5_/left_grid_pin_21_
+ cby_5__5_/left_grid_pin_22_ cby_5__5_/left_grid_pin_23_ cby_5__5_/left_grid_pin_24_
+ cby_5__5_/left_grid_pin_25_ cby_5__5_/left_grid_pin_26_ cby_5__5_/left_grid_pin_27_
+ cby_5__5_/left_grid_pin_28_ cby_5__5_/left_grid_pin_29_ cby_5__5_/left_grid_pin_30_
+ cby_5__5_/left_grid_pin_31_ cby_5__5_/prog_clk_0_N_out sb_5__4_/prog_clk_0_N_in
+ cby_5__5_/prog_clk_0_W_in cby_5__5_/prog_clk_2_N_out cby_5__5_/prog_clk_2_S_in cby_5__5_/prog_clk_2_S_out
+ cby_5__5_/prog_clk_3_N_out cby_5__5_/prog_clk_3_S_in cby_5__5_/prog_clk_3_S_out
+ cby_1__1_
.ends

