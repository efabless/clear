magic
tech sky130A
magscale 1 2
timestamp 1681685267
<< viali >>
rect 16405 54281 16439 54315
rect 18981 54281 19015 54315
rect 25329 54213 25363 54247
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9597 54145 9631 54179
rect 12173 54145 12207 54179
rect 14473 54145 14507 54179
rect 15025 54145 15059 54179
rect 15945 54145 15979 54179
rect 16865 54145 16899 54179
rect 17969 54145 18003 54179
rect 19441 54145 19475 54179
rect 20729 54145 20763 54179
rect 21281 54145 21315 54179
rect 22017 54145 22051 54179
rect 22569 54145 22603 54179
rect 23397 54145 23431 54179
rect 24685 54145 24719 54179
rect 2513 54077 2547 54111
rect 5181 54077 5215 54111
rect 7849 54077 7883 54111
rect 9873 54077 9907 54111
rect 12633 54077 12667 54111
rect 19717 54077 19751 54111
rect 23121 54077 23155 54111
rect 22201 54009 22235 54043
rect 14289 53941 14323 53975
rect 15669 53941 15703 53975
rect 17509 53941 17543 53975
rect 18613 53941 18647 53975
rect 20913 53941 20947 53975
rect 24041 53941 24075 53975
rect 13829 53737 13863 53771
rect 14933 53737 14967 53771
rect 18153 53737 18187 53771
rect 2053 53601 2087 53635
rect 4445 53601 4479 53635
rect 7113 53601 7147 53635
rect 11253 53601 11287 53635
rect 1777 53533 1811 53567
rect 4169 53533 4203 53567
rect 6837 53533 6871 53567
rect 10793 53533 10827 53567
rect 14289 53533 14323 53567
rect 15577 53533 15611 53567
rect 17049 53533 17083 53567
rect 17877 53533 17911 53567
rect 22293 53533 22327 53567
rect 23121 53533 23155 53567
rect 23765 53533 23799 53567
rect 24685 53533 24719 53567
rect 15393 53397 15427 53431
rect 16865 53397 16899 53431
rect 17693 53397 17727 53431
rect 22477 53397 22511 53431
rect 23213 53397 23247 53431
rect 23949 53397 23983 53431
rect 25329 53397 25363 53431
rect 5181 53193 5215 53227
rect 23305 53193 23339 53227
rect 23397 53193 23431 53227
rect 25053 53193 25087 53227
rect 25329 53193 25363 53227
rect 5365 53057 5399 53091
rect 23765 53057 23799 53091
rect 24501 53057 24535 53091
rect 22753 52989 22787 53023
rect 25513 52921 25547 52955
rect 23949 52853 23983 52887
rect 24685 52853 24719 52887
rect 6561 52649 6595 52683
rect 24501 52649 24535 52683
rect 23949 52581 23983 52615
rect 6745 52445 6779 52479
rect 23765 52445 23799 52479
rect 25329 52445 25363 52479
rect 24961 52377 24995 52411
rect 24133 52105 24167 52139
rect 24593 51969 24627 52003
rect 25053 51969 25087 52003
rect 24409 51765 24443 51799
rect 25237 51765 25271 51799
rect 8309 51561 8343 51595
rect 9229 51493 9263 51527
rect 7849 51357 7883 51391
rect 8493 51357 8527 51391
rect 9413 51357 9447 51391
rect 7665 51289 7699 51323
rect 24593 51289 24627 51323
rect 24961 51289 24995 51323
rect 25329 51289 25363 51323
rect 24593 50881 24627 50915
rect 24961 50881 24995 50915
rect 25053 50677 25087 50711
rect 7849 50473 7883 50507
rect 9597 50473 9631 50507
rect 8033 50405 8067 50439
rect 8401 50337 8435 50371
rect 7573 50269 7607 50303
rect 24593 50269 24627 50303
rect 9505 50201 9539 50235
rect 25237 50133 25271 50167
rect 23397 49793 23431 49827
rect 24777 49793 24811 49827
rect 24041 49725 24075 49759
rect 24501 49725 24535 49759
rect 24225 49385 24259 49419
rect 10701 49317 10735 49351
rect 11713 49317 11747 49351
rect 24685 49181 24719 49215
rect 10517 49113 10551 49147
rect 11529 49113 11563 49147
rect 25329 49045 25363 49079
rect 24777 48841 24811 48875
rect 25145 48773 25179 48807
rect 6653 48705 6687 48739
rect 6929 48637 6963 48671
rect 8401 48637 8435 48671
rect 8769 48569 8803 48603
rect 25329 48569 25363 48603
rect 8953 48501 8987 48535
rect 10368 48093 10402 48127
rect 23397 48093 23431 48127
rect 24685 48093 24719 48127
rect 10471 47957 10505 47991
rect 24041 47957 24075 47991
rect 25329 47957 25363 47991
rect 9873 47753 9907 47787
rect 24777 47753 24811 47787
rect 10149 47685 10183 47719
rect 25145 47685 25179 47719
rect 9413 47617 9447 47651
rect 25329 47481 25363 47515
rect 9505 47413 9539 47447
rect 25145 47141 25179 47175
rect 11656 47005 11690 47039
rect 24869 47005 24903 47039
rect 25329 47005 25363 47039
rect 11759 46937 11793 46971
rect 10793 46665 10827 46699
rect 11069 46665 11103 46699
rect 14749 46597 14783 46631
rect 14841 46597 14875 46631
rect 10333 46529 10367 46563
rect 12576 46529 12610 46563
rect 24869 46529 24903 46563
rect 25329 46529 25363 46563
rect 15761 46461 15795 46495
rect 10425 46325 10459 46359
rect 12679 46325 12713 46359
rect 25145 46325 25179 46359
rect 8493 46121 8527 46155
rect 8125 45985 8159 46019
rect 15669 45985 15703 46019
rect 16497 45985 16531 46019
rect 7941 45917 7975 45951
rect 13312 45917 13346 45951
rect 24869 45917 24903 45951
rect 25329 45917 25363 45951
rect 15761 45849 15795 45883
rect 13415 45781 13449 45815
rect 25145 45781 25179 45815
rect 13553 45509 13587 45543
rect 13645 45509 13679 45543
rect 24869 45441 24903 45475
rect 25329 45441 25363 45475
rect 14565 45373 14599 45407
rect 25145 45237 25179 45271
rect 10885 45033 10919 45067
rect 16497 44897 16531 44931
rect 9137 44829 9171 44863
rect 9413 44761 9447 44795
rect 11253 44761 11287 44795
rect 16566 44761 16600 44795
rect 17509 44761 17543 44795
rect 25145 44761 25179 44795
rect 11437 44693 11471 44727
rect 25237 44693 25271 44727
rect 9597 44489 9631 44523
rect 25329 44489 25363 44523
rect 9137 44353 9171 44387
rect 10609 44353 10643 44387
rect 11529 44353 11563 44387
rect 24409 44353 24443 44387
rect 24685 44353 24719 44387
rect 8953 44285 8987 44319
rect 10701 44149 10735 44183
rect 11069 44149 11103 44183
rect 20637 43809 20671 43843
rect 20361 43741 20395 43775
rect 20085 43673 20119 43707
rect 25145 43673 25179 43707
rect 22109 43605 22143 43639
rect 25237 43605 25271 43639
rect 25329 43401 25363 43435
rect 24409 43265 24443 43299
rect 24685 43265 24719 43299
rect 10241 42721 10275 42755
rect 9597 42653 9631 42687
rect 9781 42653 9815 42687
rect 24685 42653 24719 42687
rect 25329 42517 25363 42551
rect 11161 42313 11195 42347
rect 24777 42313 24811 42347
rect 25145 42245 25179 42279
rect 9413 42109 9447 42143
rect 9689 42109 9723 42143
rect 11529 41973 11563 42007
rect 11713 41973 11747 42007
rect 25237 41973 25271 42007
rect 10885 41769 10919 41803
rect 10425 41633 10459 41667
rect 10241 41565 10275 41599
rect 24685 41565 24719 41599
rect 25329 41429 25363 41463
rect 24777 41225 24811 41259
rect 25145 41157 25179 41191
rect 25237 40885 25271 40919
rect 24869 40477 24903 40511
rect 25329 40477 25363 40511
rect 25145 40341 25179 40375
rect 25145 40137 25179 40171
rect 24869 40001 24903 40035
rect 25329 40001 25363 40035
rect 24869 39389 24903 39423
rect 25329 39389 25363 39423
rect 25145 39253 25179 39287
rect 25329 38913 25363 38947
rect 24869 38709 24903 38743
rect 25145 38709 25179 38743
rect 25145 38233 25179 38267
rect 25237 38165 25271 38199
rect 8677 37961 8711 37995
rect 25329 37961 25363 37995
rect 8861 37825 8895 37859
rect 24409 37825 24443 37859
rect 24685 37825 24719 37859
rect 25329 37281 25363 37315
rect 25145 37145 25179 37179
rect 25329 36873 25363 36907
rect 24409 36737 24443 36771
rect 24685 36737 24719 36771
rect 24225 36125 24259 36159
rect 24685 36125 24719 36159
rect 25329 35989 25363 36023
rect 21189 35785 21223 35819
rect 22477 35785 22511 35819
rect 11529 35717 11563 35751
rect 20453 35717 20487 35751
rect 21097 35717 21131 35751
rect 9413 35649 9447 35683
rect 22385 35649 22419 35683
rect 24685 35649 24719 35683
rect 25329 35649 25363 35683
rect 9689 35581 9723 35615
rect 21281 35581 21315 35615
rect 22569 35581 22603 35615
rect 22017 35513 22051 35547
rect 11161 35445 11195 35479
rect 11805 35445 11839 35479
rect 20729 35445 20763 35479
rect 24501 35445 24535 35479
rect 25145 35445 25179 35479
rect 25329 35241 25363 35275
rect 23305 35105 23339 35139
rect 24225 35037 24259 35071
rect 24685 35037 24719 35071
rect 23121 34969 23155 35003
rect 23213 34969 23247 35003
rect 21925 34901 21959 34935
rect 22385 34901 22419 34935
rect 22753 34901 22787 34935
rect 21465 34697 21499 34731
rect 25145 34697 25179 34731
rect 24869 34561 24903 34595
rect 25329 34561 25363 34595
rect 9137 34153 9171 34187
rect 21912 34153 21946 34187
rect 15393 34017 15427 34051
rect 21649 34017 21683 34051
rect 9321 33949 9355 33983
rect 19441 33949 19475 33983
rect 24869 33949 24903 33983
rect 25329 33949 25363 33983
rect 14657 33881 14691 33915
rect 15853 33881 15887 33915
rect 19717 33881 19751 33915
rect 19073 33813 19107 33847
rect 21189 33813 21223 33847
rect 23397 33813 23431 33847
rect 25145 33813 25179 33847
rect 25145 33609 25179 33643
rect 19809 33541 19843 33575
rect 21557 33541 21591 33575
rect 19533 33473 19567 33507
rect 22017 33473 22051 33507
rect 25329 33473 25363 33507
rect 22293 33405 22327 33439
rect 23765 33405 23799 33439
rect 19257 33269 19291 33303
rect 21281 33269 21315 33303
rect 24409 33269 24443 33303
rect 24869 33269 24903 33303
rect 16681 33065 16715 33099
rect 21925 33065 21959 33099
rect 24041 33065 24075 33099
rect 19625 32997 19659 33031
rect 16037 32929 16071 32963
rect 16129 32929 16163 32963
rect 17049 32929 17083 32963
rect 22293 32929 22327 32963
rect 22569 32929 22603 32963
rect 25237 32929 25271 32963
rect 16773 32861 16807 32895
rect 20637 32861 20671 32895
rect 25053 32861 25087 32895
rect 15945 32793 15979 32827
rect 19901 32793 19935 32827
rect 24961 32793 24995 32827
rect 15577 32725 15611 32759
rect 24593 32725 24627 32759
rect 17049 32521 17083 32555
rect 18797 32521 18831 32555
rect 25237 32521 25271 32555
rect 15393 32453 15427 32487
rect 22845 32453 22879 32487
rect 22109 32385 22143 32419
rect 23489 32385 23523 32419
rect 16129 32317 16163 32351
rect 16865 32317 16899 32351
rect 19073 32317 19107 32351
rect 19349 32317 19383 32351
rect 23765 32317 23799 32351
rect 20821 32181 20855 32215
rect 21649 32181 21683 32215
rect 17036 31977 17070 32011
rect 18889 31977 18923 32011
rect 19073 31977 19107 32011
rect 24041 31977 24075 32011
rect 15577 31909 15611 31943
rect 21649 31909 21683 31943
rect 23029 31909 23063 31943
rect 25145 31909 25179 31943
rect 16129 31841 16163 31875
rect 18521 31841 18555 31875
rect 19717 31841 19751 31875
rect 22201 31841 22235 31875
rect 23489 31841 23523 31875
rect 23581 31841 23615 31875
rect 16037 31773 16071 31807
rect 16773 31773 16807 31807
rect 19441 31773 19475 31807
rect 22109 31773 22143 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 15945 31637 15979 31671
rect 21189 31637 21223 31671
rect 22017 31637 22051 31671
rect 22661 31637 22695 31671
rect 23397 31637 23431 31671
rect 16681 31433 16715 31467
rect 19165 31433 19199 31467
rect 20545 31433 20579 31467
rect 19441 31365 19475 31399
rect 22753 31365 22787 31399
rect 17417 31297 17451 31331
rect 19809 31297 19843 31331
rect 20453 31297 20487 31331
rect 22477 31297 22511 31331
rect 25329 31297 25363 31331
rect 13369 31229 13403 31263
rect 13645 31229 13679 31263
rect 15485 31229 15519 31263
rect 16405 31229 16439 31263
rect 17693 31229 17727 31263
rect 20637 31229 20671 31263
rect 22201 31229 22235 31263
rect 21557 31161 21591 31195
rect 15117 31093 15151 31127
rect 15761 31093 15795 31127
rect 20085 31093 20119 31127
rect 24225 31093 24259 31127
rect 25145 31093 25179 31127
rect 9137 30889 9171 30923
rect 15577 30889 15611 30923
rect 15761 30889 15795 30923
rect 18521 30889 18555 30923
rect 18889 30889 18923 30923
rect 19717 30889 19751 30923
rect 22477 30889 22511 30923
rect 25513 30889 25547 30923
rect 16773 30753 16807 30787
rect 20729 30753 20763 30787
rect 9321 30685 9355 30719
rect 14381 30685 14415 30719
rect 15117 30617 15151 30651
rect 17049 30617 17083 30651
rect 21005 30617 21039 30651
rect 24593 30617 24627 30651
rect 20085 30549 20119 30583
rect 23213 30549 23247 30583
rect 18981 30345 19015 30379
rect 20269 30345 20303 30379
rect 14105 30277 14139 30311
rect 20361 30277 20395 30311
rect 22477 30277 22511 30311
rect 23581 30277 23615 30311
rect 9137 30209 9171 30243
rect 11805 30209 11839 30243
rect 15853 30209 15887 30243
rect 21281 30209 21315 30243
rect 22385 30209 22419 30243
rect 12081 30141 12115 30175
rect 14841 30141 14875 30175
rect 15945 30141 15979 30175
rect 16037 30141 16071 30175
rect 20545 30141 20579 30175
rect 22661 30141 22695 30175
rect 23305 30141 23339 30175
rect 25053 30141 25087 30175
rect 8953 30073 8987 30107
rect 13553 30005 13587 30039
rect 15485 30005 15519 30039
rect 16681 30005 16715 30039
rect 16865 30005 16899 30039
rect 19901 30005 19935 30039
rect 22017 30005 22051 30039
rect 13461 29801 13495 29835
rect 16313 29801 16347 29835
rect 18797 29801 18831 29835
rect 25145 29801 25179 29835
rect 12909 29733 12943 29767
rect 16497 29733 16531 29767
rect 23857 29733 23891 29767
rect 11161 29665 11195 29699
rect 15853 29665 15887 29699
rect 17049 29665 17083 29699
rect 20729 29665 20763 29699
rect 15577 29597 15611 29631
rect 20637 29597 20671 29631
rect 23397 29597 23431 29631
rect 24041 29597 24075 29631
rect 25329 29597 25363 29631
rect 11437 29529 11471 29563
rect 15669 29529 15703 29563
rect 17325 29529 17359 29563
rect 22937 29529 22971 29563
rect 13277 29461 13311 29495
rect 13737 29461 13771 29495
rect 15209 29461 15243 29495
rect 19441 29461 19475 29495
rect 20177 29461 20211 29495
rect 20545 29461 20579 29495
rect 23213 29461 23247 29495
rect 24501 29461 24535 29495
rect 9505 29257 9539 29291
rect 12541 29257 12575 29291
rect 12633 29257 12667 29291
rect 15117 29257 15151 29291
rect 16037 29257 16071 29291
rect 18797 29257 18831 29291
rect 19165 29257 19199 29291
rect 23949 29257 23983 29291
rect 25421 29257 25455 29291
rect 9873 29189 9907 29223
rect 15945 29189 15979 29223
rect 19257 29189 19291 29223
rect 9965 29121 9999 29155
rect 13369 29121 13403 29155
rect 17233 29121 17267 29155
rect 17325 29121 17359 29155
rect 17877 29121 17911 29155
rect 20453 29121 20487 29155
rect 22201 29121 22235 29155
rect 24041 29121 24075 29155
rect 25329 29121 25363 29155
rect 10057 29053 10091 29087
rect 12817 29053 12851 29087
rect 16129 29053 16163 29087
rect 17417 29053 17451 29087
rect 19441 29053 19475 29087
rect 23029 29053 23063 29087
rect 24133 29053 24167 29087
rect 24777 29053 24811 29087
rect 12173 28985 12207 29019
rect 15577 28985 15611 29019
rect 16865 28985 16899 29019
rect 18061 28985 18095 29019
rect 19993 28985 20027 29019
rect 21833 28985 21867 29019
rect 23581 28985 23615 29019
rect 13632 28917 13666 28951
rect 10885 28713 10919 28747
rect 16313 28713 16347 28747
rect 18889 28713 18923 28747
rect 22385 28713 22419 28747
rect 15945 28645 15979 28679
rect 22845 28645 22879 28679
rect 24041 28645 24075 28679
rect 9137 28577 9171 28611
rect 11437 28577 11471 28611
rect 13185 28577 13219 28611
rect 15301 28577 15335 28611
rect 15393 28577 15427 28611
rect 17417 28577 17451 28611
rect 20085 28577 20119 28611
rect 23397 28577 23431 28611
rect 25053 28577 25087 28611
rect 25237 28577 25271 28611
rect 17141 28509 17175 28543
rect 20637 28509 20671 28543
rect 23305 28509 23339 28543
rect 24961 28509 24995 28543
rect 9413 28441 9447 28475
rect 11713 28441 11747 28475
rect 15209 28441 15243 28475
rect 19901 28441 19935 28475
rect 20913 28441 20947 28475
rect 13553 28373 13587 28407
rect 14841 28373 14875 28407
rect 16037 28373 16071 28407
rect 19441 28373 19475 28407
rect 19809 28373 19843 28407
rect 23213 28373 23247 28407
rect 23949 28373 23983 28407
rect 24593 28373 24627 28407
rect 13829 28169 13863 28203
rect 15577 28169 15611 28203
rect 16405 28169 16439 28203
rect 17233 28169 17267 28203
rect 18981 28169 19015 28203
rect 19717 28169 19751 28203
rect 22477 28169 22511 28203
rect 11989 28101 12023 28135
rect 18705 28101 18739 28135
rect 21097 28101 21131 28135
rect 23489 28101 23523 28135
rect 15669 28033 15703 28067
rect 20361 28033 20395 28067
rect 22385 28033 22419 28067
rect 23213 28033 23247 28067
rect 11713 27965 11747 27999
rect 15761 27965 15795 27999
rect 17325 27965 17359 27999
rect 17417 27965 17451 27999
rect 18061 27965 18095 27999
rect 22569 27965 22603 27999
rect 19349 27897 19383 27931
rect 22017 27897 22051 27931
rect 10977 27829 11011 27863
rect 13461 27829 13495 27863
rect 15209 27829 15243 27863
rect 16313 27829 16347 27863
rect 16865 27829 16899 27863
rect 18521 27829 18555 27863
rect 21557 27829 21591 27863
rect 24961 27829 24995 27863
rect 25237 27829 25271 27863
rect 25513 27829 25547 27863
rect 12633 27625 12667 27659
rect 16497 27625 16531 27659
rect 20164 27625 20198 27659
rect 23857 27625 23891 27659
rect 9137 27557 9171 27591
rect 7665 27489 7699 27523
rect 10517 27489 10551 27523
rect 10793 27489 10827 27523
rect 13553 27489 13587 27523
rect 15761 27489 15795 27523
rect 18061 27489 18095 27523
rect 19901 27489 19935 27523
rect 22109 27489 22143 27523
rect 24133 27489 24167 27523
rect 25053 27489 25087 27523
rect 25145 27489 25179 27523
rect 7389 27421 7423 27455
rect 13461 27421 13495 27455
rect 15669 27421 15703 27455
rect 17877 27421 17911 27455
rect 9045 27353 9079 27387
rect 13369 27353 13403 27387
rect 16221 27353 16255 27387
rect 17969 27353 18003 27387
rect 22385 27353 22419 27387
rect 12265 27285 12299 27319
rect 13001 27285 13035 27319
rect 15209 27285 15243 27319
rect 15577 27285 15611 27319
rect 17509 27285 17543 27319
rect 19625 27285 19659 27319
rect 21649 27285 21683 27319
rect 24593 27285 24627 27319
rect 24961 27285 24995 27319
rect 15669 27081 15703 27115
rect 22845 27081 22879 27115
rect 25329 27081 25363 27115
rect 11621 27013 11655 27047
rect 13369 27013 13403 27047
rect 15761 27013 15795 27047
rect 7665 26945 7699 26979
rect 9321 26945 9355 26979
rect 13093 26945 13127 26979
rect 17969 26945 18003 26979
rect 22753 26945 22787 26979
rect 7941 26877 7975 26911
rect 9597 26877 9631 26911
rect 11069 26877 11103 26911
rect 15853 26877 15887 26911
rect 18245 26877 18279 26911
rect 23029 26877 23063 26911
rect 23581 26877 23615 26911
rect 23857 26877 23891 26911
rect 14841 26741 14875 26775
rect 15301 26741 15335 26775
rect 19717 26741 19751 26775
rect 20085 26741 20119 26775
rect 21557 26741 21591 26775
rect 21925 26741 21959 26775
rect 22385 26741 22419 26775
rect 11345 26537 11379 26571
rect 21189 26537 21223 26571
rect 11253 26469 11287 26503
rect 15669 26469 15703 26503
rect 18981 26469 19015 26503
rect 22661 26469 22695 26503
rect 23857 26469 23891 26503
rect 24593 26469 24627 26503
rect 9137 26401 9171 26435
rect 10885 26401 10919 26435
rect 14841 26401 14875 26435
rect 15393 26401 15427 26435
rect 16221 26401 16255 26435
rect 19441 26401 19475 26435
rect 19717 26401 19751 26435
rect 23213 26401 23247 26435
rect 25145 26401 25179 26435
rect 16681 26333 16715 26367
rect 16865 26333 16899 26367
rect 22109 26333 22143 26367
rect 24041 26333 24075 26367
rect 9413 26265 9447 26299
rect 14657 26265 14691 26299
rect 16129 26265 16163 26299
rect 17049 26265 17083 26299
rect 22385 26265 22419 26299
rect 23121 26265 23155 26299
rect 24961 26265 24995 26299
rect 25053 26265 25087 26299
rect 14289 26197 14323 26231
rect 14749 26197 14783 26231
rect 16037 26197 16071 26231
rect 17233 26197 17267 26231
rect 18245 26197 18279 26231
rect 23029 26197 23063 26231
rect 9505 25993 9539 26027
rect 12173 25993 12207 26027
rect 12633 25993 12667 26027
rect 16865 25993 16899 26027
rect 17785 25993 17819 26027
rect 18153 25993 18187 26027
rect 19073 25993 19107 26027
rect 22477 25993 22511 26027
rect 13921 25925 13955 25959
rect 14013 25925 14047 25959
rect 18245 25925 18279 25959
rect 8033 25857 8067 25891
rect 12541 25857 12575 25891
rect 15209 25857 15243 25891
rect 16037 25857 16071 25891
rect 17049 25857 17083 25891
rect 22385 25857 22419 25891
rect 23489 25857 23523 25891
rect 23949 25857 23983 25891
rect 8309 25789 8343 25823
rect 12725 25789 12759 25823
rect 14105 25789 14139 25823
rect 15301 25789 15335 25823
rect 15393 25789 15427 25823
rect 18429 25789 18463 25823
rect 22661 25789 22695 25823
rect 25145 25789 25179 25823
rect 13553 25653 13587 25687
rect 14841 25653 14875 25687
rect 17417 25653 17451 25687
rect 21557 25653 21591 25687
rect 22017 25653 22051 25687
rect 23305 25653 23339 25687
rect 14289 25449 14323 25483
rect 17601 25449 17635 25483
rect 18337 25449 18371 25483
rect 20361 25449 20395 25483
rect 21557 25449 21591 25483
rect 25329 25449 25363 25483
rect 15301 25381 15335 25415
rect 16957 25381 16991 25415
rect 10885 25313 10919 25347
rect 11161 25313 11195 25347
rect 14841 25313 14875 25347
rect 16313 25313 16347 25347
rect 12909 25245 12943 25279
rect 17141 25245 17175 25279
rect 17785 25245 17819 25279
rect 18153 25245 18187 25279
rect 19809 25245 19843 25279
rect 20453 25245 20487 25279
rect 21005 25245 21039 25279
rect 21741 25245 21775 25279
rect 22661 25245 22695 25279
rect 24685 25245 24719 25279
rect 14657 25177 14691 25211
rect 16221 25177 16255 25211
rect 19349 25177 19383 25211
rect 23857 25177 23891 25211
rect 12633 25109 12667 25143
rect 14749 25109 14783 25143
rect 15761 25109 15795 25143
rect 16129 25109 16163 25143
rect 18705 25109 18739 25143
rect 19901 25109 19935 25143
rect 20821 25109 20855 25143
rect 15117 24905 15151 24939
rect 15485 24905 15519 24939
rect 17233 24905 17267 24939
rect 12081 24837 12115 24871
rect 22477 24837 22511 24871
rect 12173 24769 12207 24803
rect 13001 24769 13035 24803
rect 17325 24769 17359 24803
rect 18429 24769 18463 24803
rect 18521 24769 18555 24803
rect 19073 24769 19107 24803
rect 19717 24769 19751 24803
rect 22569 24769 22603 24803
rect 9413 24701 9447 24735
rect 9689 24701 9723 24735
rect 12265 24701 12299 24735
rect 13277 24701 13311 24735
rect 14749 24701 14783 24735
rect 15393 24701 15427 24735
rect 17417 24701 17451 24735
rect 18613 24701 18647 24735
rect 19993 24701 20027 24735
rect 21465 24701 21499 24735
rect 22753 24701 22787 24735
rect 23581 24701 23615 24735
rect 23857 24701 23891 24735
rect 25329 24701 25363 24735
rect 19257 24633 19291 24667
rect 11161 24565 11195 24599
rect 11713 24565 11747 24599
rect 16865 24565 16899 24599
rect 18061 24565 18095 24599
rect 22109 24565 22143 24599
rect 23305 24565 23339 24599
rect 21189 24361 21223 24395
rect 22188 24361 22222 24395
rect 11345 24293 11379 24327
rect 11437 24293 11471 24327
rect 25145 24293 25179 24327
rect 9413 24225 9447 24259
rect 11989 24225 12023 24259
rect 18797 24225 18831 24259
rect 19441 24225 19475 24259
rect 21925 24225 21959 24259
rect 9137 24157 9171 24191
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 24869 24157 24903 24191
rect 25329 24157 25363 24191
rect 12265 24089 12299 24123
rect 15945 24089 15979 24123
rect 19717 24089 19751 24123
rect 10885 24021 10919 24055
rect 13737 24021 13771 24055
rect 14105 24021 14139 24055
rect 18153 24021 18187 24055
rect 18613 24021 18647 24055
rect 21557 24021 21591 24055
rect 23673 24021 23707 24055
rect 9781 23817 9815 23851
rect 10425 23817 10459 23851
rect 10793 23817 10827 23851
rect 14473 23817 14507 23851
rect 14933 23817 14967 23851
rect 17325 23817 17359 23851
rect 18705 23817 18739 23851
rect 18889 23817 18923 23851
rect 20913 23817 20947 23851
rect 22201 23817 22235 23851
rect 24961 23817 24995 23851
rect 25421 23817 25455 23851
rect 11621 23749 11655 23783
rect 13645 23749 13679 23783
rect 8033 23681 8067 23715
rect 13737 23681 13771 23715
rect 14841 23681 14875 23715
rect 17233 23681 17267 23715
rect 18245 23681 18279 23715
rect 18613 23681 18647 23715
rect 19625 23681 19659 23715
rect 20821 23681 20855 23715
rect 22385 23681 22419 23715
rect 8309 23613 8343 23647
rect 10885 23613 10919 23647
rect 10977 23613 11011 23647
rect 13829 23613 13863 23647
rect 15025 23613 15059 23647
rect 15669 23613 15703 23647
rect 17417 23613 17451 23647
rect 19717 23613 19751 23647
rect 19901 23613 19935 23647
rect 21005 23613 21039 23647
rect 23213 23613 23247 23647
rect 23489 23613 23523 23647
rect 18061 23545 18095 23579
rect 10057 23477 10091 23511
rect 13277 23477 13311 23511
rect 16865 23477 16899 23511
rect 19257 23477 19291 23511
rect 20453 23477 20487 23511
rect 21925 23477 21959 23511
rect 22845 23477 22879 23511
rect 25329 23477 25363 23511
rect 10793 23273 10827 23307
rect 15853 23273 15887 23307
rect 14749 23205 14783 23239
rect 17877 23205 17911 23239
rect 19533 23205 19567 23239
rect 9689 23137 9723 23171
rect 11713 23137 11747 23171
rect 11805 23137 11839 23171
rect 13553 23137 13587 23171
rect 15301 23137 15335 23171
rect 18521 23137 18555 23171
rect 18981 23137 19015 23171
rect 20177 23137 20211 23171
rect 20729 23137 20763 23171
rect 25237 23137 25271 23171
rect 9321 23069 9355 23103
rect 11621 23069 11655 23103
rect 14381 23069 14415 23103
rect 15117 23069 15151 23103
rect 18245 23069 18279 23103
rect 19901 23069 19935 23103
rect 19993 23069 20027 23103
rect 21833 23069 21867 23103
rect 22845 23069 22879 23103
rect 25053 23069 25087 23103
rect 13369 23001 13403 23035
rect 15209 23001 15243 23035
rect 23857 23001 23891 23035
rect 24961 23001 24995 23035
rect 11253 22933 11287 22967
rect 13001 22933 13035 22967
rect 13461 22933 13495 22967
rect 14197 22933 14231 22967
rect 18337 22933 18371 22967
rect 21649 22933 21683 22967
rect 24593 22933 24627 22967
rect 10149 22729 10183 22763
rect 14473 22729 14507 22763
rect 16865 22729 16899 22763
rect 18797 22729 18831 22763
rect 18889 22729 18923 22763
rect 19717 22729 19751 22763
rect 21189 22729 21223 22763
rect 25145 22661 25179 22695
rect 8125 22593 8159 22627
rect 12357 22593 12391 22627
rect 17049 22593 17083 22627
rect 21097 22593 21131 22627
rect 22109 22593 22143 22627
rect 23949 22593 23983 22627
rect 8401 22525 8435 22559
rect 12633 22525 12667 22559
rect 21281 22525 21315 22559
rect 23305 22525 23339 22559
rect 20361 22457 20395 22491
rect 9873 22389 9907 22423
rect 14105 22389 14139 22423
rect 14657 22389 14691 22423
rect 20729 22389 20763 22423
rect 21820 22185 21854 22219
rect 23305 22185 23339 22219
rect 9689 22049 9723 22083
rect 11345 22049 11379 22083
rect 12449 22049 12483 22083
rect 12541 22049 12575 22083
rect 15301 22049 15335 22083
rect 15393 22049 15427 22083
rect 16129 22049 16163 22083
rect 20361 22049 20395 22083
rect 21557 22049 21591 22083
rect 25053 22049 25087 22083
rect 25237 22049 25271 22083
rect 11161 21981 11195 22015
rect 18153 21981 18187 22015
rect 23857 21981 23891 22015
rect 9597 21913 9631 21947
rect 16405 21913 16439 21947
rect 24961 21913 24995 21947
rect 9137 21845 9171 21879
rect 9505 21845 9539 21879
rect 10425 21845 10459 21879
rect 10701 21845 10735 21879
rect 11069 21845 11103 21879
rect 11989 21845 12023 21879
rect 12357 21845 12391 21879
rect 14841 21845 14875 21879
rect 15209 21845 15243 21879
rect 17877 21845 17911 21879
rect 19717 21845 19751 21879
rect 20085 21845 20119 21879
rect 20177 21845 20211 21879
rect 20913 21845 20947 21879
rect 24593 21845 24627 21879
rect 10425 21641 10459 21675
rect 10793 21641 10827 21675
rect 11713 21641 11747 21675
rect 15209 21641 15243 21675
rect 19165 21641 19199 21675
rect 19993 21641 20027 21675
rect 21189 21641 21223 21675
rect 22477 21641 22511 21675
rect 25053 21641 25087 21675
rect 10885 21573 10919 21607
rect 21373 21573 21407 21607
rect 9597 21505 9631 21539
rect 13093 21505 13127 21539
rect 15669 21505 15703 21539
rect 18889 21505 18923 21539
rect 19901 21505 19935 21539
rect 20729 21505 20763 21539
rect 22385 21505 22419 21539
rect 23305 21505 23339 21539
rect 6929 21437 6963 21471
rect 7205 21437 7239 21471
rect 9689 21437 9723 21471
rect 9781 21437 9815 21471
rect 11069 21437 11103 21471
rect 13369 21437 13403 21471
rect 14841 21437 14875 21471
rect 20085 21437 20119 21471
rect 22661 21437 22695 21471
rect 23581 21437 23615 21471
rect 21649 21369 21683 21403
rect 8677 21301 8711 21335
rect 9229 21301 9263 21335
rect 15761 21301 15795 21335
rect 18705 21301 18739 21335
rect 19533 21301 19567 21335
rect 22017 21301 22051 21335
rect 25329 21301 25363 21335
rect 12449 21097 12483 21131
rect 16957 21097 16991 21131
rect 19441 21029 19475 21063
rect 20821 21029 20855 21063
rect 24593 21029 24627 21063
rect 9965 20961 9999 20995
rect 15209 20961 15243 20995
rect 19993 20961 20027 20995
rect 22017 20961 22051 20995
rect 23857 20961 23891 20995
rect 25145 20961 25179 20995
rect 10701 20893 10735 20927
rect 19809 20893 19843 20927
rect 20453 20893 20487 20927
rect 21005 20893 21039 20927
rect 22661 20893 22695 20927
rect 25053 20893 25087 20927
rect 9229 20825 9263 20859
rect 10977 20825 11011 20859
rect 15485 20825 15519 20859
rect 19901 20825 19935 20859
rect 21281 20825 21315 20859
rect 24961 20825 24995 20859
rect 9045 20757 9079 20791
rect 12817 20757 12851 20791
rect 14657 20757 14691 20791
rect 17325 20757 17359 20791
rect 18797 20757 18831 20791
rect 21465 20757 21499 20791
rect 10425 20553 10459 20587
rect 10793 20553 10827 20587
rect 15485 20553 15519 20587
rect 20913 20553 20947 20587
rect 22937 20553 22971 20587
rect 25329 20553 25363 20587
rect 8033 20485 8067 20519
rect 17141 20485 17175 20519
rect 12725 20417 12759 20451
rect 15393 20417 15427 20451
rect 16865 20417 16899 20451
rect 19257 20417 19291 20451
rect 19901 20417 19935 20451
rect 20821 20417 20855 20451
rect 21465 20417 21499 20451
rect 22201 20417 22235 20451
rect 23121 20417 23155 20451
rect 7757 20349 7791 20383
rect 9781 20349 9815 20383
rect 10885 20349 10919 20383
rect 10977 20349 11011 20383
rect 13001 20349 13035 20383
rect 15577 20349 15611 20383
rect 18613 20349 18647 20383
rect 21097 20349 21131 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 20453 20281 20487 20315
rect 22017 20281 22051 20315
rect 10149 20213 10183 20247
rect 14473 20213 14507 20247
rect 15025 20213 15059 20247
rect 19073 20213 19107 20247
rect 19717 20213 19751 20247
rect 22477 20213 22511 20247
rect 8493 20009 8527 20043
rect 11345 20009 11379 20043
rect 14552 20009 14586 20043
rect 16037 20009 16071 20043
rect 16957 20009 16991 20043
rect 23857 20009 23891 20043
rect 25329 20009 25363 20043
rect 21649 19941 21683 19975
rect 11989 19873 12023 19907
rect 14289 19873 14323 19907
rect 17969 19873 18003 19907
rect 18061 19873 18095 19907
rect 19901 19873 19935 19907
rect 22109 19873 22143 19907
rect 22385 19873 22419 19907
rect 9137 19805 9171 19839
rect 16681 19805 16715 19839
rect 18889 19805 18923 19839
rect 24777 19805 24811 19839
rect 9413 19737 9447 19771
rect 11805 19737 11839 19771
rect 17877 19737 17911 19771
rect 20177 19737 20211 19771
rect 10885 19669 10919 19703
rect 11713 19669 11747 19703
rect 16497 19669 16531 19703
rect 17509 19669 17543 19703
rect 18705 19669 18739 19703
rect 19533 19669 19567 19703
rect 24133 19669 24167 19703
rect 24593 19669 24627 19703
rect 8769 19465 8803 19499
rect 10977 19465 11011 19499
rect 11713 19465 11747 19499
rect 15025 19465 15059 19499
rect 16865 19465 16899 19499
rect 17233 19465 17267 19499
rect 17325 19465 17359 19499
rect 18981 19465 19015 19499
rect 20453 19465 20487 19499
rect 20545 19465 20579 19499
rect 22661 19465 22695 19499
rect 25145 19465 25179 19499
rect 9137 19397 9171 19431
rect 23673 19397 23707 19431
rect 12541 19329 12575 19363
rect 15209 19329 15243 19363
rect 16129 19329 16163 19363
rect 19165 19329 19199 19363
rect 21281 19329 21315 19363
rect 22569 19329 22603 19363
rect 23397 19329 23431 19363
rect 6561 19261 6595 19295
rect 6837 19261 6871 19295
rect 9229 19261 9263 19295
rect 9321 19261 9355 19295
rect 12817 19261 12851 19295
rect 17417 19261 17451 19295
rect 17877 19261 17911 19295
rect 20637 19261 20671 19295
rect 22753 19261 22787 19295
rect 18061 19193 18095 19227
rect 22201 19193 22235 19227
rect 8309 19125 8343 19159
rect 11161 19125 11195 19159
rect 14289 19125 14323 19159
rect 14565 19125 14599 19159
rect 15945 19125 15979 19159
rect 20085 19125 20119 19159
rect 21833 19125 21867 19159
rect 8677 18921 8711 18955
rect 10057 18921 10091 18955
rect 11161 18921 11195 18955
rect 11529 18921 11563 18955
rect 12725 18921 12759 18955
rect 18153 18853 18187 18887
rect 6929 18785 6963 18819
rect 10609 18785 10643 18819
rect 12081 18785 12115 18819
rect 13277 18785 13311 18819
rect 17325 18785 17359 18819
rect 17509 18785 17543 18819
rect 18705 18785 18739 18819
rect 23489 18785 23523 18819
rect 6653 18717 6687 18751
rect 10517 18717 10551 18751
rect 17233 18717 17267 18751
rect 21465 18717 21499 18751
rect 22201 18717 22235 18751
rect 22845 18717 22879 18751
rect 25145 18717 25179 18751
rect 11989 18649 12023 18683
rect 13093 18649 13127 18683
rect 18521 18649 18555 18683
rect 24685 18649 24719 18683
rect 24869 18649 24903 18683
rect 8401 18581 8435 18615
rect 9689 18581 9723 18615
rect 10425 18581 10459 18615
rect 11897 18581 11931 18615
rect 13185 18581 13219 18615
rect 13829 18581 13863 18615
rect 14289 18581 14323 18615
rect 16865 18581 16899 18615
rect 18613 18581 18647 18615
rect 21281 18581 21315 18615
rect 22017 18581 22051 18615
rect 9505 18377 9539 18411
rect 10425 18377 10459 18411
rect 11069 18377 11103 18411
rect 11253 18377 11287 18411
rect 13829 18377 13863 18411
rect 14197 18377 14231 18411
rect 14933 18377 14967 18411
rect 8033 18309 8067 18343
rect 13185 18309 13219 18343
rect 23305 18309 23339 18343
rect 10333 18241 10367 18275
rect 12449 18241 12483 18275
rect 16865 18241 16899 18275
rect 19993 18241 20027 18275
rect 21281 18241 21315 18275
rect 22109 18241 22143 18275
rect 23949 18241 23983 18275
rect 7757 18173 7791 18207
rect 10517 18173 10551 18207
rect 14289 18173 14323 18207
rect 14381 18173 14415 18207
rect 17141 18173 17175 18207
rect 24685 18173 24719 18207
rect 9965 18105 9999 18139
rect 19809 18105 19843 18139
rect 18613 18037 18647 18071
rect 18889 18037 18923 18071
rect 21097 18037 21131 18071
rect 7849 17833 7883 17867
rect 18429 17833 18463 17867
rect 18981 17833 19015 17867
rect 21649 17833 21683 17867
rect 12265 17765 12299 17799
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 12909 17697 12943 17731
rect 16405 17697 16439 17731
rect 17969 17697 18003 17731
rect 19625 17697 19659 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 9781 17629 9815 17663
rect 11805 17629 11839 17663
rect 12633 17629 12667 17663
rect 16129 17629 16163 17663
rect 17785 17629 17819 17663
rect 18797 17629 18831 17663
rect 19901 17629 19935 17663
rect 21097 17629 21131 17663
rect 22017 17629 22051 17663
rect 22845 17629 22879 17663
rect 8217 17561 8251 17595
rect 14197 17561 14231 17595
rect 17877 17561 17911 17595
rect 18613 17561 18647 17595
rect 22201 17561 22235 17595
rect 7205 17493 7239 17527
rect 8309 17493 8343 17527
rect 9137 17493 9171 17527
rect 12725 17493 12759 17527
rect 13461 17493 13495 17527
rect 15485 17493 15519 17527
rect 17417 17493 17451 17527
rect 20913 17493 20947 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 8033 17289 8067 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 11621 17289 11655 17323
rect 13185 17289 13219 17323
rect 20361 17289 20395 17323
rect 22753 17289 22787 17323
rect 10977 17221 11011 17255
rect 16957 17221 16991 17255
rect 17969 17221 18003 17255
rect 23765 17221 23799 17255
rect 10241 17153 10275 17187
rect 14565 17153 14599 17187
rect 21281 17153 21315 17187
rect 22661 17153 22695 17187
rect 23489 17153 23523 17187
rect 8125 17085 8159 17119
rect 8309 17085 8343 17119
rect 8769 17085 8803 17119
rect 9505 17085 9539 17119
rect 9597 17085 9631 17119
rect 11897 17085 11931 17119
rect 12541 17085 12575 17119
rect 13277 17085 13311 17119
rect 13461 17085 13495 17119
rect 14841 17085 14875 17119
rect 16313 17085 16347 17119
rect 18613 17085 18647 17119
rect 18889 17085 18923 17119
rect 22937 17085 22971 17119
rect 25237 17085 25271 17119
rect 7665 17017 7699 17051
rect 17141 17017 17175 17051
rect 18153 17017 18187 17051
rect 7297 16949 7331 16983
rect 12081 16949 12115 16983
rect 12817 16949 12851 16983
rect 17509 16949 17543 16983
rect 21925 16949 21959 16983
rect 22293 16949 22327 16983
rect 8585 16745 8619 16779
rect 11253 16745 11287 16779
rect 13921 16745 13955 16779
rect 15761 16745 15795 16779
rect 16865 16745 16899 16779
rect 19993 16745 20027 16779
rect 22293 16745 22327 16779
rect 24593 16745 24627 16779
rect 10701 16609 10735 16643
rect 10885 16609 10919 16643
rect 11805 16609 11839 16643
rect 15117 16609 15151 16643
rect 16313 16609 16347 16643
rect 17969 16609 18003 16643
rect 14933 16541 14967 16575
rect 18889 16541 18923 16575
rect 20269 16541 20303 16575
rect 22661 16541 22695 16575
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 10609 16473 10643 16507
rect 12081 16473 12115 16507
rect 17233 16473 17267 16507
rect 20545 16473 20579 16507
rect 9965 16405 9999 16439
rect 10241 16405 10275 16439
rect 13553 16405 13587 16439
rect 14289 16405 14323 16439
rect 14565 16405 14599 16439
rect 15025 16405 15059 16439
rect 16129 16405 16163 16439
rect 16221 16405 16255 16439
rect 18705 16405 18739 16439
rect 19257 16405 19291 16439
rect 22017 16405 22051 16439
rect 8309 16201 8343 16235
rect 8677 16201 8711 16235
rect 13369 16201 13403 16235
rect 13829 16201 13863 16235
rect 14565 16201 14599 16235
rect 15761 16201 15795 16235
rect 16865 16201 16899 16235
rect 21189 16201 21223 16235
rect 11805 16133 11839 16167
rect 12541 16133 12575 16167
rect 20085 16133 20119 16167
rect 6561 16065 6595 16099
rect 12633 16065 12667 16099
rect 13737 16065 13771 16099
rect 14933 16065 14967 16099
rect 17233 16065 17267 16099
rect 18061 16065 18095 16099
rect 18705 16065 18739 16099
rect 19257 16065 19291 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 6837 15997 6871 16031
rect 12725 15997 12759 16031
rect 14013 15997 14047 16031
rect 15025 15997 15059 16031
rect 15117 15997 15151 16031
rect 21373 15997 21407 16031
rect 22293 15997 22327 16031
rect 24501 15997 24535 16031
rect 24777 15997 24811 16031
rect 12173 15929 12207 15963
rect 16221 15861 16255 15895
rect 17325 15861 17359 15895
rect 17877 15861 17911 15895
rect 18521 15861 18555 15895
rect 20729 15861 20763 15895
rect 23765 15861 23799 15895
rect 9137 15657 9171 15691
rect 10149 15657 10183 15691
rect 11621 15657 11655 15691
rect 15485 15657 15519 15691
rect 9689 15521 9723 15555
rect 12265 15521 12299 15555
rect 12633 15521 12667 15555
rect 16405 15521 16439 15555
rect 16681 15521 16715 15555
rect 19441 15521 19475 15555
rect 22293 15521 22327 15555
rect 22569 15521 22603 15555
rect 24593 15521 24627 15555
rect 13185 15453 13219 15487
rect 21833 15453 21867 15487
rect 9597 15385 9631 15419
rect 11989 15385 12023 15419
rect 19717 15385 19751 15419
rect 9505 15317 9539 15351
rect 12081 15317 12115 15351
rect 14289 15317 14323 15351
rect 14749 15317 14783 15351
rect 15761 15317 15795 15351
rect 18153 15317 18187 15351
rect 18429 15317 18463 15351
rect 18981 15317 19015 15351
rect 21189 15317 21223 15351
rect 21649 15317 21683 15351
rect 24041 15317 24075 15351
rect 10149 15113 10183 15147
rect 11345 15113 11379 15147
rect 14105 15113 14139 15147
rect 15945 15113 15979 15147
rect 17509 15113 17543 15147
rect 20085 15113 20119 15147
rect 18705 15045 18739 15079
rect 23305 15045 23339 15079
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 16037 14977 16071 15011
rect 19993 14977 20027 15011
rect 21005 14977 21039 15011
rect 21557 14977 21591 15011
rect 22109 14977 22143 15011
rect 24133 14977 24167 15011
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 9689 14909 9723 14943
rect 10701 14909 10735 14943
rect 14197 14909 14231 14943
rect 14381 14909 14415 14943
rect 16221 14909 16255 14943
rect 20269 14909 20303 14943
rect 24777 14909 24811 14943
rect 13369 14841 13403 14875
rect 13737 14841 13771 14875
rect 15577 14841 15611 14875
rect 19625 14841 19659 14875
rect 12081 14773 12115 14807
rect 12541 14773 12575 14807
rect 15209 14773 15243 14807
rect 18797 14773 18831 14807
rect 20821 14773 20855 14807
rect 8217 14569 8251 14603
rect 8585 14569 8619 14603
rect 9597 14569 9631 14603
rect 10228 14569 10262 14603
rect 12449 14569 12483 14603
rect 21465 14501 21499 14535
rect 6469 14433 6503 14467
rect 11989 14433 12023 14467
rect 13001 14433 13035 14467
rect 14749 14433 14783 14467
rect 14841 14433 14875 14467
rect 16957 14433 16991 14467
rect 17049 14433 17083 14467
rect 21925 14433 21959 14467
rect 22109 14433 22143 14467
rect 23857 14433 23891 14467
rect 9965 14365 9999 14399
rect 13829 14365 13863 14399
rect 14657 14365 14691 14399
rect 15393 14365 15427 14399
rect 20453 14365 20487 14399
rect 22845 14365 22879 14399
rect 25053 14365 25087 14399
rect 6745 14297 6779 14331
rect 12909 14297 12943 14331
rect 16865 14297 16899 14331
rect 17693 14297 17727 14331
rect 12817 14229 12851 14263
rect 13553 14229 13587 14263
rect 14289 14229 14323 14263
rect 16497 14229 16531 14263
rect 20269 14229 20303 14263
rect 21833 14229 21867 14263
rect 24869 14229 24903 14263
rect 12633 14025 12667 14059
rect 13001 14025 13035 14059
rect 19625 14025 19659 14059
rect 20177 14025 20211 14059
rect 8033 13957 8067 13991
rect 10241 13957 10275 13991
rect 15945 13957 15979 13991
rect 19073 13957 19107 13991
rect 19533 13957 19567 13991
rect 22569 13957 22603 13991
rect 7757 13889 7791 13923
rect 10977 13889 11011 13923
rect 20361 13889 20395 13923
rect 21097 13889 21131 13923
rect 22201 13889 22235 13923
rect 25237 13889 25271 13923
rect 9781 13821 9815 13855
rect 11713 13821 11747 13855
rect 13093 13821 13127 13855
rect 13277 13821 13311 13855
rect 13829 13821 13863 13855
rect 15577 13821 15611 13855
rect 16865 13821 16899 13855
rect 17141 13821 17175 13855
rect 18613 13821 18647 13855
rect 22845 13821 22879 13855
rect 23121 13821 23155 13855
rect 24593 13821 24627 13855
rect 20913 13753 20947 13787
rect 22017 13753 22051 13787
rect 12265 13685 12299 13719
rect 14092 13685 14126 13719
rect 18981 13685 19015 13719
rect 25053 13685 25087 13719
rect 8309 13481 8343 13515
rect 8585 13481 8619 13515
rect 9229 13481 9263 13515
rect 10688 13481 10722 13515
rect 13829 13481 13863 13515
rect 17417 13481 17451 13515
rect 21005 13481 21039 13515
rect 24593 13481 24627 13515
rect 6561 13345 6595 13379
rect 9781 13345 9815 13379
rect 10425 13345 10459 13379
rect 13461 13345 13495 13379
rect 14657 13345 14691 13379
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 18797 13345 18831 13379
rect 21649 13345 21683 13379
rect 12633 13277 12667 13311
rect 17877 13277 17911 13311
rect 19441 13277 19475 13311
rect 20821 13277 20855 13311
rect 21373 13277 21407 13311
rect 22845 13277 22879 13311
rect 23857 13277 23891 13311
rect 24777 13277 24811 13311
rect 6837 13209 6871 13243
rect 9597 13209 9631 13243
rect 15577 13209 15611 13243
rect 16221 13209 16255 13243
rect 18613 13209 18647 13243
rect 20269 13209 20303 13243
rect 20729 13209 20763 13243
rect 9689 13141 9723 13175
rect 12173 13141 12207 13175
rect 14841 13141 14875 13175
rect 15209 13141 15243 13175
rect 17969 13141 18003 13175
rect 6653 12937 6687 12971
rect 9045 12937 9079 12971
rect 9413 12937 9447 12971
rect 9505 12937 9539 12971
rect 10425 12937 10459 12971
rect 10793 12937 10827 12971
rect 11897 12937 11931 12971
rect 12265 12937 12299 12971
rect 12633 12937 12667 12971
rect 13093 12937 13127 12971
rect 13829 12937 13863 12971
rect 15393 12937 15427 12971
rect 16129 12937 16163 12971
rect 16865 12937 16899 12971
rect 17325 12937 17359 12971
rect 19993 12937 20027 12971
rect 21097 12937 21131 12971
rect 21189 12937 21223 12971
rect 22017 12937 22051 12971
rect 22845 12937 22879 12971
rect 13001 12869 13035 12903
rect 19257 12869 19291 12903
rect 23397 12869 23431 12903
rect 7021 12801 7055 12835
rect 8217 12801 8251 12835
rect 10885 12801 10919 12835
rect 11529 12801 11563 12835
rect 14197 12801 14231 12835
rect 14289 12801 14323 12835
rect 17233 12801 17267 12835
rect 18245 12801 18279 12835
rect 19165 12801 19199 12835
rect 20177 12801 20211 12835
rect 22201 12801 22235 12835
rect 7113 12733 7147 12767
rect 7205 12733 7239 12767
rect 8309 12733 8343 12767
rect 8493 12733 8527 12767
rect 9597 12733 9631 12767
rect 11069 12733 11103 12767
rect 13185 12733 13219 12767
rect 14381 12733 14415 12767
rect 15485 12733 15519 12767
rect 15669 12733 15703 12767
rect 17509 12733 17543 12767
rect 19441 12733 19475 12767
rect 21373 12733 21407 12767
rect 22477 12733 22511 12767
rect 23121 12733 23155 12767
rect 15025 12665 15059 12699
rect 18061 12665 18095 12699
rect 7849 12597 7883 12631
rect 12081 12597 12115 12631
rect 18797 12597 18831 12631
rect 20729 12597 20763 12631
rect 24869 12597 24903 12631
rect 10241 12393 10275 12427
rect 11437 12393 11471 12427
rect 12633 12393 12667 12427
rect 16313 12393 16347 12427
rect 24593 12393 24627 12427
rect 14289 12325 14323 12359
rect 15393 12325 15427 12359
rect 7389 12257 7423 12291
rect 8217 12257 8251 12291
rect 10793 12257 10827 12291
rect 11989 12257 12023 12291
rect 13277 12257 13311 12291
rect 14841 12257 14875 12291
rect 15577 12257 15611 12291
rect 18705 12257 18739 12291
rect 19993 12257 20027 12291
rect 20453 12257 20487 12291
rect 11805 12189 11839 12223
rect 14749 12189 14783 12223
rect 17325 12189 17359 12223
rect 19533 12189 19567 12223
rect 22845 12189 22879 12223
rect 24777 12189 24811 12223
rect 11897 12121 11931 12155
rect 13093 12121 13127 12155
rect 13737 12121 13771 12155
rect 18153 12121 18187 12155
rect 20729 12121 20763 12155
rect 23857 12121 23891 12155
rect 8953 12053 8987 12087
rect 10609 12053 10643 12087
rect 10701 12053 10735 12087
rect 13001 12053 13035 12087
rect 13921 12053 13955 12087
rect 14657 12053 14691 12087
rect 15761 12053 15795 12087
rect 16681 12053 16715 12087
rect 19625 12053 19659 12087
rect 22201 12053 22235 12087
rect 9045 11849 9079 11883
rect 9873 11849 9907 11883
rect 11897 11849 11931 11883
rect 13093 11849 13127 11883
rect 13461 11849 13495 11883
rect 14289 11849 14323 11883
rect 17325 11849 17359 11883
rect 18061 11849 18095 11883
rect 18429 11849 18463 11883
rect 21373 11849 21407 11883
rect 21649 11849 21683 11883
rect 9505 11781 9539 11815
rect 10241 11781 10275 11815
rect 10333 11781 10367 11815
rect 19349 11781 19383 11815
rect 20085 11781 20119 11815
rect 21281 11781 21315 11815
rect 23305 11781 23339 11815
rect 25145 11781 25179 11815
rect 11621 11713 11655 11747
rect 12265 11713 12299 11747
rect 12357 11713 12391 11747
rect 14657 11713 14691 11747
rect 17233 11713 17267 11747
rect 20269 11713 20303 11747
rect 22293 11713 22327 11747
rect 24133 11713 24167 11747
rect 7297 11645 7331 11679
rect 7573 11645 7607 11679
rect 10425 11645 10459 11679
rect 12449 11645 12483 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 14749 11645 14783 11679
rect 14933 11645 14967 11679
rect 15577 11645 15611 11679
rect 17417 11645 17451 11679
rect 18521 11645 18555 11679
rect 18705 11645 18739 11679
rect 20729 11645 20763 11679
rect 16865 11577 16899 11611
rect 9413 11509 9447 11543
rect 11253 11509 11287 11543
rect 15301 11509 15335 11543
rect 19441 11509 19475 11543
rect 12633 11305 12667 11339
rect 17601 11305 17635 11339
rect 21557 11305 21591 11339
rect 25053 11305 25087 11339
rect 11437 11237 11471 11271
rect 13737 11237 13771 11271
rect 16681 11237 16715 11271
rect 18153 11237 18187 11271
rect 19625 11237 19659 11271
rect 22109 11237 22143 11271
rect 22293 11237 22327 11271
rect 9413 11169 9447 11203
rect 11989 11169 12023 11203
rect 13277 11169 13311 11203
rect 14933 11169 14967 11203
rect 17785 11169 17819 11203
rect 18797 11169 18831 11203
rect 20269 11169 20303 11203
rect 21097 11169 21131 11203
rect 9137 11101 9171 11135
rect 13001 11101 13035 11135
rect 17141 11101 17175 11135
rect 18613 11101 18647 11135
rect 19257 11101 19291 11135
rect 19993 11101 20027 11135
rect 21741 11101 21775 11135
rect 22845 11101 22879 11135
rect 25237 11101 25271 11135
rect 11897 11033 11931 11067
rect 13093 11033 13127 11067
rect 15209 11033 15243 11067
rect 16957 11033 16991 11067
rect 18521 11033 18555 11067
rect 20913 11033 20947 11067
rect 23581 11033 23615 11067
rect 10885 10965 10919 10999
rect 11805 10965 11839 10999
rect 14289 10965 14323 10999
rect 20085 10965 20119 10999
rect 9965 10761 9999 10795
rect 12357 10761 12391 10795
rect 12817 10761 12851 10795
rect 13829 10761 13863 10795
rect 14197 10761 14231 10795
rect 15577 10761 15611 10795
rect 15945 10761 15979 10795
rect 16865 10761 16899 10795
rect 18245 10761 18279 10795
rect 22845 10761 22879 10795
rect 8493 10693 8527 10727
rect 12725 10693 12759 10727
rect 17601 10693 17635 10727
rect 21097 10693 21131 10727
rect 21189 10693 21223 10727
rect 22477 10693 22511 10727
rect 23397 10693 23431 10727
rect 17049 10625 17083 10659
rect 18429 10625 18463 10659
rect 19073 10625 19107 10659
rect 19901 10625 19935 10659
rect 22201 10625 22235 10659
rect 23121 10625 23155 10659
rect 8217 10557 8251 10591
rect 11713 10557 11747 10591
rect 12909 10557 12943 10591
rect 14289 10557 14323 10591
rect 14473 10557 14507 10591
rect 16037 10557 16071 10591
rect 16221 10557 16255 10591
rect 19993 10557 20027 10591
rect 20177 10557 20211 10591
rect 21281 10557 21315 10591
rect 22017 10489 22051 10523
rect 7849 10421 7883 10455
rect 10425 10421 10459 10455
rect 10977 10421 11011 10455
rect 11253 10421 11287 10455
rect 13461 10421 13495 10455
rect 15301 10421 15335 10455
rect 17693 10421 17727 10455
rect 18889 10421 18923 10455
rect 19533 10421 19567 10455
rect 20729 10421 20763 10455
rect 24869 10421 24903 10455
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 12817 10217 12851 10251
rect 14565 10217 14599 10251
rect 15669 10217 15703 10251
rect 22293 10217 22327 10251
rect 24593 10217 24627 10251
rect 23857 10149 23891 10183
rect 9321 10081 9355 10115
rect 12173 10081 12207 10115
rect 13461 10081 13495 10115
rect 14289 10081 14323 10115
rect 15117 10081 15151 10115
rect 18429 10081 18463 10115
rect 18613 10081 18647 10115
rect 23305 10081 23339 10115
rect 23397 10081 23431 10115
rect 13185 10013 13219 10047
rect 14933 10013 14967 10047
rect 20545 10013 20579 10047
rect 23213 10013 23247 10047
rect 24777 10013 24811 10047
rect 9597 9945 9631 9979
rect 11989 9945 12023 9979
rect 16129 9945 16163 9979
rect 16865 9945 16899 9979
rect 19533 9945 19567 9979
rect 20821 9945 20855 9979
rect 12081 9877 12115 9911
rect 13277 9877 13311 9911
rect 13829 9877 13863 9911
rect 15025 9877 15059 9911
rect 16957 9877 16991 9911
rect 17969 9877 18003 9911
rect 18337 9877 18371 9911
rect 18981 9877 19015 9911
rect 19625 9877 19659 9911
rect 19993 9877 20027 9911
rect 20177 9877 20211 9911
rect 22845 9877 22879 9911
rect 13921 9673 13955 9707
rect 24409 9673 24443 9707
rect 14289 9605 14323 9639
rect 16129 9605 16163 9639
rect 11713 9537 11747 9571
rect 15485 9537 15519 9571
rect 20085 9537 20119 9571
rect 25053 9537 25087 9571
rect 11989 9469 12023 9503
rect 13461 9469 13495 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 15577 9469 15611 9503
rect 15761 9469 15795 9503
rect 17325 9469 17359 9503
rect 17601 9469 17635 9503
rect 21281 9469 21315 9503
rect 22017 9469 22051 9503
rect 22661 9469 22695 9503
rect 22937 9469 22971 9503
rect 15117 9401 15151 9435
rect 11345 9333 11379 9367
rect 16405 9333 16439 9367
rect 19073 9333 19107 9367
rect 19441 9333 19475 9367
rect 19809 9333 19843 9367
rect 24869 9333 24903 9367
rect 14289 9129 14323 9163
rect 21373 9129 21407 9163
rect 24593 9129 24627 9163
rect 13001 9061 13035 9095
rect 15945 9061 15979 9095
rect 17233 9061 17267 9095
rect 19349 9061 19383 9095
rect 25053 9061 25087 9095
rect 9137 8993 9171 9027
rect 13645 8993 13679 9027
rect 14841 8993 14875 9027
rect 15301 8993 15335 9027
rect 16497 8993 16531 9027
rect 19625 8993 19659 9027
rect 13461 8925 13495 8959
rect 16313 8925 16347 8959
rect 17693 8925 17727 8959
rect 21925 8925 21959 8959
rect 22661 8925 22695 8959
rect 24777 8925 24811 8959
rect 9413 8857 9447 8891
rect 11161 8857 11195 8891
rect 13369 8857 13403 8891
rect 14657 8857 14691 8891
rect 15485 8857 15519 8891
rect 18705 8857 18739 8891
rect 19901 8857 19935 8891
rect 23857 8857 23891 8891
rect 10885 8789 10919 8823
rect 12725 8789 12759 8823
rect 14749 8789 14783 8823
rect 16405 8789 16439 8823
rect 16957 8789 16991 8823
rect 22017 8789 22051 8823
rect 12909 8585 12943 8619
rect 14473 8585 14507 8619
rect 13921 8517 13955 8551
rect 21281 8517 21315 8551
rect 15117 8449 15151 8483
rect 17417 8449 17451 8483
rect 18245 8449 18279 8483
rect 20269 8449 20303 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 11713 8381 11747 8415
rect 13185 8381 13219 8415
rect 14841 8381 14875 8415
rect 16129 8381 16163 8415
rect 16773 8381 16807 8415
rect 17509 8381 17543 8415
rect 17601 8381 17635 8415
rect 18705 8381 18739 8415
rect 22569 8381 22603 8415
rect 24777 8381 24811 8415
rect 14105 8313 14139 8347
rect 17049 8313 17083 8347
rect 11069 8041 11103 8075
rect 14289 8041 14323 8075
rect 15853 8041 15887 8075
rect 24777 8041 24811 8075
rect 25329 7973 25363 8007
rect 11621 7905 11655 7939
rect 13461 7905 13495 7939
rect 13553 7905 13587 7939
rect 14841 7905 14875 7939
rect 16405 7905 16439 7939
rect 22109 7905 22143 7939
rect 25145 7905 25179 7939
rect 11437 7837 11471 7871
rect 13369 7837 13403 7871
rect 14657 7837 14691 7871
rect 16221 7837 16255 7871
rect 17693 7837 17727 7871
rect 19533 7837 19567 7871
rect 20453 7837 20487 7871
rect 14749 7769 14783 7803
rect 18705 7769 18739 7803
rect 19717 7769 19751 7803
rect 21465 7769 21499 7803
rect 22385 7769 22419 7803
rect 24685 7769 24719 7803
rect 11529 7701 11563 7735
rect 12357 7701 12391 7735
rect 13001 7701 13035 7735
rect 15393 7701 15427 7735
rect 15577 7701 15611 7735
rect 16313 7701 16347 7735
rect 16865 7701 16899 7735
rect 23857 7701 23891 7735
rect 24133 7701 24167 7735
rect 11161 7497 11195 7531
rect 11897 7497 11931 7531
rect 12265 7497 12299 7531
rect 12633 7497 12667 7531
rect 15485 7497 15519 7531
rect 17233 7497 17267 7531
rect 17325 7497 17359 7531
rect 18061 7497 18095 7531
rect 16129 7429 16163 7463
rect 23305 7429 23339 7463
rect 25145 7429 25179 7463
rect 9045 7361 9079 7395
rect 18521 7361 18555 7395
rect 21097 7361 21131 7395
rect 22293 7361 22327 7395
rect 23949 7361 23983 7395
rect 9321 7293 9355 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 13737 7293 13771 7327
rect 14013 7293 14047 7327
rect 17509 7293 17543 7327
rect 20269 7293 20303 7327
rect 21189 7293 21223 7327
rect 21281 7293 21315 7327
rect 16313 7225 16347 7259
rect 10793 7157 10827 7191
rect 16865 7157 16899 7191
rect 17969 7157 18003 7191
rect 18784 7157 18818 7191
rect 20729 7157 20763 7191
rect 12817 6953 12851 6987
rect 10793 6817 10827 6851
rect 12541 6817 12575 6851
rect 14381 6817 14415 6851
rect 19993 6817 20027 6851
rect 20453 6817 20487 6851
rect 24409 6817 24443 6851
rect 25145 6817 25179 6851
rect 13737 6749 13771 6783
rect 14841 6749 14875 6783
rect 15485 6749 15519 6783
rect 17141 6749 17175 6783
rect 20821 6749 20855 6783
rect 22661 6749 22695 6783
rect 24961 6749 24995 6783
rect 11069 6681 11103 6715
rect 16497 6681 16531 6715
rect 17417 6681 17451 6715
rect 19901 6681 19935 6715
rect 22017 6681 22051 6715
rect 23857 6681 23891 6715
rect 13553 6613 13587 6647
rect 14657 6613 14691 6647
rect 18889 6613 18923 6647
rect 19441 6613 19475 6647
rect 19809 6613 19843 6647
rect 24593 6613 24627 6647
rect 25053 6613 25087 6647
rect 10425 6409 10459 6443
rect 11713 6409 11747 6443
rect 13369 6409 13403 6443
rect 17325 6409 17359 6443
rect 23765 6409 23799 6443
rect 12173 6341 12207 6375
rect 12725 6341 12759 6375
rect 22293 6341 22327 6375
rect 24317 6341 24351 6375
rect 10793 6273 10827 6307
rect 12081 6273 12115 6307
rect 13737 6273 13771 6307
rect 15117 6273 15151 6307
rect 17233 6273 17267 6307
rect 17969 6273 18003 6307
rect 18245 6273 18279 6307
rect 20269 6273 20303 6307
rect 22017 6273 22051 6307
rect 25053 6273 25087 6307
rect 10885 6205 10919 6239
rect 10977 6205 11011 6239
rect 12265 6205 12299 6239
rect 13001 6205 13035 6239
rect 13829 6205 13863 6239
rect 13921 6205 13955 6239
rect 16129 6205 16163 6239
rect 17417 6205 17451 6239
rect 19441 6205 19475 6239
rect 21281 6205 21315 6239
rect 25237 6205 25271 6239
rect 16865 6137 16899 6171
rect 24501 6137 24535 6171
rect 14381 6069 14415 6103
rect 11805 5865 11839 5899
rect 13553 5865 13587 5899
rect 14197 5865 14231 5899
rect 14749 5865 14783 5899
rect 17693 5865 17727 5899
rect 24133 5865 24167 5899
rect 25145 5865 25179 5899
rect 12909 5797 12943 5831
rect 24869 5797 24903 5831
rect 10333 5729 10367 5763
rect 12265 5729 12299 5763
rect 15393 5729 15427 5763
rect 18613 5729 18647 5763
rect 18797 5729 18831 5763
rect 19901 5729 19935 5763
rect 22201 5729 22235 5763
rect 23673 5729 23707 5763
rect 10057 5661 10091 5695
rect 13093 5661 13127 5695
rect 13737 5661 13771 5695
rect 15945 5661 15979 5695
rect 19625 5661 19659 5695
rect 21281 5661 21315 5695
rect 23581 5661 23615 5695
rect 24685 5661 24719 5695
rect 25329 5661 25363 5695
rect 14473 5593 14507 5627
rect 15209 5593 15243 5627
rect 16221 5593 16255 5627
rect 18521 5593 18555 5627
rect 23489 5593 23523 5627
rect 15117 5525 15151 5559
rect 18153 5525 18187 5559
rect 23121 5525 23155 5559
rect 11529 5321 11563 5355
rect 12541 5321 12575 5355
rect 14933 5321 14967 5355
rect 21373 5321 21407 5355
rect 13461 5253 13495 5287
rect 10609 5185 10643 5219
rect 12725 5185 12759 5219
rect 16681 5185 16715 5219
rect 16865 5185 16899 5219
rect 17049 5185 17083 5219
rect 17417 5185 17451 5219
rect 19625 5185 19659 5219
rect 22201 5185 22235 5219
rect 24041 5185 24075 5219
rect 10333 5117 10367 5151
rect 11805 5117 11839 5151
rect 12081 5117 12115 5151
rect 13185 5117 13219 5151
rect 15485 5117 15519 5151
rect 15761 5117 15795 5151
rect 19901 5117 19935 5151
rect 22937 5117 22971 5151
rect 24317 5117 24351 5151
rect 6101 4981 6135 5015
rect 7205 4981 7239 5015
rect 18705 4981 18739 5015
rect 18981 4777 19015 4811
rect 21281 4777 21315 4811
rect 24777 4777 24811 4811
rect 1593 4709 1627 4743
rect 16865 4709 16899 4743
rect 5089 4641 5123 4675
rect 9689 4641 9723 4675
rect 9965 4641 9999 4675
rect 14473 4641 14507 4675
rect 15117 4641 15151 4675
rect 15393 4641 15427 4675
rect 19533 4641 19567 4675
rect 22201 4641 22235 4675
rect 1777 4573 1811 4607
rect 2789 4573 2823 4607
rect 3433 4573 3467 4607
rect 3985 4573 4019 4607
rect 7849 4573 7883 4607
rect 11069 4573 11103 4607
rect 11345 4573 11379 4607
rect 12541 4573 12575 4607
rect 14197 4573 14231 4607
rect 17509 4573 17543 4607
rect 21925 4573 21959 4607
rect 24685 4573 24719 4607
rect 25145 4573 25179 4607
rect 4629 4505 4663 4539
rect 5365 4505 5399 4539
rect 7113 4505 7147 4539
rect 13277 4505 13311 4539
rect 18521 4505 18555 4539
rect 19809 4505 19843 4539
rect 23673 4505 23707 4539
rect 24133 4505 24167 4539
rect 25329 4505 25363 4539
rect 7481 4437 7515 4471
rect 7757 4437 7791 4471
rect 8033 4437 8067 4471
rect 8309 4437 8343 4471
rect 8585 4437 8619 4471
rect 8769 4437 8803 4471
rect 23765 4437 23799 4471
rect 7205 4233 7239 4267
rect 10011 4233 10045 4267
rect 21557 4233 21591 4267
rect 22109 4233 22143 4267
rect 22753 4233 22787 4267
rect 14197 4165 14231 4199
rect 1593 4097 1627 4131
rect 2881 4097 2915 4131
rect 4353 4097 4387 4131
rect 4997 4097 5031 4131
rect 5365 4097 5399 4131
rect 6009 4097 6043 4131
rect 6745 4097 6779 4131
rect 7389 4097 7423 4131
rect 8033 4097 8067 4131
rect 8677 4097 8711 4131
rect 9321 4097 9355 4131
rect 11069 4097 11103 4131
rect 11345 4097 11379 4131
rect 12265 4097 12299 4131
rect 13921 4097 13955 4131
rect 16313 4097 16347 4131
rect 17049 4097 17083 4131
rect 18889 4097 18923 4131
rect 20913 4097 20947 4131
rect 22293 4097 22327 4131
rect 23581 4097 23615 4131
rect 24225 4097 24259 4131
rect 24685 4097 24719 4131
rect 3249 4029 3283 4063
rect 9781 4029 9815 4063
rect 13277 4029 13311 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 21005 4029 21039 4063
rect 21189 4029 21223 4063
rect 2237 3961 2271 3995
rect 3341 3961 3375 3995
rect 4169 3961 4203 3995
rect 6561 3961 6595 3995
rect 7849 3961 7883 3995
rect 8493 3961 8527 3995
rect 9137 3961 9171 3995
rect 15669 3961 15703 3995
rect 23397 3961 23431 3995
rect 2697 3893 2731 3927
rect 3525 3893 3559 3927
rect 3893 3893 3927 3927
rect 4813 3893 4847 3927
rect 5549 3893 5583 3927
rect 5825 3893 5859 3927
rect 10885 3893 10919 3927
rect 11621 3893 11655 3927
rect 11805 3893 11839 3927
rect 16129 3893 16163 3927
rect 20545 3893 20579 3927
rect 24041 3893 24075 3927
rect 25329 3893 25363 3927
rect 2605 3689 2639 3723
rect 3065 3689 3099 3723
rect 4261 3689 4295 3723
rect 7021 3689 7055 3723
rect 7481 3689 7515 3723
rect 8401 3689 8435 3723
rect 9137 3689 9171 3723
rect 9781 3689 9815 3723
rect 10425 3689 10459 3723
rect 18291 3689 18325 3723
rect 22937 3689 22971 3723
rect 24041 3689 24075 3723
rect 3985 3553 4019 3587
rect 4905 3553 4939 3587
rect 5181 3553 5215 3587
rect 6101 3553 6135 3587
rect 11069 3553 11103 3587
rect 12817 3553 12851 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 18061 3553 18095 3587
rect 21741 3553 21775 3587
rect 1961 3485 1995 3519
rect 3249 3485 3283 3519
rect 3617 3485 3651 3519
rect 4445 3485 4479 3519
rect 6377 3485 6411 3519
rect 7665 3485 7699 3519
rect 8585 3485 8619 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 10609 3485 10643 3519
rect 11345 3485 11379 3519
rect 12449 3485 12483 3519
rect 14473 3485 14507 3519
rect 16313 3485 16347 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 23397 3485 23431 3519
rect 24593 3485 24627 3519
rect 8125 3417 8159 3451
rect 20361 3417 20395 3451
rect 1501 3349 1535 3383
rect 25237 3349 25271 3383
rect 7297 3145 7331 3179
rect 9413 3145 9447 3179
rect 10333 3145 10367 3179
rect 21281 3145 21315 3179
rect 22937 3145 22971 3179
rect 23673 3145 23707 3179
rect 24225 3145 24259 3179
rect 24593 3145 24627 3179
rect 22293 3077 22327 3111
rect 22845 3077 22879 3111
rect 25053 3077 25087 3111
rect 2421 3009 2455 3043
rect 3433 3009 3467 3043
rect 3709 3009 3743 3043
rect 5457 3009 5491 3043
rect 6653 3009 6687 3043
rect 7849 3009 7883 3043
rect 9873 3009 9907 3043
rect 10517 3009 10551 3043
rect 11161 3009 11195 3043
rect 11713 3009 11747 3043
rect 13185 3009 13219 3043
rect 14841 3009 14875 3043
rect 17049 3009 17083 3043
rect 18889 3009 18923 3043
rect 20637 3009 20671 3043
rect 22109 3009 22143 3043
rect 23581 3009 23615 3043
rect 24777 3009 24811 3043
rect 25237 3009 25271 3043
rect 1777 2941 1811 2975
rect 2145 2941 2179 2975
rect 4721 2941 4755 2975
rect 5181 2941 5215 2975
rect 8125 2941 8159 2975
rect 9229 2941 9263 2975
rect 11989 2941 12023 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 24041 2941 24075 2975
rect 1685 2873 1719 2907
rect 9045 2873 9079 2907
rect 9689 2873 9723 2907
rect 4905 2805 4939 2839
rect 10977 2805 11011 2839
rect 20729 2805 20763 2839
rect 4629 2601 4663 2635
rect 7297 2601 7331 2635
rect 8401 2601 8435 2635
rect 18705 2601 18739 2635
rect 16313 2533 16347 2567
rect 2329 2465 2363 2499
rect 2605 2465 2639 2499
rect 2881 2465 2915 2499
rect 5457 2465 5491 2499
rect 14197 2465 14231 2499
rect 14933 2465 14967 2499
rect 16129 2465 16163 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 25237 2465 25271 2499
rect 1869 2397 1903 2431
rect 3985 2397 4019 2431
rect 5181 2397 5215 2431
rect 6653 2397 6687 2431
rect 7941 2397 7975 2431
rect 8585 2397 8619 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 14473 2397 14507 2431
rect 16865 2397 16899 2431
rect 18889 2397 18923 2431
rect 19625 2397 19659 2431
rect 21465 2397 21499 2431
rect 22017 2397 22051 2431
rect 22937 2397 22971 2431
rect 24593 2397 24627 2431
rect 10977 2329 11011 2363
rect 13277 2329 13311 2363
rect 23857 2329 23891 2363
rect 1685 2261 1719 2295
rect 7757 2261 7791 2295
rect 9137 2261 9171 2295
rect 11713 2261 11747 2295
rect 21281 2261 21315 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 16206 54272 16212 54324
rect 16264 54312 16270 54324
rect 16393 54315 16451 54321
rect 16393 54312 16405 54315
rect 16264 54284 16405 54312
rect 16264 54272 16270 54284
rect 16393 54281 16405 54284
rect 16439 54281 16451 54315
rect 16393 54275 16451 54281
rect 16500 54284 18184 54312
rect 8570 54204 8576 54256
rect 8628 54244 8634 54256
rect 16500 54244 16528 54284
rect 8628 54216 16528 54244
rect 8628 54204 8634 54216
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 4062 54176 4068 54188
rect 2271 54148 4068 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4062 54136 4068 54148
rect 4120 54136 4126 54188
rect 4798 54136 4804 54188
rect 4856 54136 4862 54188
rect 7374 54136 7380 54188
rect 7432 54136 7438 54188
rect 9582 54136 9588 54188
rect 9640 54136 9646 54188
rect 11698 54136 11704 54188
rect 11756 54176 11762 54188
rect 12161 54179 12219 54185
rect 12161 54176 12173 54179
rect 11756 54148 12173 54176
rect 11756 54136 11762 54148
rect 12161 54145 12173 54148
rect 12207 54145 12219 54179
rect 12161 54139 12219 54145
rect 14458 54136 14464 54188
rect 14516 54136 14522 54188
rect 14826 54136 14832 54188
rect 14884 54176 14890 54188
rect 15013 54179 15071 54185
rect 15013 54176 15025 54179
rect 14884 54148 15025 54176
rect 14884 54136 14890 54148
rect 15013 54145 15025 54148
rect 15059 54176 15071 54179
rect 15933 54179 15991 54185
rect 15933 54176 15945 54179
rect 15059 54148 15945 54176
rect 15059 54145 15071 54148
rect 15013 54139 15071 54145
rect 15933 54145 15945 54148
rect 15979 54145 15991 54179
rect 15933 54139 15991 54145
rect 16206 54136 16212 54188
rect 16264 54176 16270 54188
rect 16853 54179 16911 54185
rect 16853 54176 16865 54179
rect 16264 54148 16865 54176
rect 16264 54136 16270 54148
rect 16853 54145 16865 54148
rect 16899 54145 16911 54179
rect 16853 54139 16911 54145
rect 17954 54136 17960 54188
rect 18012 54136 18018 54188
rect 2406 54068 2412 54120
rect 2464 54108 2470 54120
rect 2501 54111 2559 54117
rect 2501 54108 2513 54111
rect 2464 54080 2513 54108
rect 2464 54068 2470 54080
rect 2501 54077 2513 54080
rect 2547 54077 2559 54111
rect 2501 54071 2559 54077
rect 5166 54068 5172 54120
rect 5224 54068 5230 54120
rect 7834 54068 7840 54120
rect 7892 54068 7898 54120
rect 9306 54068 9312 54120
rect 9364 54108 9370 54120
rect 9861 54111 9919 54117
rect 9861 54108 9873 54111
rect 9364 54080 9873 54108
rect 9364 54068 9370 54080
rect 9861 54077 9873 54080
rect 9907 54077 9919 54111
rect 9861 54071 9919 54077
rect 12342 54068 12348 54120
rect 12400 54108 12406 54120
rect 12621 54111 12679 54117
rect 12621 54108 12633 54111
rect 12400 54080 12633 54108
rect 12400 54068 12406 54080
rect 12621 54077 12633 54080
rect 12667 54077 12679 54111
rect 18156 54108 18184 54284
rect 18966 54272 18972 54324
rect 19024 54272 19030 54324
rect 18984 54176 19012 54272
rect 25317 54247 25375 54253
rect 25317 54244 25329 54247
rect 23400 54216 25329 54244
rect 19429 54179 19487 54185
rect 19429 54176 19441 54179
rect 18984 54148 19441 54176
rect 19429 54145 19441 54148
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 21269 54179 21327 54185
rect 21269 54176 21281 54179
rect 20772 54148 21281 54176
rect 20772 54136 20778 54148
rect 21269 54145 21281 54148
rect 21315 54145 21327 54179
rect 21269 54139 21327 54145
rect 21726 54136 21732 54188
rect 21784 54176 21790 54188
rect 23400 54185 23428 54216
rect 25317 54213 25329 54216
rect 25363 54213 25375 54247
rect 25317 54207 25375 54213
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21784 54148 22017 54176
rect 21784 54136 21790 54148
rect 22005 54145 22017 54148
rect 22051 54176 22063 54179
rect 22557 54179 22615 54185
rect 22557 54176 22569 54179
rect 22051 54148 22569 54176
rect 22051 54145 22063 54148
rect 22005 54139 22063 54145
rect 22557 54145 22569 54148
rect 22603 54145 22615 54179
rect 22557 54139 22615 54145
rect 23385 54179 23443 54185
rect 23385 54145 23397 54179
rect 23431 54145 23443 54179
rect 23385 54139 23443 54145
rect 24673 54179 24731 54185
rect 24673 54145 24685 54179
rect 24719 54176 24731 54179
rect 25866 54176 25872 54188
rect 24719 54148 25872 54176
rect 24719 54145 24731 54148
rect 24673 54139 24731 54145
rect 19705 54111 19763 54117
rect 19705 54108 19717 54111
rect 18156 54080 19717 54108
rect 12621 54071 12679 54077
rect 19705 54077 19717 54080
rect 19751 54077 19763 54111
rect 19705 54071 19763 54077
rect 23109 54111 23167 54117
rect 23109 54077 23121 54111
rect 23155 54108 23167 54111
rect 24688 54108 24716 54139
rect 25866 54136 25872 54148
rect 25924 54136 25930 54188
rect 23155 54080 24716 54108
rect 23155 54077 23167 54080
rect 23109 54071 23167 54077
rect 16758 54000 16764 54052
rect 16816 54040 16822 54052
rect 16816 54012 18736 54040
rect 16816 54000 16822 54012
rect 13538 53932 13544 53984
rect 13596 53972 13602 53984
rect 14277 53975 14335 53981
rect 14277 53972 14289 53975
rect 13596 53944 14289 53972
rect 13596 53932 13602 53944
rect 14277 53941 14289 53944
rect 14323 53941 14335 53975
rect 14277 53935 14335 53941
rect 15562 53932 15568 53984
rect 15620 53972 15626 53984
rect 15657 53975 15715 53981
rect 15657 53972 15669 53975
rect 15620 53944 15669 53972
rect 15620 53932 15626 53944
rect 15657 53941 15669 53944
rect 15703 53941 15715 53975
rect 15657 53935 15715 53941
rect 17034 53932 17040 53984
rect 17092 53972 17098 53984
rect 17497 53975 17555 53981
rect 17497 53972 17509 53975
rect 17092 53944 17509 53972
rect 17092 53932 17098 53944
rect 17497 53941 17509 53944
rect 17543 53941 17555 53975
rect 17497 53935 17555 53941
rect 18598 53932 18604 53984
rect 18656 53932 18662 53984
rect 18708 53972 18736 54012
rect 18782 54000 18788 54052
rect 18840 54040 18846 54052
rect 22189 54043 22247 54049
rect 22189 54040 22201 54043
rect 18840 54012 22201 54040
rect 18840 54000 18846 54012
rect 22189 54009 22201 54012
rect 22235 54009 22247 54043
rect 22189 54003 22247 54009
rect 20901 53975 20959 53981
rect 20901 53972 20913 53975
rect 18708 53944 20913 53972
rect 20901 53941 20913 53944
rect 20947 53941 20959 53975
rect 20901 53935 20959 53941
rect 24029 53975 24087 53981
rect 24029 53941 24041 53975
rect 24075 53972 24087 53975
rect 24670 53972 24676 53984
rect 24075 53944 24676 53972
rect 24075 53941 24087 53944
rect 24029 53935 24087 53941
rect 24670 53932 24676 53944
rect 24728 53932 24734 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 13446 53728 13452 53780
rect 13504 53768 13510 53780
rect 13817 53771 13875 53777
rect 13817 53768 13829 53771
rect 13504 53740 13829 53768
rect 13504 53728 13510 53740
rect 13817 53737 13829 53740
rect 13863 53737 13875 53771
rect 13817 53731 13875 53737
rect 10686 53660 10692 53712
rect 10744 53660 10750 53712
rect 1026 53592 1032 53644
rect 1084 53632 1090 53644
rect 2041 53635 2099 53641
rect 2041 53632 2053 53635
rect 1084 53604 2053 53632
rect 1084 53592 1090 53604
rect 2041 53601 2053 53604
rect 2087 53601 2099 53635
rect 2041 53595 2099 53601
rect 3786 53592 3792 53644
rect 3844 53632 3850 53644
rect 4433 53635 4491 53641
rect 4433 53632 4445 53635
rect 3844 53604 4445 53632
rect 3844 53592 3850 53604
rect 4433 53601 4445 53604
rect 4479 53601 4491 53635
rect 4433 53595 4491 53601
rect 6546 53592 6552 53644
rect 6604 53632 6610 53644
rect 7101 53635 7159 53641
rect 7101 53632 7113 53635
rect 6604 53604 7113 53632
rect 6604 53592 6610 53604
rect 7101 53601 7113 53604
rect 7147 53601 7159 53635
rect 10704 53632 10732 53660
rect 11241 53635 11299 53641
rect 11241 53632 11253 53635
rect 10704 53604 11253 53632
rect 7101 53595 7159 53601
rect 11241 53601 11253 53604
rect 11287 53601 11299 53635
rect 11241 53595 11299 53601
rect 1765 53567 1823 53573
rect 1765 53533 1777 53567
rect 1811 53533 1823 53567
rect 1765 53527 1823 53533
rect 1780 53496 1808 53527
rect 4154 53524 4160 53576
rect 4212 53524 4218 53576
rect 6825 53567 6883 53573
rect 6825 53533 6837 53567
rect 6871 53564 6883 53567
rect 7834 53564 7840 53576
rect 6871 53536 7840 53564
rect 6871 53533 6883 53536
rect 6825 53527 6883 53533
rect 7834 53524 7840 53536
rect 7892 53524 7898 53576
rect 10686 53524 10692 53576
rect 10744 53564 10750 53576
rect 10781 53567 10839 53573
rect 10781 53564 10793 53567
rect 10744 53536 10793 53564
rect 10744 53524 10750 53536
rect 10781 53533 10793 53536
rect 10827 53533 10839 53567
rect 13832 53564 13860 53731
rect 14458 53728 14464 53780
rect 14516 53768 14522 53780
rect 14921 53771 14979 53777
rect 14921 53768 14933 53771
rect 14516 53740 14933 53768
rect 14516 53728 14522 53740
rect 14921 53737 14933 53740
rect 14967 53737 14979 53771
rect 14921 53731 14979 53737
rect 17862 53728 17868 53780
rect 17920 53768 17926 53780
rect 18141 53771 18199 53777
rect 18141 53768 18153 53771
rect 17920 53740 18153 53768
rect 17920 53728 17926 53740
rect 18141 53737 18153 53740
rect 18187 53737 18199 53771
rect 18141 53731 18199 53737
rect 23290 53592 23296 53644
rect 23348 53632 23354 53644
rect 23348 53604 23796 53632
rect 23348 53592 23354 53604
rect 14277 53567 14335 53573
rect 14277 53564 14289 53567
rect 13832 53536 14289 53564
rect 10781 53527 10839 53533
rect 14277 53533 14289 53536
rect 14323 53533 14335 53567
rect 14277 53527 14335 53533
rect 15562 53524 15568 53576
rect 15620 53524 15626 53576
rect 17034 53524 17040 53576
rect 17092 53524 17098 53576
rect 17865 53567 17923 53573
rect 17865 53533 17877 53567
rect 17911 53564 17923 53567
rect 18598 53564 18604 53576
rect 17911 53536 18604 53564
rect 17911 53533 17923 53536
rect 17865 53527 17923 53533
rect 18598 53524 18604 53536
rect 18656 53524 18662 53576
rect 22278 53524 22284 53576
rect 22336 53524 22342 53576
rect 23109 53567 23167 53573
rect 23109 53533 23121 53567
rect 23155 53564 23167 53567
rect 23382 53564 23388 53576
rect 23155 53536 23388 53564
rect 23155 53533 23167 53536
rect 23109 53527 23167 53533
rect 23382 53524 23388 53536
rect 23440 53524 23446 53576
rect 23768 53573 23796 53604
rect 23753 53567 23811 53573
rect 23753 53533 23765 53567
rect 23799 53533 23811 53567
rect 23753 53527 23811 53533
rect 24670 53524 24676 53576
rect 24728 53524 24734 53576
rect 5534 53496 5540 53508
rect 1780 53468 5540 53496
rect 5534 53456 5540 53468
rect 5592 53456 5598 53508
rect 21450 53456 21456 53508
rect 21508 53496 21514 53508
rect 21508 53468 22600 53496
rect 21508 53456 21514 53468
rect 14734 53388 14740 53440
rect 14792 53428 14798 53440
rect 15381 53431 15439 53437
rect 15381 53428 15393 53431
rect 14792 53400 15393 53428
rect 14792 53388 14798 53400
rect 15381 53397 15393 53400
rect 15427 53397 15439 53431
rect 15381 53391 15439 53397
rect 15654 53388 15660 53440
rect 15712 53428 15718 53440
rect 16853 53431 16911 53437
rect 16853 53428 16865 53431
rect 15712 53400 16865 53428
rect 15712 53388 15718 53400
rect 16853 53397 16865 53400
rect 16899 53397 16911 53431
rect 16853 53391 16911 53397
rect 17678 53388 17684 53440
rect 17736 53388 17742 53440
rect 19978 53388 19984 53440
rect 20036 53428 20042 53440
rect 22465 53431 22523 53437
rect 22465 53428 22477 53431
rect 20036 53400 22477 53428
rect 20036 53388 20042 53400
rect 22465 53397 22477 53400
rect 22511 53397 22523 53431
rect 22572 53428 22600 53468
rect 23201 53431 23259 53437
rect 23201 53428 23213 53431
rect 22572 53400 23213 53428
rect 22465 53391 22523 53397
rect 23201 53397 23213 53400
rect 23247 53397 23259 53431
rect 23201 53391 23259 53397
rect 23934 53388 23940 53440
rect 23992 53388 23998 53440
rect 24578 53388 24584 53440
rect 24636 53428 24642 53440
rect 25317 53431 25375 53437
rect 25317 53428 25329 53431
rect 24636 53400 25329 53428
rect 24636 53388 24642 53400
rect 25317 53397 25329 53400
rect 25363 53397 25375 53431
rect 25317 53391 25375 53397
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 4062 53184 4068 53236
rect 4120 53224 4126 53236
rect 5169 53227 5227 53233
rect 5169 53224 5181 53227
rect 4120 53196 5181 53224
rect 4120 53184 4126 53196
rect 5169 53193 5181 53196
rect 5215 53193 5227 53227
rect 5169 53187 5227 53193
rect 23290 53184 23296 53236
rect 23348 53184 23354 53236
rect 23382 53184 23388 53236
rect 23440 53184 23446 53236
rect 24762 53184 24768 53236
rect 24820 53224 24826 53236
rect 25041 53227 25099 53233
rect 25041 53224 25053 53227
rect 24820 53196 25053 53224
rect 24820 53184 24826 53196
rect 25041 53193 25053 53196
rect 25087 53193 25099 53227
rect 25041 53187 25099 53193
rect 25314 53184 25320 53236
rect 25372 53184 25378 53236
rect 24780 53156 24808 53184
rect 23768 53128 24808 53156
rect 5353 53091 5411 53097
rect 5353 53057 5365 53091
rect 5399 53088 5411 53091
rect 7742 53088 7748 53100
rect 5399 53060 7748 53088
rect 5399 53057 5411 53060
rect 5353 53051 5411 53057
rect 7742 53048 7748 53060
rect 7800 53048 7806 53100
rect 23768 53097 23796 53128
rect 23753 53091 23811 53097
rect 23753 53057 23765 53091
rect 23799 53057 23811 53091
rect 23753 53051 23811 53057
rect 24489 53091 24547 53097
rect 24489 53057 24501 53091
rect 24535 53088 24547 53091
rect 25332 53088 25360 53184
rect 24535 53060 25360 53088
rect 24535 53057 24547 53060
rect 24489 53051 24547 53057
rect 22278 52980 22284 53032
rect 22336 53020 22342 53032
rect 22741 53023 22799 53029
rect 22741 53020 22753 53023
rect 22336 52992 22753 53020
rect 22336 52980 22342 52992
rect 22741 52989 22753 52992
rect 22787 53020 22799 53023
rect 24854 53020 24860 53032
rect 22787 52992 24860 53020
rect 22787 52989 22799 52992
rect 22741 52983 22799 52989
rect 24854 52980 24860 52992
rect 24912 52980 24918 53032
rect 25498 52912 25504 52964
rect 25556 52912 25562 52964
rect 23658 52844 23664 52896
rect 23716 52884 23722 52896
rect 23937 52887 23995 52893
rect 23937 52884 23949 52887
rect 23716 52856 23949 52884
rect 23716 52844 23722 52856
rect 23937 52853 23949 52856
rect 23983 52853 23995 52887
rect 23937 52847 23995 52853
rect 24670 52844 24676 52896
rect 24728 52844 24734 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 4154 52640 4160 52692
rect 4212 52680 4218 52692
rect 6549 52683 6607 52689
rect 6549 52680 6561 52683
rect 4212 52652 6561 52680
rect 4212 52640 4218 52652
rect 6549 52649 6561 52652
rect 6595 52649 6607 52683
rect 6549 52643 6607 52649
rect 24486 52640 24492 52692
rect 24544 52640 24550 52692
rect 23842 52572 23848 52624
rect 23900 52612 23906 52624
rect 23937 52615 23995 52621
rect 23937 52612 23949 52615
rect 23900 52584 23949 52612
rect 23900 52572 23906 52584
rect 23937 52581 23949 52584
rect 23983 52581 23995 52615
rect 23937 52575 23995 52581
rect 6733 52479 6791 52485
rect 6733 52445 6745 52479
rect 6779 52476 6791 52479
rect 9490 52476 9496 52488
rect 6779 52448 9496 52476
rect 6779 52445 6791 52448
rect 6733 52439 6791 52445
rect 9490 52436 9496 52448
rect 9548 52436 9554 52488
rect 23753 52479 23811 52485
rect 23753 52445 23765 52479
rect 23799 52476 23811 52479
rect 24486 52476 24492 52488
rect 23799 52448 24492 52476
rect 23799 52445 23811 52448
rect 23753 52439 23811 52445
rect 24486 52436 24492 52448
rect 24544 52436 24550 52488
rect 25317 52479 25375 52485
rect 25317 52445 25329 52479
rect 25363 52476 25375 52479
rect 25958 52476 25964 52488
rect 25363 52448 25964 52476
rect 25363 52445 25375 52448
rect 25317 52439 25375 52445
rect 25958 52436 25964 52448
rect 26016 52436 26022 52488
rect 24946 52368 24952 52420
rect 25004 52368 25010 52420
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 24121 52139 24179 52145
rect 24121 52105 24133 52139
rect 24167 52136 24179 52139
rect 24946 52136 24952 52148
rect 24167 52108 24952 52136
rect 24167 52105 24179 52108
rect 24121 52099 24179 52105
rect 24946 52096 24952 52108
rect 25004 52096 25010 52148
rect 24578 51960 24584 52012
rect 24636 51960 24642 52012
rect 25041 52003 25099 52009
rect 25041 51969 25053 52003
rect 25087 52000 25099 52003
rect 25498 52000 25504 52012
rect 25087 51972 25504 52000
rect 25087 51969 25099 51972
rect 25041 51963 25099 51969
rect 25498 51960 25504 51972
rect 25556 51960 25562 52012
rect 24397 51799 24455 51805
rect 24397 51765 24409 51799
rect 24443 51796 24455 51799
rect 24578 51796 24584 51808
rect 24443 51768 24584 51796
rect 24443 51765 24455 51768
rect 24397 51759 24455 51765
rect 24578 51756 24584 51768
rect 24636 51756 24642 51808
rect 25222 51756 25228 51808
rect 25280 51756 25286 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 7374 51552 7380 51604
rect 7432 51592 7438 51604
rect 8297 51595 8355 51601
rect 8297 51592 8309 51595
rect 7432 51564 8309 51592
rect 7432 51552 7438 51564
rect 8297 51561 8309 51564
rect 8343 51561 8355 51595
rect 8297 51555 8355 51561
rect 7834 51484 7840 51536
rect 7892 51524 7898 51536
rect 9217 51527 9275 51533
rect 9217 51524 9229 51527
rect 7892 51496 9229 51524
rect 7892 51484 7898 51496
rect 9217 51493 9229 51496
rect 9263 51493 9275 51527
rect 9217 51487 9275 51493
rect 4798 51348 4804 51400
rect 4856 51388 4862 51400
rect 7837 51391 7895 51397
rect 7837 51388 7849 51391
rect 4856 51360 7849 51388
rect 4856 51348 4862 51360
rect 7837 51357 7849 51360
rect 7883 51357 7895 51391
rect 7837 51351 7895 51357
rect 8478 51348 8484 51400
rect 8536 51348 8542 51400
rect 9401 51391 9459 51397
rect 9401 51357 9413 51391
rect 9447 51388 9459 51391
rect 10502 51388 10508 51400
rect 9447 51360 10508 51388
rect 9447 51357 9459 51360
rect 9401 51351 9459 51357
rect 10502 51348 10508 51360
rect 10560 51348 10566 51400
rect 7653 51323 7711 51329
rect 7653 51289 7665 51323
rect 7699 51320 7711 51323
rect 10778 51320 10784 51332
rect 7699 51292 10784 51320
rect 7699 51289 7711 51292
rect 7653 51283 7711 51289
rect 10778 51280 10784 51292
rect 10836 51280 10842 51332
rect 24581 51323 24639 51329
rect 24581 51289 24593 51323
rect 24627 51320 24639 51323
rect 24946 51320 24952 51332
rect 24627 51292 24952 51320
rect 24627 51289 24639 51292
rect 24581 51283 24639 51289
rect 24946 51280 24952 51292
rect 25004 51280 25010 51332
rect 25317 51323 25375 51329
rect 25317 51289 25329 51323
rect 25363 51320 25375 51323
rect 25774 51320 25780 51332
rect 25363 51292 25780 51320
rect 25363 51289 25375 51292
rect 25317 51283 25375 51289
rect 25774 51280 25780 51292
rect 25832 51280 25838 51332
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 24581 50915 24639 50921
rect 24581 50881 24593 50915
rect 24627 50912 24639 50915
rect 24949 50915 25007 50921
rect 24949 50912 24961 50915
rect 24627 50884 24961 50912
rect 24627 50881 24639 50884
rect 24581 50875 24639 50881
rect 24949 50881 24961 50884
rect 24995 50912 25007 50915
rect 25038 50912 25044 50924
rect 24995 50884 25044 50912
rect 24995 50881 25007 50884
rect 24949 50875 25007 50881
rect 25038 50872 25044 50884
rect 25096 50872 25102 50924
rect 24946 50668 24952 50720
rect 25004 50708 25010 50720
rect 25041 50711 25099 50717
rect 25041 50708 25053 50711
rect 25004 50680 25053 50708
rect 25004 50668 25010 50680
rect 25041 50677 25053 50680
rect 25087 50677 25099 50711
rect 25041 50671 25099 50677
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 5534 50464 5540 50516
rect 5592 50504 5598 50516
rect 7837 50507 7895 50513
rect 7837 50504 7849 50507
rect 5592 50476 7849 50504
rect 5592 50464 5598 50476
rect 7837 50473 7849 50476
rect 7883 50504 7895 50507
rect 8386 50504 8392 50516
rect 7883 50476 8392 50504
rect 7883 50473 7895 50476
rect 7837 50467 7895 50473
rect 8386 50464 8392 50476
rect 8444 50464 8450 50516
rect 9582 50464 9588 50516
rect 9640 50464 9646 50516
rect 7742 50396 7748 50448
rect 7800 50436 7806 50448
rect 8021 50439 8079 50445
rect 8021 50436 8033 50439
rect 7800 50408 8033 50436
rect 7800 50396 7806 50408
rect 8021 50405 8033 50408
rect 8067 50405 8079 50439
rect 8021 50399 8079 50405
rect 8389 50371 8447 50377
rect 8389 50337 8401 50371
rect 8435 50368 8447 50371
rect 8570 50368 8576 50380
rect 8435 50340 8576 50368
rect 8435 50337 8447 50340
rect 8389 50331 8447 50337
rect 7561 50303 7619 50309
rect 7561 50269 7573 50303
rect 7607 50300 7619 50303
rect 8404 50300 8432 50331
rect 8570 50328 8576 50340
rect 8628 50328 8634 50380
rect 7607 50272 8432 50300
rect 7607 50269 7619 50272
rect 7561 50263 7619 50269
rect 24578 50260 24584 50312
rect 24636 50260 24642 50312
rect 9493 50235 9551 50241
rect 9493 50201 9505 50235
rect 9539 50232 9551 50235
rect 9582 50232 9588 50244
rect 9539 50204 9588 50232
rect 9539 50201 9551 50204
rect 9493 50195 9551 50201
rect 9582 50192 9588 50204
rect 9640 50192 9646 50244
rect 23382 50124 23388 50176
rect 23440 50164 23446 50176
rect 25225 50167 25283 50173
rect 25225 50164 25237 50167
rect 23440 50136 25237 50164
rect 23440 50124 23446 50136
rect 25225 50133 25237 50136
rect 25271 50133 25283 50167
rect 25225 50127 25283 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 19794 49852 19800 49904
rect 19852 49892 19858 49904
rect 19852 49864 24808 49892
rect 19852 49852 19858 49864
rect 23385 49827 23443 49833
rect 23385 49793 23397 49827
rect 23431 49824 23443 49827
rect 24210 49824 24216 49836
rect 23431 49796 24216 49824
rect 23431 49793 23443 49796
rect 23385 49787 23443 49793
rect 24210 49784 24216 49796
rect 24268 49784 24274 49836
rect 24780 49833 24808 49864
rect 24765 49827 24823 49833
rect 24765 49793 24777 49827
rect 24811 49793 24823 49827
rect 24765 49787 24823 49793
rect 24029 49759 24087 49765
rect 24029 49725 24041 49759
rect 24075 49756 24087 49759
rect 24489 49759 24547 49765
rect 24489 49756 24501 49759
rect 24075 49728 24501 49756
rect 24075 49725 24087 49728
rect 24029 49719 24087 49725
rect 24489 49725 24501 49728
rect 24535 49725 24547 49759
rect 24489 49719 24547 49725
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 24210 49376 24216 49428
rect 24268 49416 24274 49428
rect 24762 49416 24768 49428
rect 24268 49388 24768 49416
rect 24268 49376 24274 49388
rect 24762 49376 24768 49388
rect 24820 49376 24826 49428
rect 10686 49308 10692 49360
rect 10744 49308 10750 49360
rect 11698 49308 11704 49360
rect 11756 49308 11762 49360
rect 24673 49215 24731 49221
rect 24673 49181 24685 49215
rect 24719 49212 24731 49215
rect 24854 49212 24860 49224
rect 24719 49184 24860 49212
rect 24719 49181 24731 49184
rect 24673 49175 24731 49181
rect 24854 49172 24860 49184
rect 24912 49172 24918 49224
rect 10226 49104 10232 49156
rect 10284 49144 10290 49156
rect 10505 49147 10563 49153
rect 10505 49144 10517 49147
rect 10284 49116 10517 49144
rect 10284 49104 10290 49116
rect 10505 49113 10517 49116
rect 10551 49113 10563 49147
rect 10505 49107 10563 49113
rect 10870 49104 10876 49156
rect 10928 49144 10934 49156
rect 11517 49147 11575 49153
rect 11517 49144 11529 49147
rect 10928 49116 11529 49144
rect 10928 49104 10934 49116
rect 11517 49113 11529 49116
rect 11563 49113 11575 49147
rect 11517 49107 11575 49113
rect 25130 49036 25136 49088
rect 25188 49076 25194 49088
rect 25317 49079 25375 49085
rect 25317 49076 25329 49079
rect 25188 49048 25329 49076
rect 25188 49036 25194 49048
rect 25317 49045 25329 49048
rect 25363 49045 25375 49079
rect 25317 49039 25375 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 9122 48872 9128 48884
rect 6656 48844 9128 48872
rect 6656 48745 6684 48844
rect 9122 48832 9128 48844
rect 9180 48832 9186 48884
rect 24765 48875 24823 48881
rect 24765 48841 24777 48875
rect 24811 48872 24823 48875
rect 24854 48872 24860 48884
rect 24811 48844 24860 48872
rect 24811 48841 24823 48844
rect 24765 48835 24823 48841
rect 24854 48832 24860 48844
rect 24912 48832 24918 48884
rect 25130 48764 25136 48816
rect 25188 48764 25194 48816
rect 6641 48739 6699 48745
rect 6641 48705 6653 48739
rect 6687 48705 6699 48739
rect 8050 48708 8800 48736
rect 6641 48699 6699 48705
rect 6917 48671 6975 48677
rect 6917 48637 6929 48671
rect 6963 48668 6975 48671
rect 8294 48668 8300 48680
rect 6963 48640 8300 48668
rect 6963 48637 6975 48640
rect 6917 48631 6975 48637
rect 8294 48628 8300 48640
rect 8352 48628 8358 48680
rect 8386 48628 8392 48680
rect 8444 48628 8450 48680
rect 8772 48609 8800 48708
rect 8757 48603 8815 48609
rect 8757 48569 8769 48603
rect 8803 48600 8815 48603
rect 9950 48600 9956 48612
rect 8803 48572 9956 48600
rect 8803 48569 8815 48572
rect 8757 48563 8815 48569
rect 9950 48560 9956 48572
rect 10008 48560 10014 48612
rect 25317 48603 25375 48609
rect 25317 48569 25329 48603
rect 25363 48600 25375 48603
rect 26142 48600 26148 48612
rect 25363 48572 26148 48600
rect 25363 48569 25375 48572
rect 25317 48563 25375 48569
rect 26142 48560 26148 48572
rect 26200 48560 26206 48612
rect 8941 48535 8999 48541
rect 8941 48501 8953 48535
rect 8987 48532 8999 48535
rect 9122 48532 9128 48544
rect 8987 48504 9128 48532
rect 8987 48501 8999 48504
rect 8941 48495 8999 48501
rect 9122 48492 9128 48504
rect 9180 48492 9186 48544
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 7742 48084 7748 48136
rect 7800 48124 7806 48136
rect 10356 48127 10414 48133
rect 10356 48124 10368 48127
rect 7800 48096 10368 48124
rect 7800 48084 7806 48096
rect 10356 48093 10368 48096
rect 10402 48093 10414 48127
rect 10356 48087 10414 48093
rect 23382 48084 23388 48136
rect 23440 48084 23446 48136
rect 24673 48127 24731 48133
rect 24673 48093 24685 48127
rect 24719 48124 24731 48127
rect 24854 48124 24860 48136
rect 24719 48096 24860 48124
rect 24719 48093 24731 48096
rect 24673 48087 24731 48093
rect 24854 48084 24860 48096
rect 24912 48084 24918 48136
rect 10459 47991 10517 47997
rect 10459 47957 10471 47991
rect 10505 47988 10517 47991
rect 13722 47988 13728 48000
rect 10505 47960 13728 47988
rect 10505 47957 10517 47960
rect 10459 47951 10517 47957
rect 13722 47948 13728 47960
rect 13780 47948 13786 48000
rect 24026 47948 24032 48000
rect 24084 47948 24090 48000
rect 25130 47948 25136 48000
rect 25188 47988 25194 48000
rect 25317 47991 25375 47997
rect 25317 47988 25329 47991
rect 25188 47960 25329 47988
rect 25188 47948 25194 47960
rect 25317 47957 25329 47960
rect 25363 47957 25375 47991
rect 25317 47951 25375 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9214 47744 9220 47796
rect 9272 47784 9278 47796
rect 9490 47784 9496 47796
rect 9272 47756 9496 47784
rect 9272 47744 9278 47756
rect 9490 47744 9496 47756
rect 9548 47784 9554 47796
rect 9861 47787 9919 47793
rect 9861 47784 9873 47787
rect 9548 47756 9873 47784
rect 9548 47744 9554 47756
rect 9861 47753 9873 47756
rect 9907 47753 9919 47787
rect 9861 47747 9919 47753
rect 24765 47787 24823 47793
rect 24765 47753 24777 47787
rect 24811 47784 24823 47787
rect 24854 47784 24860 47796
rect 24811 47756 24860 47784
rect 24811 47753 24823 47756
rect 24765 47747 24823 47753
rect 24854 47744 24860 47756
rect 24912 47744 24918 47796
rect 8570 47676 8576 47728
rect 8628 47716 8634 47728
rect 10137 47719 10195 47725
rect 10137 47716 10149 47719
rect 8628 47688 10149 47716
rect 8628 47676 8634 47688
rect 9416 47657 9444 47688
rect 10137 47685 10149 47688
rect 10183 47716 10195 47719
rect 10962 47716 10968 47728
rect 10183 47688 10968 47716
rect 10183 47685 10195 47688
rect 10137 47679 10195 47685
rect 10962 47676 10968 47688
rect 11020 47676 11026 47728
rect 25130 47676 25136 47728
rect 25188 47676 25194 47728
rect 9401 47651 9459 47657
rect 9401 47617 9413 47651
rect 9447 47648 9459 47651
rect 9447 47620 9481 47648
rect 9447 47617 9459 47620
rect 9401 47611 9459 47617
rect 16206 47540 16212 47592
rect 16264 47580 16270 47592
rect 25222 47580 25228 47592
rect 16264 47552 25228 47580
rect 16264 47540 16270 47552
rect 25222 47540 25228 47552
rect 25280 47540 25286 47592
rect 25317 47515 25375 47521
rect 25317 47481 25329 47515
rect 25363 47512 25375 47515
rect 25682 47512 25688 47524
rect 25363 47484 25688 47512
rect 25363 47481 25375 47484
rect 25317 47475 25375 47481
rect 25682 47472 25688 47484
rect 25740 47472 25746 47524
rect 8294 47404 8300 47456
rect 8352 47444 8358 47456
rect 9490 47444 9496 47456
rect 8352 47416 9496 47444
rect 8352 47404 8358 47416
rect 9490 47404 9496 47416
rect 9548 47404 9554 47456
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 25133 47175 25191 47181
rect 25133 47141 25145 47175
rect 25179 47172 25191 47175
rect 26510 47172 26516 47184
rect 25179 47144 26516 47172
rect 25179 47141 25191 47144
rect 25133 47135 25191 47141
rect 26510 47132 26516 47144
rect 26568 47132 26574 47184
rect 9214 46996 9220 47048
rect 9272 47036 9278 47048
rect 11644 47039 11702 47045
rect 11644 47036 11656 47039
rect 9272 47008 11656 47036
rect 9272 46996 9278 47008
rect 11644 47005 11656 47008
rect 11690 47005 11702 47039
rect 11644 46999 11702 47005
rect 24857 47039 24915 47045
rect 24857 47005 24869 47039
rect 24903 47036 24915 47039
rect 25314 47036 25320 47048
rect 24903 47008 25320 47036
rect 24903 47005 24915 47008
rect 24857 46999 24915 47005
rect 25314 46996 25320 47008
rect 25372 46996 25378 47048
rect 11747 46971 11805 46977
rect 11747 46937 11759 46971
rect 11793 46968 11805 46971
rect 13630 46968 13636 46980
rect 11793 46940 13636 46968
rect 11793 46937 11805 46940
rect 11747 46931 11805 46937
rect 13630 46928 13636 46940
rect 13688 46928 13694 46980
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 10778 46656 10784 46708
rect 10836 46656 10842 46708
rect 10962 46656 10968 46708
rect 11020 46696 11026 46708
rect 11057 46699 11115 46705
rect 11057 46696 11069 46699
rect 11020 46668 11069 46696
rect 11020 46656 11026 46668
rect 11057 46665 11069 46668
rect 11103 46665 11115 46699
rect 11057 46659 11115 46665
rect 13630 46656 13636 46708
rect 13688 46696 13694 46708
rect 13688 46668 14872 46696
rect 13688 46656 13694 46668
rect 10980 46628 11008 46656
rect 10336 46600 11008 46628
rect 10336 46569 10364 46600
rect 10321 46563 10379 46569
rect 10321 46529 10333 46563
rect 10367 46529 10379 46563
rect 10321 46523 10379 46529
rect 10704 46424 10732 46600
rect 14734 46588 14740 46640
rect 14792 46588 14798 46640
rect 14844 46637 14872 46668
rect 14829 46631 14887 46637
rect 14829 46597 14841 46631
rect 14875 46597 14887 46631
rect 14829 46591 14887 46597
rect 10778 46520 10784 46572
rect 10836 46560 10842 46572
rect 12564 46563 12622 46569
rect 12564 46560 12576 46563
rect 10836 46532 12576 46560
rect 10836 46520 10842 46532
rect 12564 46529 12576 46532
rect 12610 46529 12622 46563
rect 12564 46523 12622 46529
rect 24857 46563 24915 46569
rect 24857 46529 24869 46563
rect 24903 46560 24915 46563
rect 25314 46560 25320 46572
rect 24903 46532 25320 46560
rect 24903 46529 24915 46532
rect 24857 46523 24915 46529
rect 25314 46520 25320 46532
rect 25372 46520 25378 46572
rect 15746 46452 15752 46504
rect 15804 46452 15810 46504
rect 10778 46424 10784 46436
rect 10704 46396 10784 46424
rect 10778 46384 10784 46396
rect 10836 46384 10842 46436
rect 10410 46316 10416 46368
rect 10468 46316 10474 46368
rect 12667 46359 12725 46365
rect 12667 46325 12679 46359
rect 12713 46356 12725 46359
rect 15470 46356 15476 46368
rect 12713 46328 15476 46356
rect 12713 46325 12725 46328
rect 12667 46319 12725 46325
rect 15470 46316 15476 46328
rect 15528 46316 15534 46368
rect 21174 46316 21180 46368
rect 21232 46356 21238 46368
rect 25133 46359 25191 46365
rect 25133 46356 25145 46359
rect 21232 46328 25145 46356
rect 21232 46316 21238 46328
rect 25133 46325 25145 46328
rect 25179 46325 25191 46359
rect 25133 46319 25191 46325
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 8478 46112 8484 46164
rect 8536 46112 8542 46164
rect 7742 45976 7748 46028
rect 7800 46016 7806 46028
rect 8113 46019 8171 46025
rect 8113 46016 8125 46019
rect 7800 45988 8125 46016
rect 7800 45976 7806 45988
rect 8113 45985 8125 45988
rect 8159 45985 8171 46019
rect 8113 45979 8171 45985
rect 15654 45976 15660 46028
rect 15712 45976 15718 46028
rect 16482 45976 16488 46028
rect 16540 45976 16546 46028
rect 7834 45908 7840 45960
rect 7892 45948 7898 45960
rect 7929 45951 7987 45957
rect 7929 45948 7941 45951
rect 7892 45920 7941 45948
rect 7892 45908 7898 45920
rect 7929 45917 7941 45920
rect 7975 45917 7987 45951
rect 7929 45911 7987 45917
rect 12802 45908 12808 45960
rect 12860 45948 12866 45960
rect 13300 45951 13358 45957
rect 13300 45948 13312 45951
rect 12860 45920 13312 45948
rect 12860 45908 12866 45920
rect 13300 45917 13312 45920
rect 13346 45917 13358 45951
rect 13300 45911 13358 45917
rect 24857 45951 24915 45957
rect 24857 45917 24869 45951
rect 24903 45948 24915 45951
rect 25314 45948 25320 45960
rect 24903 45920 25320 45948
rect 24903 45917 24915 45920
rect 24857 45911 24915 45917
rect 25314 45908 25320 45920
rect 25372 45908 25378 45960
rect 15470 45840 15476 45892
rect 15528 45880 15534 45892
rect 15749 45883 15807 45889
rect 15749 45880 15761 45883
rect 15528 45852 15761 45880
rect 15528 45840 15534 45852
rect 15749 45849 15761 45852
rect 15795 45849 15807 45883
rect 15749 45843 15807 45849
rect 13403 45815 13461 45821
rect 13403 45781 13415 45815
rect 13449 45812 13461 45815
rect 14918 45812 14924 45824
rect 13449 45784 14924 45812
rect 13449 45781 13461 45784
rect 13403 45775 13461 45781
rect 14918 45772 14924 45784
rect 14976 45772 14982 45824
rect 25038 45772 25044 45824
rect 25096 45812 25102 45824
rect 25133 45815 25191 45821
rect 25133 45812 25145 45815
rect 25096 45784 25145 45812
rect 25096 45772 25102 45784
rect 25133 45781 25145 45784
rect 25179 45781 25191 45815
rect 25133 45775 25191 45781
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 10502 45500 10508 45552
rect 10560 45540 10566 45552
rect 12802 45540 12808 45552
rect 10560 45512 12808 45540
rect 10560 45500 10566 45512
rect 12802 45500 12808 45512
rect 12860 45500 12866 45552
rect 13538 45500 13544 45552
rect 13596 45500 13602 45552
rect 13633 45543 13691 45549
rect 13633 45509 13645 45543
rect 13679 45540 13691 45543
rect 13722 45540 13728 45552
rect 13679 45512 13728 45540
rect 13679 45509 13691 45512
rect 13633 45503 13691 45509
rect 13722 45500 13728 45512
rect 13780 45500 13786 45552
rect 24857 45475 24915 45481
rect 24857 45441 24869 45475
rect 24903 45472 24915 45475
rect 25317 45475 25375 45481
rect 25317 45472 25329 45475
rect 24903 45444 25329 45472
rect 24903 45441 24915 45444
rect 24857 45435 24915 45441
rect 25317 45441 25329 45444
rect 25363 45472 25375 45475
rect 25406 45472 25412 45484
rect 25363 45444 25412 45472
rect 25363 45441 25375 45444
rect 25317 45435 25375 45441
rect 25406 45432 25412 45444
rect 25464 45432 25470 45484
rect 14550 45364 14556 45416
rect 14608 45364 14614 45416
rect 25133 45271 25191 45277
rect 25133 45237 25145 45271
rect 25179 45268 25191 45271
rect 25222 45268 25228 45280
rect 25179 45240 25228 45268
rect 25179 45237 25191 45240
rect 25133 45231 25191 45237
rect 25222 45228 25228 45240
rect 25280 45228 25286 45280
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 9490 45024 9496 45076
rect 9548 45064 9554 45076
rect 10873 45067 10931 45073
rect 10873 45064 10885 45067
rect 9548 45036 10885 45064
rect 9548 45024 9554 45036
rect 10873 45033 10885 45036
rect 10919 45033 10931 45067
rect 10873 45027 10931 45033
rect 16022 44956 16028 45008
rect 16080 44996 16086 45008
rect 24946 44996 24952 45008
rect 16080 44968 24952 44996
rect 16080 44956 16086 44968
rect 24946 44956 24952 44968
rect 25004 44956 25010 45008
rect 9950 44888 9956 44940
rect 10008 44928 10014 44940
rect 16485 44931 16543 44937
rect 10008 44900 10640 44928
rect 10008 44888 10014 44900
rect 9122 44820 9128 44872
rect 9180 44820 9186 44872
rect 9401 44795 9459 44801
rect 9401 44761 9413 44795
rect 9447 44792 9459 44795
rect 9674 44792 9680 44804
rect 9447 44764 9680 44792
rect 9447 44761 9459 44764
rect 9401 44755 9459 44761
rect 9674 44752 9680 44764
rect 9732 44752 9738 44804
rect 10612 44792 10640 44900
rect 16485 44897 16497 44931
rect 16531 44928 16543 44931
rect 17678 44928 17684 44940
rect 16531 44900 17684 44928
rect 16531 44897 16543 44900
rect 16485 44891 16543 44897
rect 17678 44888 17684 44900
rect 17736 44888 17742 44940
rect 11241 44795 11299 44801
rect 11241 44792 11253 44795
rect 10612 44778 11253 44792
rect 10626 44764 11253 44778
rect 11241 44761 11253 44764
rect 11287 44792 11299 44795
rect 11514 44792 11520 44804
rect 11287 44764 11520 44792
rect 11287 44761 11299 44764
rect 11241 44755 11299 44761
rect 11514 44752 11520 44764
rect 11572 44752 11578 44804
rect 14918 44752 14924 44804
rect 14976 44792 14982 44804
rect 16554 44795 16612 44801
rect 16554 44792 16566 44795
rect 14976 44764 16566 44792
rect 14976 44752 14982 44764
rect 16554 44761 16566 44764
rect 16600 44761 16612 44795
rect 16554 44755 16612 44761
rect 17494 44752 17500 44804
rect 17552 44752 17558 44804
rect 25133 44795 25191 44801
rect 25133 44761 25145 44795
rect 25179 44792 25191 44795
rect 25314 44792 25320 44804
rect 25179 44764 25320 44792
rect 25179 44761 25191 44764
rect 25133 44755 25191 44761
rect 25314 44752 25320 44764
rect 25372 44752 25378 44804
rect 9692 44724 9720 44752
rect 10410 44724 10416 44736
rect 9692 44696 10416 44724
rect 10410 44684 10416 44696
rect 10468 44684 10474 44736
rect 11425 44727 11483 44733
rect 11425 44693 11437 44727
rect 11471 44724 11483 44727
rect 11698 44724 11704 44736
rect 11471 44696 11704 44724
rect 11471 44693 11483 44696
rect 11425 44687 11483 44693
rect 11698 44684 11704 44696
rect 11756 44684 11762 44736
rect 25225 44727 25283 44733
rect 25225 44693 25237 44727
rect 25271 44724 25283 44727
rect 25498 44724 25504 44736
rect 25271 44696 25504 44724
rect 25271 44693 25283 44696
rect 25225 44687 25283 44693
rect 25498 44684 25504 44696
rect 25556 44684 25562 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 9582 44480 9588 44532
rect 9640 44480 9646 44532
rect 13814 44480 13820 44532
rect 13872 44520 13878 44532
rect 17494 44520 17500 44532
rect 13872 44492 17500 44520
rect 13872 44480 13878 44492
rect 17494 44480 17500 44492
rect 17552 44480 17558 44532
rect 25314 44480 25320 44532
rect 25372 44480 25378 44532
rect 9125 44387 9183 44393
rect 9125 44353 9137 44387
rect 9171 44384 9183 44387
rect 9214 44384 9220 44396
rect 9171 44356 9220 44384
rect 9171 44353 9183 44356
rect 9125 44347 9183 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 10597 44387 10655 44393
rect 10597 44353 10609 44387
rect 10643 44384 10655 44387
rect 10778 44384 10784 44396
rect 10643 44356 10784 44384
rect 10643 44353 10655 44356
rect 10597 44347 10655 44353
rect 10778 44344 10784 44356
rect 10836 44384 10842 44396
rect 11517 44387 11575 44393
rect 11517 44384 11529 44387
rect 10836 44356 11529 44384
rect 10836 44344 10842 44356
rect 11517 44353 11529 44356
rect 11563 44353 11575 44387
rect 11517 44347 11575 44353
rect 24397 44387 24455 44393
rect 24397 44353 24409 44387
rect 24443 44384 24455 44387
rect 24670 44384 24676 44396
rect 24443 44356 24676 44384
rect 24443 44353 24455 44356
rect 24397 44347 24455 44353
rect 24670 44344 24676 44356
rect 24728 44344 24734 44396
rect 8941 44319 8999 44325
rect 8941 44285 8953 44319
rect 8987 44316 8999 44319
rect 9306 44316 9312 44328
rect 8987 44288 9312 44316
rect 8987 44285 8999 44288
rect 8941 44279 8999 44285
rect 9306 44276 9312 44288
rect 9364 44276 9370 44328
rect 10502 44208 10508 44260
rect 10560 44248 10566 44260
rect 10560 44220 11008 44248
rect 10560 44208 10566 44220
rect 10980 44192 11008 44220
rect 10686 44140 10692 44192
rect 10744 44140 10750 44192
rect 10962 44140 10968 44192
rect 11020 44180 11026 44192
rect 11057 44183 11115 44189
rect 11057 44180 11069 44183
rect 11020 44152 11069 44180
rect 11020 44140 11026 44152
rect 11057 44149 11069 44152
rect 11103 44149 11115 44183
rect 11057 44143 11115 44149
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 20625 43843 20683 43849
rect 20625 43809 20637 43843
rect 20671 43840 20683 43843
rect 24026 43840 24032 43852
rect 20671 43812 24032 43840
rect 20671 43809 20683 43812
rect 20625 43803 20683 43809
rect 24026 43800 24032 43812
rect 24084 43800 24090 43852
rect 19518 43732 19524 43784
rect 19576 43772 19582 43784
rect 20349 43775 20407 43781
rect 20349 43772 20361 43775
rect 19576 43744 20361 43772
rect 19576 43732 19582 43744
rect 20349 43741 20361 43744
rect 20395 43741 20407 43775
rect 20349 43735 20407 43741
rect 20073 43707 20131 43713
rect 20073 43673 20085 43707
rect 20119 43704 20131 43707
rect 21082 43704 21088 43716
rect 20119 43676 21088 43704
rect 20119 43673 20131 43676
rect 20073 43667 20131 43673
rect 21082 43664 21088 43676
rect 21140 43664 21146 43716
rect 25133 43707 25191 43713
rect 25133 43673 25145 43707
rect 25179 43704 25191 43707
rect 25314 43704 25320 43716
rect 25179 43676 25320 43704
rect 25179 43673 25191 43676
rect 25133 43667 25191 43673
rect 25314 43664 25320 43676
rect 25372 43664 25378 43716
rect 21358 43596 21364 43648
rect 21416 43636 21422 43648
rect 22097 43639 22155 43645
rect 22097 43636 22109 43639
rect 21416 43608 22109 43636
rect 21416 43596 21422 43608
rect 22097 43605 22109 43608
rect 22143 43605 22155 43639
rect 22097 43599 22155 43605
rect 24854 43596 24860 43648
rect 24912 43636 24918 43648
rect 25225 43639 25283 43645
rect 25225 43636 25237 43639
rect 24912 43608 25237 43636
rect 24912 43596 24918 43608
rect 25225 43605 25237 43608
rect 25271 43605 25283 43639
rect 25225 43599 25283 43605
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 25314 43392 25320 43444
rect 25372 43392 25378 43444
rect 24397 43299 24455 43305
rect 24397 43265 24409 43299
rect 24443 43296 24455 43299
rect 24673 43299 24731 43305
rect 24673 43296 24685 43299
rect 24443 43268 24685 43296
rect 24443 43265 24455 43268
rect 24397 43259 24455 43265
rect 24673 43265 24685 43268
rect 24719 43296 24731 43299
rect 24946 43296 24952 43308
rect 24719 43268 24952 43296
rect 24719 43265 24731 43268
rect 24673 43259 24731 43265
rect 24946 43256 24952 43268
rect 25004 43256 25010 43308
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 24854 42780 24860 42832
rect 24912 42780 24918 42832
rect 10226 42712 10232 42764
rect 10284 42712 10290 42764
rect 21266 42712 21272 42764
rect 21324 42752 21330 42764
rect 24872 42752 24900 42780
rect 21324 42724 24900 42752
rect 21324 42712 21330 42724
rect 8938 42644 8944 42696
rect 8996 42684 9002 42696
rect 9585 42687 9643 42693
rect 9585 42684 9597 42687
rect 8996 42656 9597 42684
rect 8996 42644 9002 42656
rect 9585 42653 9597 42656
rect 9631 42653 9643 42687
rect 9585 42647 9643 42653
rect 9769 42687 9827 42693
rect 9769 42653 9781 42687
rect 9815 42684 9827 42687
rect 10594 42684 10600 42696
rect 9815 42656 10600 42684
rect 9815 42653 9827 42656
rect 9769 42647 9827 42653
rect 10594 42644 10600 42656
rect 10652 42644 10658 42696
rect 24673 42687 24731 42693
rect 24673 42653 24685 42687
rect 24719 42684 24731 42687
rect 24854 42684 24860 42696
rect 24719 42656 24860 42684
rect 24719 42653 24731 42656
rect 24673 42647 24731 42653
rect 24854 42644 24860 42656
rect 24912 42644 24918 42696
rect 25130 42508 25136 42560
rect 25188 42548 25194 42560
rect 25317 42551 25375 42557
rect 25317 42548 25329 42551
rect 25188 42520 25329 42548
rect 25188 42508 25194 42520
rect 25317 42517 25329 42520
rect 25363 42517 25375 42551
rect 25317 42511 25375 42517
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 9674 42304 9680 42356
rect 9732 42344 9738 42356
rect 11149 42347 11207 42353
rect 11149 42344 11161 42347
rect 9732 42316 11161 42344
rect 9732 42304 9738 42316
rect 11149 42313 11161 42316
rect 11195 42313 11207 42347
rect 11149 42307 11207 42313
rect 24765 42347 24823 42353
rect 24765 42313 24777 42347
rect 24811 42344 24823 42347
rect 24854 42344 24860 42356
rect 24811 42316 24860 42344
rect 24811 42313 24823 42316
rect 24765 42307 24823 42313
rect 24854 42304 24860 42316
rect 24912 42304 24918 42356
rect 11514 42276 11520 42288
rect 10902 42248 11520 42276
rect 11514 42236 11520 42248
rect 11572 42236 11578 42288
rect 25130 42236 25136 42288
rect 25188 42236 25194 42288
rect 9122 42100 9128 42152
rect 9180 42140 9186 42152
rect 9401 42143 9459 42149
rect 9401 42140 9413 42143
rect 9180 42112 9413 42140
rect 9180 42100 9186 42112
rect 9401 42109 9413 42112
rect 9447 42109 9459 42143
rect 9401 42103 9459 42109
rect 9416 42004 9444 42103
rect 9674 42100 9680 42152
rect 9732 42140 9738 42152
rect 10686 42140 10692 42152
rect 9732 42112 10692 42140
rect 9732 42100 9738 42112
rect 10686 42100 10692 42112
rect 10744 42100 10750 42152
rect 10704 42044 11744 42072
rect 10704 42004 10732 42044
rect 11716 42016 11744 42044
rect 15838 42032 15844 42084
rect 15896 42072 15902 42084
rect 24486 42072 24492 42084
rect 15896 42044 24492 42072
rect 15896 42032 15902 42044
rect 24486 42032 24492 42044
rect 24544 42032 24550 42084
rect 9416 41976 10732 42004
rect 11514 41964 11520 42016
rect 11572 41964 11578 42016
rect 11698 41964 11704 42016
rect 11756 41964 11762 42016
rect 21726 41964 21732 42016
rect 21784 42004 21790 42016
rect 25225 42007 25283 42013
rect 25225 42004 25237 42007
rect 21784 41976 25237 42004
rect 21784 41964 21790 41976
rect 25225 41973 25237 41976
rect 25271 41973 25283 42007
rect 25225 41967 25283 41973
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 10870 41760 10876 41812
rect 10928 41760 10934 41812
rect 10413 41667 10471 41673
rect 10413 41633 10425 41667
rect 10459 41664 10471 41667
rect 10962 41664 10968 41676
rect 10459 41636 10968 41664
rect 10459 41633 10471 41636
rect 10413 41627 10471 41633
rect 10962 41624 10968 41636
rect 11020 41624 11026 41676
rect 10226 41556 10232 41608
rect 10284 41556 10290 41608
rect 16850 41556 16856 41608
rect 16908 41596 16914 41608
rect 21450 41596 21456 41608
rect 16908 41568 21456 41596
rect 16908 41556 16914 41568
rect 21450 41556 21456 41568
rect 21508 41556 21514 41608
rect 24673 41599 24731 41605
rect 24673 41565 24685 41599
rect 24719 41596 24731 41599
rect 24854 41596 24860 41608
rect 24719 41568 24860 41596
rect 24719 41565 24731 41568
rect 24673 41559 24731 41565
rect 24854 41556 24860 41568
rect 24912 41556 24918 41608
rect 25314 41420 25320 41472
rect 25372 41420 25378 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 24762 41216 24768 41268
rect 24820 41216 24826 41268
rect 25133 41191 25191 41197
rect 25133 41157 25145 41191
rect 25179 41188 25191 41191
rect 25314 41188 25320 41200
rect 25179 41160 25320 41188
rect 25179 41157 25191 41160
rect 25133 41151 25191 41157
rect 25314 41148 25320 41160
rect 25372 41148 25378 41200
rect 24854 40876 24860 40928
rect 24912 40916 24918 40928
rect 25225 40919 25283 40925
rect 25225 40916 25237 40919
rect 24912 40888 25237 40916
rect 24912 40876 24918 40888
rect 25225 40885 25237 40888
rect 25271 40885 25283 40919
rect 25225 40879 25283 40885
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 24857 40511 24915 40517
rect 24857 40477 24869 40511
rect 24903 40508 24915 40511
rect 25314 40508 25320 40520
rect 24903 40480 25320 40508
rect 24903 40477 24915 40480
rect 24857 40471 24915 40477
rect 25314 40468 25320 40480
rect 25372 40468 25378 40520
rect 25133 40375 25191 40381
rect 25133 40341 25145 40375
rect 25179 40372 25191 40375
rect 25406 40372 25412 40384
rect 25179 40344 25412 40372
rect 25179 40341 25191 40344
rect 25133 40335 25191 40341
rect 25406 40332 25412 40344
rect 25464 40332 25470 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 23290 40128 23296 40180
rect 23348 40168 23354 40180
rect 25133 40171 25191 40177
rect 25133 40168 25145 40171
rect 23348 40140 25145 40168
rect 23348 40128 23354 40140
rect 25133 40137 25145 40140
rect 25179 40137 25191 40171
rect 25133 40131 25191 40137
rect 24857 40035 24915 40041
rect 24857 40001 24869 40035
rect 24903 40032 24915 40035
rect 25314 40032 25320 40044
rect 24903 40004 25320 40032
rect 24903 40001 24915 40004
rect 24857 39995 24915 40001
rect 25314 39992 25320 40004
rect 25372 39992 25378 40044
rect 17034 39924 17040 39976
rect 17092 39964 17098 39976
rect 23658 39964 23664 39976
rect 17092 39936 23664 39964
rect 17092 39924 17098 39936
rect 23658 39924 23664 39936
rect 23716 39924 23722 39976
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 10686 39584 10692 39636
rect 10744 39624 10750 39636
rect 13814 39624 13820 39636
rect 10744 39596 13820 39624
rect 10744 39584 10750 39596
rect 13814 39584 13820 39596
rect 13872 39584 13878 39636
rect 24857 39423 24915 39429
rect 24857 39389 24869 39423
rect 24903 39420 24915 39423
rect 25314 39420 25320 39432
rect 24903 39392 25320 39420
rect 24903 39389 24915 39392
rect 24857 39383 24915 39389
rect 25314 39380 25320 39392
rect 25372 39380 25378 39432
rect 24118 39244 24124 39296
rect 24176 39284 24182 39296
rect 25133 39287 25191 39293
rect 25133 39284 25145 39287
rect 24176 39256 25145 39284
rect 24176 39244 24182 39256
rect 25133 39253 25145 39256
rect 25179 39253 25191 39287
rect 25133 39247 25191 39253
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 25317 38947 25375 38953
rect 25317 38944 25329 38947
rect 24872 38916 25329 38944
rect 24762 38700 24768 38752
rect 24820 38740 24826 38752
rect 24872 38749 24900 38916
rect 25317 38913 25329 38916
rect 25363 38913 25375 38947
rect 25317 38907 25375 38913
rect 24857 38743 24915 38749
rect 24857 38740 24869 38743
rect 24820 38712 24869 38740
rect 24820 38700 24826 38712
rect 24857 38709 24869 38712
rect 24903 38709 24915 38743
rect 24857 38703 24915 38709
rect 25038 38700 25044 38752
rect 25096 38740 25102 38752
rect 25133 38743 25191 38749
rect 25133 38740 25145 38743
rect 25096 38712 25145 38740
rect 25096 38700 25102 38712
rect 25133 38709 25145 38712
rect 25179 38709 25191 38743
rect 25133 38703 25191 38709
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 16942 38496 16948 38548
rect 17000 38536 17006 38548
rect 19978 38536 19984 38548
rect 17000 38508 19984 38536
rect 17000 38496 17006 38508
rect 19978 38496 19984 38508
rect 20036 38496 20042 38548
rect 25133 38267 25191 38273
rect 25133 38233 25145 38267
rect 25179 38264 25191 38267
rect 25314 38264 25320 38276
rect 25179 38236 25320 38264
rect 25179 38233 25191 38236
rect 25133 38227 25191 38233
rect 25314 38224 25320 38236
rect 25372 38224 25378 38276
rect 25225 38199 25283 38205
rect 25225 38165 25237 38199
rect 25271 38196 25283 38199
rect 25866 38196 25872 38208
rect 25271 38168 25872 38196
rect 25271 38165 25283 38168
rect 25225 38159 25283 38165
rect 25866 38156 25872 38168
rect 25924 38156 25930 38208
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 7834 37952 7840 38004
rect 7892 37992 7898 38004
rect 8665 37995 8723 38001
rect 8665 37992 8677 37995
rect 7892 37964 8677 37992
rect 7892 37952 7898 37964
rect 8665 37961 8677 37964
rect 8711 37961 8723 37995
rect 8665 37955 8723 37961
rect 25314 37952 25320 38004
rect 25372 37952 25378 38004
rect 9030 37884 9036 37936
rect 9088 37924 9094 37936
rect 15746 37924 15752 37936
rect 9088 37896 15752 37924
rect 9088 37884 9094 37896
rect 15746 37884 15752 37896
rect 15804 37884 15810 37936
rect 8846 37816 8852 37868
rect 8904 37816 8910 37868
rect 24397 37859 24455 37865
rect 24397 37825 24409 37859
rect 24443 37856 24455 37859
rect 24673 37859 24731 37865
rect 24673 37856 24685 37859
rect 24443 37828 24685 37856
rect 24443 37825 24455 37828
rect 24397 37819 24455 37825
rect 24673 37825 24685 37828
rect 24719 37856 24731 37859
rect 24854 37856 24860 37868
rect 24719 37828 24860 37856
rect 24719 37825 24731 37828
rect 24673 37819 24731 37825
rect 24854 37816 24860 37828
rect 24912 37816 24918 37868
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 25317 37315 25375 37321
rect 25317 37281 25329 37315
rect 25363 37312 25375 37315
rect 25590 37312 25596 37324
rect 25363 37284 25596 37312
rect 25363 37281 25375 37284
rect 25317 37275 25375 37281
rect 25590 37272 25596 37284
rect 25648 37272 25654 37324
rect 25133 37179 25191 37185
rect 25133 37145 25145 37179
rect 25179 37176 25191 37179
rect 25314 37176 25320 37188
rect 25179 37148 25320 37176
rect 25179 37145 25191 37148
rect 25133 37139 25191 37145
rect 25314 37136 25320 37148
rect 25372 37136 25378 37188
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 25314 36864 25320 36916
rect 25372 36864 25378 36916
rect 24397 36771 24455 36777
rect 24397 36737 24409 36771
rect 24443 36768 24455 36771
rect 24673 36771 24731 36777
rect 24673 36768 24685 36771
rect 24443 36740 24685 36768
rect 24443 36737 24455 36740
rect 24397 36731 24455 36737
rect 24673 36737 24685 36740
rect 24719 36768 24731 36771
rect 24946 36768 24952 36780
rect 24719 36740 24952 36768
rect 24719 36737 24731 36740
rect 24673 36731 24731 36737
rect 24946 36728 24952 36740
rect 25004 36728 25010 36780
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 24213 36159 24271 36165
rect 24213 36125 24225 36159
rect 24259 36156 24271 36159
rect 24673 36159 24731 36165
rect 24673 36156 24685 36159
rect 24259 36128 24685 36156
rect 24259 36125 24271 36128
rect 24213 36119 24271 36125
rect 24673 36125 24685 36128
rect 24719 36156 24731 36159
rect 24762 36156 24768 36168
rect 24719 36128 24768 36156
rect 24719 36125 24731 36128
rect 24673 36119 24731 36125
rect 24762 36116 24768 36128
rect 24820 36116 24826 36168
rect 24670 35980 24676 36032
rect 24728 36020 24734 36032
rect 25317 36023 25375 36029
rect 25317 36020 25329 36023
rect 24728 35992 25329 36020
rect 24728 35980 24734 35992
rect 25317 35989 25329 35992
rect 25363 35989 25375 36023
rect 25317 35983 25375 35989
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 11698 35816 11704 35828
rect 9416 35788 11704 35816
rect 9416 35689 9444 35788
rect 11698 35776 11704 35788
rect 11756 35776 11762 35828
rect 21174 35776 21180 35828
rect 21232 35776 21238 35828
rect 22465 35819 22523 35825
rect 22465 35785 22477 35819
rect 22511 35816 22523 35819
rect 25130 35816 25136 35828
rect 22511 35788 25136 35816
rect 22511 35785 22523 35788
rect 22465 35779 22523 35785
rect 25130 35776 25136 35788
rect 25188 35776 25194 35828
rect 11514 35748 11520 35760
rect 10902 35720 11520 35748
rect 11514 35708 11520 35720
rect 11572 35748 11578 35760
rect 12342 35748 12348 35760
rect 11572 35720 12348 35748
rect 11572 35708 11578 35720
rect 12342 35708 12348 35720
rect 12400 35708 12406 35760
rect 20441 35751 20499 35757
rect 20441 35717 20453 35751
rect 20487 35748 20499 35751
rect 21085 35751 21143 35757
rect 21085 35748 21097 35751
rect 20487 35720 21097 35748
rect 20487 35717 20499 35720
rect 20441 35711 20499 35717
rect 21085 35717 21097 35720
rect 21131 35748 21143 35751
rect 22094 35748 22100 35760
rect 21131 35720 22100 35748
rect 21131 35717 21143 35720
rect 21085 35711 21143 35717
rect 22094 35708 22100 35720
rect 22152 35708 22158 35760
rect 9401 35683 9459 35689
rect 9401 35649 9413 35683
rect 9447 35649 9459 35683
rect 9401 35643 9459 35649
rect 22002 35640 22008 35692
rect 22060 35680 22066 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 22060 35652 22385 35680
rect 22060 35640 22066 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 24670 35640 24676 35692
rect 24728 35640 24734 35692
rect 25314 35640 25320 35692
rect 25372 35640 25378 35692
rect 9677 35615 9735 35621
rect 9677 35581 9689 35615
rect 9723 35612 9735 35615
rect 10042 35612 10048 35624
rect 9723 35584 10048 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 10042 35572 10048 35584
rect 10100 35572 10106 35624
rect 21174 35572 21180 35624
rect 21232 35612 21238 35624
rect 21269 35615 21327 35621
rect 21269 35612 21281 35615
rect 21232 35584 21281 35612
rect 21232 35572 21238 35584
rect 21269 35581 21281 35584
rect 21315 35581 21327 35615
rect 21269 35575 21327 35581
rect 22554 35572 22560 35624
rect 22612 35572 22618 35624
rect 19058 35504 19064 35556
rect 19116 35544 19122 35556
rect 19116 35516 20484 35544
rect 19116 35504 19122 35516
rect 9674 35436 9680 35488
rect 9732 35476 9738 35488
rect 11149 35479 11207 35485
rect 11149 35476 11161 35479
rect 9732 35448 11161 35476
rect 9732 35436 9738 35448
rect 11149 35445 11161 35448
rect 11195 35445 11207 35479
rect 11149 35439 11207 35445
rect 11790 35436 11796 35488
rect 11848 35436 11854 35488
rect 20456 35476 20484 35516
rect 20622 35504 20628 35556
rect 20680 35544 20686 35556
rect 22005 35547 22063 35553
rect 22005 35544 22017 35547
rect 20680 35516 22017 35544
rect 20680 35504 20686 35516
rect 22005 35513 22017 35516
rect 22051 35513 22063 35547
rect 22005 35507 22063 35513
rect 20717 35479 20775 35485
rect 20717 35476 20729 35479
rect 20456 35448 20729 35476
rect 20717 35445 20729 35448
rect 20763 35445 20775 35479
rect 20717 35439 20775 35445
rect 24489 35479 24547 35485
rect 24489 35445 24501 35479
rect 24535 35476 24547 35479
rect 24578 35476 24584 35488
rect 24535 35448 24584 35476
rect 24535 35445 24547 35448
rect 24489 35439 24547 35445
rect 24578 35436 24584 35448
rect 24636 35436 24642 35488
rect 25133 35479 25191 35485
rect 25133 35445 25145 35479
rect 25179 35476 25191 35479
rect 26050 35476 26056 35488
rect 25179 35448 26056 35476
rect 25179 35445 25191 35448
rect 25133 35439 25191 35445
rect 26050 35436 26056 35448
rect 26108 35436 26114 35488
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 25314 35232 25320 35284
rect 25372 35232 25378 35284
rect 22738 35096 22744 35148
rect 22796 35136 22802 35148
rect 23293 35139 23351 35145
rect 23293 35136 23305 35139
rect 22796 35108 23305 35136
rect 22796 35096 22802 35108
rect 23293 35105 23305 35108
rect 23339 35105 23351 35139
rect 23293 35099 23351 35105
rect 24213 35071 24271 35077
rect 24213 35037 24225 35071
rect 24259 35068 24271 35071
rect 24673 35071 24731 35077
rect 24673 35068 24685 35071
rect 24259 35040 24685 35068
rect 24259 35037 24271 35040
rect 24213 35031 24271 35037
rect 24673 35037 24685 35040
rect 24719 35068 24731 35071
rect 24854 35068 24860 35080
rect 24719 35040 24860 35068
rect 24719 35037 24731 35040
rect 24673 35031 24731 35037
rect 24854 35028 24860 35040
rect 24912 35028 24918 35080
rect 23109 35003 23167 35009
rect 23109 35000 23121 35003
rect 22388 34972 23121 35000
rect 21913 34935 21971 34941
rect 21913 34901 21925 34935
rect 21959 34932 21971 34935
rect 22002 34932 22008 34944
rect 21959 34904 22008 34932
rect 21959 34901 21971 34904
rect 21913 34895 21971 34901
rect 22002 34892 22008 34904
rect 22060 34892 22066 34944
rect 22186 34892 22192 34944
rect 22244 34932 22250 34944
rect 22388 34941 22416 34972
rect 23109 34969 23121 34972
rect 23155 34969 23167 35003
rect 23109 34963 23167 34969
rect 23201 35003 23259 35009
rect 23201 34969 23213 35003
rect 23247 35000 23259 35003
rect 25222 35000 25228 35012
rect 23247 34972 25228 35000
rect 23247 34969 23259 34972
rect 23201 34963 23259 34969
rect 25222 34960 25228 34972
rect 25280 34960 25286 35012
rect 22373 34935 22431 34941
rect 22373 34932 22385 34935
rect 22244 34904 22385 34932
rect 22244 34892 22250 34904
rect 22373 34901 22385 34904
rect 22419 34901 22431 34935
rect 22373 34895 22431 34901
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22741 34935 22799 34941
rect 22741 34932 22753 34935
rect 22520 34904 22753 34932
rect 22520 34892 22526 34904
rect 22741 34901 22753 34904
rect 22787 34901 22799 34935
rect 22741 34895 22799 34901
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 21082 34688 21088 34740
rect 21140 34728 21146 34740
rect 21453 34731 21511 34737
rect 21453 34728 21465 34731
rect 21140 34700 21465 34728
rect 21140 34688 21146 34700
rect 21453 34697 21465 34700
rect 21499 34697 21511 34731
rect 21453 34691 21511 34697
rect 25133 34731 25191 34737
rect 25133 34697 25145 34731
rect 25179 34728 25191 34731
rect 25222 34728 25228 34740
rect 25179 34700 25228 34728
rect 25179 34697 25191 34700
rect 25133 34691 25191 34697
rect 25222 34688 25228 34700
rect 25280 34688 25286 34740
rect 24857 34595 24915 34601
rect 24857 34561 24869 34595
rect 24903 34592 24915 34595
rect 25314 34592 25320 34604
rect 24903 34564 25320 34592
rect 24903 34561 24915 34564
rect 24857 34555 24915 34561
rect 25314 34552 25320 34564
rect 25372 34552 25378 34604
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 9125 34187 9183 34193
rect 9125 34153 9137 34187
rect 9171 34184 9183 34187
rect 9306 34184 9312 34196
rect 9171 34156 9312 34184
rect 9171 34153 9183 34156
rect 9125 34147 9183 34153
rect 9306 34144 9312 34156
rect 9364 34144 9370 34196
rect 21900 34187 21958 34193
rect 21900 34153 21912 34187
rect 21946 34184 21958 34187
rect 23014 34184 23020 34196
rect 21946 34156 23020 34184
rect 21946 34153 21958 34156
rect 21900 34147 21958 34153
rect 23014 34144 23020 34156
rect 23072 34144 23078 34196
rect 11790 34008 11796 34060
rect 11848 34048 11854 34060
rect 15381 34051 15439 34057
rect 15381 34048 15393 34051
rect 11848 34020 15393 34048
rect 11848 34008 11854 34020
rect 15381 34017 15393 34020
rect 15427 34017 15439 34051
rect 15381 34011 15439 34017
rect 19702 34008 19708 34060
rect 19760 34048 19766 34060
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 19760 34020 21649 34048
rect 19760 34008 19766 34020
rect 21637 34017 21649 34020
rect 21683 34048 21695 34051
rect 22278 34048 22284 34060
rect 21683 34020 22284 34048
rect 21683 34017 21695 34020
rect 21637 34011 21695 34017
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 9214 33940 9220 33992
rect 9272 33980 9278 33992
rect 9309 33983 9367 33989
rect 9309 33980 9321 33983
rect 9272 33952 9321 33980
rect 9272 33940 9278 33952
rect 9309 33949 9321 33952
rect 9355 33949 9367 33983
rect 9309 33943 9367 33949
rect 19426 33940 19432 33992
rect 19484 33940 19490 33992
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33980 24915 33983
rect 25314 33980 25320 33992
rect 24903 33952 25320 33980
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 14645 33915 14703 33921
rect 14645 33881 14657 33915
rect 14691 33912 14703 33915
rect 15378 33912 15384 33924
rect 14691 33884 15384 33912
rect 14691 33881 14703 33884
rect 14645 33875 14703 33881
rect 15378 33872 15384 33884
rect 15436 33912 15442 33924
rect 15841 33915 15899 33921
rect 15841 33912 15853 33915
rect 15436 33884 15853 33912
rect 15436 33872 15442 33884
rect 15841 33881 15853 33884
rect 15887 33881 15899 33915
rect 15841 33875 15899 33881
rect 19705 33915 19763 33921
rect 19705 33881 19717 33915
rect 19751 33912 19763 33915
rect 19978 33912 19984 33924
rect 19751 33884 19984 33912
rect 19751 33881 19763 33884
rect 19705 33875 19763 33881
rect 19978 33872 19984 33884
rect 20036 33872 20042 33924
rect 21082 33912 21088 33924
rect 20930 33884 21088 33912
rect 21082 33872 21088 33884
rect 21140 33912 21146 33924
rect 22370 33912 22376 33924
rect 21140 33884 22376 33912
rect 21140 33872 21146 33884
rect 22370 33872 22376 33884
rect 22428 33872 22434 33924
rect 19061 33847 19119 33853
rect 19061 33813 19073 33847
rect 19107 33844 19119 33847
rect 19242 33844 19248 33856
rect 19107 33816 19248 33844
rect 19107 33813 19119 33816
rect 19061 33807 19119 33813
rect 19242 33804 19248 33816
rect 19300 33804 19306 33856
rect 21174 33804 21180 33856
rect 21232 33804 21238 33856
rect 23198 33804 23204 33856
rect 23256 33844 23262 33856
rect 23385 33847 23443 33853
rect 23385 33844 23397 33847
rect 23256 33816 23397 33844
rect 23256 33804 23262 33816
rect 23385 33813 23397 33816
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 24210 33804 24216 33856
rect 24268 33844 24274 33856
rect 25133 33847 25191 33853
rect 25133 33844 25145 33847
rect 24268 33816 25145 33844
rect 24268 33804 24274 33816
rect 25133 33813 25145 33816
rect 25179 33813 25191 33847
rect 25133 33807 25191 33813
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 22554 33640 22560 33652
rect 19812 33612 22560 33640
rect 19812 33581 19840 33612
rect 22554 33600 22560 33612
rect 22612 33640 22618 33652
rect 23198 33640 23204 33652
rect 22612 33612 23204 33640
rect 22612 33600 22618 33612
rect 23198 33600 23204 33612
rect 23256 33600 23262 33652
rect 23566 33600 23572 33652
rect 23624 33640 23630 33652
rect 25133 33643 25191 33649
rect 25133 33640 25145 33643
rect 23624 33612 25145 33640
rect 23624 33600 23630 33612
rect 25133 33609 25145 33612
rect 25179 33609 25191 33643
rect 25133 33603 25191 33609
rect 19797 33575 19855 33581
rect 19797 33541 19809 33575
rect 19843 33541 19855 33575
rect 21082 33572 21088 33584
rect 21022 33544 21088 33572
rect 19797 33535 19855 33541
rect 21082 33532 21088 33544
rect 21140 33572 21146 33584
rect 21545 33575 21603 33581
rect 21545 33572 21557 33575
rect 21140 33544 21557 33572
rect 21140 33532 21146 33544
rect 21545 33541 21557 33544
rect 21591 33572 21603 33575
rect 21910 33572 21916 33584
rect 21591 33544 21916 33572
rect 21591 33541 21603 33544
rect 21545 33535 21603 33541
rect 21910 33532 21916 33544
rect 21968 33532 21974 33584
rect 22278 33572 22284 33584
rect 22020 33544 22284 33572
rect 19518 33464 19524 33516
rect 19576 33464 19582 33516
rect 22020 33513 22048 33544
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 22370 33532 22376 33584
rect 22428 33572 22434 33584
rect 22428 33544 22770 33572
rect 22428 33532 22434 33544
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33473 22063 33507
rect 25317 33507 25375 33513
rect 25317 33504 25329 33507
rect 22005 33467 22063 33473
rect 24872 33476 25329 33504
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 22370 33436 22376 33448
rect 22327 33408 22376 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 23014 33396 23020 33448
rect 23072 33436 23078 33448
rect 23753 33439 23811 33445
rect 23753 33436 23765 33439
rect 23072 33408 23765 33436
rect 23072 33396 23078 33408
rect 23753 33405 23765 33408
rect 23799 33405 23811 33439
rect 23753 33399 23811 33405
rect 19242 33260 19248 33312
rect 19300 33260 19306 33312
rect 19978 33260 19984 33312
rect 20036 33300 20042 33312
rect 20530 33300 20536 33312
rect 20036 33272 20536 33300
rect 20036 33260 20042 33272
rect 20530 33260 20536 33272
rect 20588 33300 20594 33312
rect 21269 33303 21327 33309
rect 21269 33300 21281 33303
rect 20588 33272 21281 33300
rect 20588 33260 20594 33272
rect 21269 33269 21281 33272
rect 21315 33269 21327 33303
rect 21269 33263 21327 33269
rect 23842 33260 23848 33312
rect 23900 33300 23906 33312
rect 24397 33303 24455 33309
rect 24397 33300 24409 33303
rect 23900 33272 24409 33300
rect 23900 33260 23906 33272
rect 24397 33269 24409 33272
rect 24443 33269 24455 33303
rect 24397 33263 24455 33269
rect 24762 33260 24768 33312
rect 24820 33300 24826 33312
rect 24872 33309 24900 33476
rect 25317 33473 25329 33476
rect 25363 33473 25375 33507
rect 25317 33467 25375 33473
rect 24857 33303 24915 33309
rect 24857 33300 24869 33303
rect 24820 33272 24869 33300
rect 24820 33260 24826 33272
rect 24857 33269 24869 33272
rect 24903 33269 24915 33303
rect 24857 33263 24915 33269
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 16574 33096 16580 33108
rect 16040 33068 16580 33096
rect 16040 32969 16068 33068
rect 16574 33056 16580 33068
rect 16632 33056 16638 33108
rect 16669 33099 16727 33105
rect 16669 33065 16681 33099
rect 16715 33096 16727 33099
rect 21358 33096 21364 33108
rect 16715 33068 21364 33096
rect 16715 33065 16727 33068
rect 16669 33059 16727 33065
rect 16025 32963 16083 32969
rect 16025 32929 16037 32963
rect 16071 32929 16083 32963
rect 16025 32923 16083 32929
rect 16114 32920 16120 32972
rect 16172 32960 16178 32972
rect 16684 32960 16712 33059
rect 21358 33056 21364 33068
rect 21416 33056 21422 33108
rect 21910 33056 21916 33108
rect 21968 33056 21974 33108
rect 22370 33056 22376 33108
rect 22428 33096 22434 33108
rect 22738 33096 22744 33108
rect 22428 33068 22744 33096
rect 22428 33056 22434 33068
rect 22738 33056 22744 33068
rect 22796 33096 22802 33108
rect 24029 33099 24087 33105
rect 24029 33096 24041 33099
rect 22796 33068 24041 33096
rect 22796 33056 22802 33068
rect 24029 33065 24041 33068
rect 24075 33065 24087 33099
rect 24029 33059 24087 33065
rect 19613 33031 19671 33037
rect 19613 32997 19625 33031
rect 19659 33028 19671 33031
rect 19886 33028 19892 33040
rect 19659 33000 19892 33028
rect 19659 32997 19671 33000
rect 19613 32991 19671 32997
rect 19886 32988 19892 33000
rect 19944 33028 19950 33040
rect 21818 33028 21824 33040
rect 19944 33000 21824 33028
rect 19944 32988 19950 33000
rect 21818 32988 21824 33000
rect 21876 32988 21882 33040
rect 16172 32932 16712 32960
rect 17037 32963 17095 32969
rect 16172 32920 16178 32932
rect 17037 32929 17049 32963
rect 17083 32960 17095 32963
rect 17083 32932 21864 32960
rect 17083 32929 17095 32932
rect 17037 32923 17095 32929
rect 16574 32852 16580 32904
rect 16632 32892 16638 32904
rect 16761 32895 16819 32901
rect 16761 32892 16773 32895
rect 16632 32864 16773 32892
rect 16632 32852 16638 32864
rect 16761 32861 16773 32864
rect 16807 32892 16819 32895
rect 17310 32892 17316 32904
rect 16807 32864 17316 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 17310 32852 17316 32864
rect 17368 32852 17374 32904
rect 15933 32827 15991 32833
rect 15933 32793 15945 32827
rect 15979 32824 15991 32827
rect 17218 32824 17224 32836
rect 15979 32796 17224 32824
rect 15979 32793 15991 32796
rect 15933 32787 15991 32793
rect 17218 32784 17224 32796
rect 17276 32824 17282 32836
rect 17420 32824 17448 32932
rect 19426 32852 19432 32904
rect 19484 32892 19490 32904
rect 20625 32895 20683 32901
rect 20625 32892 20637 32895
rect 19484 32864 20637 32892
rect 19484 32852 19490 32864
rect 20625 32861 20637 32864
rect 20671 32861 20683 32895
rect 20625 32855 20683 32861
rect 17276 32796 17448 32824
rect 17276 32784 17282 32796
rect 17494 32784 17500 32836
rect 17552 32824 17558 32836
rect 19886 32824 19892 32836
rect 17552 32796 19892 32824
rect 17552 32784 17558 32796
rect 19886 32784 19892 32796
rect 19944 32784 19950 32836
rect 12618 32716 12624 32768
rect 12676 32756 12682 32768
rect 15565 32759 15623 32765
rect 15565 32756 15577 32759
rect 12676 32728 15577 32756
rect 12676 32716 12682 32728
rect 15565 32725 15577 32728
rect 15611 32725 15623 32759
rect 21836 32756 21864 32932
rect 22278 32920 22284 32972
rect 22336 32920 22342 32972
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 25130 32960 25136 32972
rect 22603 32932 25136 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 25130 32920 25136 32932
rect 25188 32920 25194 32972
rect 25222 32920 25228 32972
rect 25280 32920 25286 32972
rect 25041 32895 25099 32901
rect 25041 32861 25053 32895
rect 25087 32892 25099 32895
rect 25406 32892 25412 32904
rect 25087 32864 25412 32892
rect 25087 32861 25099 32864
rect 25041 32855 25099 32861
rect 25406 32852 25412 32864
rect 25464 32852 25470 32904
rect 21910 32784 21916 32836
rect 21968 32824 21974 32836
rect 21968 32796 23046 32824
rect 21968 32784 21974 32796
rect 23842 32784 23848 32836
rect 23900 32824 23906 32836
rect 24949 32827 25007 32833
rect 24949 32824 24961 32827
rect 23900 32796 24961 32824
rect 23900 32784 23906 32796
rect 24949 32793 24961 32796
rect 24995 32793 25007 32827
rect 24949 32787 25007 32793
rect 23474 32756 23480 32768
rect 21836 32728 23480 32756
rect 15565 32719 15623 32725
rect 23474 32716 23480 32728
rect 23532 32716 23538 32768
rect 24581 32759 24639 32765
rect 24581 32725 24593 32759
rect 24627 32756 24639 32759
rect 24854 32756 24860 32768
rect 24627 32728 24860 32756
rect 24627 32725 24639 32728
rect 24581 32719 24639 32725
rect 24854 32716 24860 32728
rect 24912 32716 24918 32768
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 17037 32555 17095 32561
rect 17037 32521 17049 32555
rect 17083 32552 17095 32555
rect 17494 32552 17500 32564
rect 17083 32524 17500 32552
rect 17083 32521 17095 32524
rect 17037 32515 17095 32521
rect 15378 32444 15384 32496
rect 15436 32484 15442 32496
rect 15436 32456 16574 32484
rect 15436 32444 15442 32456
rect 16546 32416 16574 32456
rect 17052 32416 17080 32515
rect 17494 32512 17500 32524
rect 17552 32512 17558 32564
rect 18785 32555 18843 32561
rect 18785 32521 18797 32555
rect 18831 32552 18843 32555
rect 19242 32552 19248 32564
rect 18831 32524 19248 32552
rect 18831 32521 18843 32524
rect 18785 32515 18843 32521
rect 19242 32512 19248 32524
rect 19300 32552 19306 32564
rect 19300 32524 20668 32552
rect 19300 32512 19306 32524
rect 17586 32444 17592 32496
rect 17644 32484 17650 32496
rect 19610 32484 19616 32496
rect 17644 32456 19616 32484
rect 17644 32444 17650 32456
rect 19610 32444 19616 32456
rect 19668 32444 19674 32496
rect 20640 32484 20668 32524
rect 25130 32512 25136 32564
rect 25188 32552 25194 32564
rect 25225 32555 25283 32561
rect 25225 32552 25237 32555
rect 25188 32524 25237 32552
rect 25188 32512 25194 32524
rect 25225 32521 25237 32524
rect 25271 32552 25283 32555
rect 25406 32552 25412 32564
rect 25271 32524 25412 32552
rect 25271 32521 25283 32524
rect 25225 32515 25283 32521
rect 25406 32512 25412 32524
rect 25464 32512 25470 32564
rect 21082 32484 21088 32496
rect 20562 32456 21088 32484
rect 21082 32444 21088 32456
rect 21140 32444 21146 32496
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 22833 32487 22891 32493
rect 22833 32484 22845 32487
rect 22336 32456 22845 32484
rect 22336 32444 22342 32456
rect 22833 32453 22845 32456
rect 22879 32484 22891 32487
rect 22879 32456 23520 32484
rect 22879 32453 22891 32456
rect 22833 32447 22891 32453
rect 16546 32388 17080 32416
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 23492 32425 23520 32456
rect 24026 32444 24032 32496
rect 24084 32484 24090 32496
rect 24084 32456 24242 32484
rect 24084 32444 24090 32456
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 21876 32388 22109 32416
rect 21876 32376 21882 32388
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 13354 32308 13360 32360
rect 13412 32348 13418 32360
rect 16117 32351 16175 32357
rect 16117 32348 16129 32351
rect 13412 32320 16129 32348
rect 13412 32308 13418 32320
rect 16117 32317 16129 32320
rect 16163 32348 16175 32351
rect 16758 32348 16764 32360
rect 16163 32320 16764 32348
rect 16163 32317 16175 32320
rect 16117 32311 16175 32317
rect 16758 32308 16764 32320
rect 16816 32308 16822 32360
rect 16853 32351 16911 32357
rect 16853 32317 16865 32351
rect 16899 32348 16911 32351
rect 17126 32348 17132 32360
rect 16899 32320 17132 32348
rect 16899 32317 16911 32320
rect 16853 32311 16911 32317
rect 17126 32308 17132 32320
rect 17184 32308 17190 32360
rect 19061 32351 19119 32357
rect 19061 32317 19073 32351
rect 19107 32317 19119 32351
rect 19061 32311 19119 32317
rect 19337 32351 19395 32357
rect 19337 32317 19349 32351
rect 19383 32348 19395 32351
rect 21174 32348 21180 32360
rect 19383 32320 21180 32348
rect 19383 32317 19395 32320
rect 19337 32311 19395 32317
rect 19076 32212 19104 32311
rect 21174 32308 21180 32320
rect 21232 32308 21238 32360
rect 23753 32351 23811 32357
rect 23753 32317 23765 32351
rect 23799 32348 23811 32351
rect 25222 32348 25228 32360
rect 23799 32320 25228 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 20364 32252 21956 32280
rect 19426 32212 19432 32224
rect 19076 32184 19432 32212
rect 19426 32172 19432 32184
rect 19484 32172 19490 32224
rect 19702 32172 19708 32224
rect 19760 32212 19766 32224
rect 20364 32212 20392 32252
rect 19760 32184 20392 32212
rect 20809 32215 20867 32221
rect 19760 32172 19766 32184
rect 20809 32181 20821 32215
rect 20855 32212 20867 32215
rect 20898 32212 20904 32224
rect 20855 32184 20904 32212
rect 20855 32181 20867 32184
rect 20809 32175 20867 32181
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21637 32215 21695 32221
rect 21637 32181 21649 32215
rect 21683 32212 21695 32215
rect 21818 32212 21824 32224
rect 21683 32184 21824 32212
rect 21683 32181 21695 32184
rect 21637 32175 21695 32181
rect 21818 32172 21824 32184
rect 21876 32172 21882 32224
rect 21928 32212 21956 32252
rect 25958 32212 25964 32224
rect 21928 32184 25964 32212
rect 25958 32172 25964 32184
rect 26016 32172 26022 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 9490 31968 9496 32020
rect 9548 32008 9554 32020
rect 16482 32008 16488 32020
rect 9548 31980 16488 32008
rect 9548 31968 9554 31980
rect 16482 31968 16488 31980
rect 16540 31968 16546 32020
rect 17024 32011 17082 32017
rect 17024 31977 17036 32011
rect 17070 32008 17082 32011
rect 18506 32008 18512 32020
rect 17070 31980 18512 32008
rect 17070 31977 17082 31980
rect 17024 31971 17082 31977
rect 18506 31968 18512 31980
rect 18564 31968 18570 32020
rect 18877 32011 18935 32017
rect 18877 31977 18889 32011
rect 18923 32008 18935 32011
rect 19061 32011 19119 32017
rect 19061 32008 19073 32011
rect 18923 31980 19073 32008
rect 18923 31977 18935 31980
rect 18877 31971 18935 31977
rect 19061 31977 19073 31980
rect 19107 32008 19119 32011
rect 19242 32008 19248 32020
rect 19107 31980 19248 32008
rect 19107 31977 19119 31980
rect 19061 31971 19119 31977
rect 19242 31968 19248 31980
rect 19300 31968 19306 32020
rect 24026 31968 24032 32020
rect 24084 31968 24090 32020
rect 24854 31968 24860 32020
rect 24912 32008 24918 32020
rect 25314 32008 25320 32020
rect 24912 31980 25320 32008
rect 24912 31968 24918 31980
rect 25314 31968 25320 31980
rect 25372 31968 25378 32020
rect 12526 31900 12532 31952
rect 12584 31940 12590 31952
rect 15565 31943 15623 31949
rect 15565 31940 15577 31943
rect 12584 31912 15577 31940
rect 12584 31900 12590 31912
rect 15565 31909 15577 31912
rect 15611 31909 15623 31943
rect 15565 31903 15623 31909
rect 20806 31900 20812 31952
rect 20864 31940 20870 31952
rect 21637 31943 21695 31949
rect 21637 31940 21649 31943
rect 20864 31912 21649 31940
rect 20864 31900 20870 31912
rect 21637 31909 21649 31912
rect 21683 31909 21695 31943
rect 21637 31903 21695 31909
rect 22738 31900 22744 31952
rect 22796 31940 22802 31952
rect 23017 31943 23075 31949
rect 23017 31940 23029 31943
rect 22796 31912 23029 31940
rect 22796 31900 22802 31912
rect 23017 31909 23029 31912
rect 23063 31909 23075 31943
rect 24118 31940 24124 31952
rect 23017 31903 23075 31909
rect 23124 31912 24124 31940
rect 16114 31832 16120 31884
rect 16172 31832 16178 31884
rect 16666 31872 16672 31884
rect 16546 31844 16672 31872
rect 16025 31807 16083 31813
rect 16025 31773 16037 31807
rect 16071 31804 16083 31807
rect 16546 31804 16574 31844
rect 16666 31832 16672 31844
rect 16724 31872 16730 31884
rect 17586 31872 17592 31884
rect 16724 31844 17592 31872
rect 16724 31832 16730 31844
rect 17586 31832 17592 31844
rect 17644 31832 17650 31884
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 18509 31875 18567 31881
rect 18509 31872 18521 31875
rect 17736 31844 18521 31872
rect 17736 31832 17742 31844
rect 18509 31841 18521 31844
rect 18555 31841 18567 31875
rect 18509 31835 18567 31841
rect 19702 31832 19708 31884
rect 19760 31872 19766 31884
rect 22189 31875 22247 31881
rect 22189 31872 22201 31875
rect 19760 31844 22201 31872
rect 19760 31832 19766 31844
rect 22189 31841 22201 31844
rect 22235 31841 22247 31875
rect 23124 31872 23152 31912
rect 24118 31900 24124 31912
rect 24176 31900 24182 31952
rect 25038 31900 25044 31952
rect 25096 31940 25102 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 25096 31912 25145 31940
rect 25096 31900 25102 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 25133 31903 25191 31909
rect 22189 31835 22247 31841
rect 22940 31844 23152 31872
rect 16071 31776 16574 31804
rect 16071 31773 16083 31776
rect 16025 31767 16083 31773
rect 16758 31764 16764 31816
rect 16816 31764 16822 31816
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 21082 31804 21088 31816
rect 20838 31776 21088 31804
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 22097 31807 22155 31813
rect 22097 31773 22109 31807
rect 22143 31804 22155 31807
rect 22940 31804 22968 31844
rect 23290 31832 23296 31884
rect 23348 31872 23354 31884
rect 23477 31875 23535 31881
rect 23477 31872 23489 31875
rect 23348 31844 23489 31872
rect 23348 31832 23354 31844
rect 23477 31841 23489 31844
rect 23523 31841 23535 31875
rect 23477 31835 23535 31841
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31841 23627 31875
rect 23569 31835 23627 31841
rect 22143 31776 22968 31804
rect 22143 31773 22155 31776
rect 22097 31767 22155 31773
rect 23014 31764 23020 31816
rect 23072 31804 23078 31816
rect 23584 31804 23612 31835
rect 23072 31776 23612 31804
rect 24857 31807 24915 31813
rect 23072 31764 23078 31776
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 19242 31736 19248 31748
rect 18262 31708 19248 31736
rect 19242 31696 19248 31708
rect 19300 31696 19306 31748
rect 15933 31671 15991 31677
rect 15933 31637 15945 31671
rect 15979 31668 15991 31671
rect 17126 31668 17132 31680
rect 15979 31640 17132 31668
rect 15979 31637 15991 31640
rect 15933 31631 15991 31637
rect 17126 31628 17132 31640
rect 17184 31628 17190 31680
rect 20990 31628 20996 31680
rect 21048 31668 21054 31680
rect 21177 31671 21235 31677
rect 21177 31668 21189 31671
rect 21048 31640 21189 31668
rect 21048 31628 21054 31640
rect 21177 31637 21189 31640
rect 21223 31637 21235 31671
rect 21177 31631 21235 31637
rect 22002 31628 22008 31680
rect 22060 31628 22066 31680
rect 22094 31628 22100 31680
rect 22152 31668 22158 31680
rect 22554 31668 22560 31680
rect 22152 31640 22560 31668
rect 22152 31628 22158 31640
rect 22554 31628 22560 31640
rect 22612 31668 22618 31680
rect 22649 31671 22707 31677
rect 22649 31668 22661 31671
rect 22612 31640 22661 31668
rect 22612 31628 22618 31640
rect 22649 31637 22661 31640
rect 22695 31668 22707 31671
rect 23385 31671 23443 31677
rect 23385 31668 23397 31671
rect 22695 31640 23397 31668
rect 22695 31637 22707 31640
rect 22649 31631 22707 31637
rect 23385 31637 23397 31640
rect 23431 31637 23443 31671
rect 23385 31631 23443 31637
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 16666 31424 16672 31476
rect 16724 31424 16730 31476
rect 19153 31467 19211 31473
rect 19153 31433 19165 31467
rect 19199 31464 19211 31467
rect 19702 31464 19708 31476
rect 19199 31436 19708 31464
rect 19199 31433 19211 31436
rect 19153 31427 19211 31433
rect 19702 31424 19708 31436
rect 19760 31424 19766 31476
rect 20533 31467 20591 31473
rect 20533 31433 20545 31467
rect 20579 31464 20591 31467
rect 25130 31464 25136 31476
rect 20579 31436 25136 31464
rect 20579 31433 20591 31436
rect 20533 31427 20591 31433
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 25498 31424 25504 31476
rect 25556 31464 25562 31476
rect 26142 31464 26148 31476
rect 25556 31436 26148 31464
rect 25556 31424 25562 31436
rect 26142 31424 26148 31436
rect 26200 31424 26206 31476
rect 15010 31396 15016 31408
rect 14858 31368 15016 31396
rect 15010 31356 15016 31368
rect 15068 31356 15074 31408
rect 19242 31396 19248 31408
rect 18906 31368 19248 31396
rect 19242 31356 19248 31368
rect 19300 31396 19306 31408
rect 19429 31399 19487 31405
rect 19429 31396 19441 31399
rect 19300 31368 19441 31396
rect 19300 31356 19306 31368
rect 19429 31365 19441 31368
rect 19475 31365 19487 31399
rect 19429 31359 19487 31365
rect 22646 31356 22652 31408
rect 22704 31396 22710 31408
rect 22741 31399 22799 31405
rect 22741 31396 22753 31399
rect 22704 31368 22753 31396
rect 22704 31356 22710 31368
rect 22741 31365 22753 31368
rect 22787 31396 22799 31399
rect 23014 31396 23020 31408
rect 22787 31368 23020 31396
rect 22787 31365 22799 31368
rect 22741 31359 22799 31365
rect 23014 31356 23020 31368
rect 23072 31356 23078 31408
rect 24026 31396 24032 31408
rect 23966 31368 24032 31396
rect 24026 31356 24032 31368
rect 24084 31356 24090 31408
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 17405 31331 17463 31337
rect 17405 31328 17417 31331
rect 16816 31300 17417 31328
rect 16816 31288 16822 31300
rect 17405 31297 17417 31300
rect 17451 31297 17463 31331
rect 17405 31291 17463 31297
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31328 19855 31331
rect 20441 31331 20499 31337
rect 20441 31328 20453 31331
rect 19843 31300 20453 31328
rect 19843 31297 19855 31300
rect 19797 31291 19855 31297
rect 20441 31297 20453 31300
rect 20487 31328 20499 31331
rect 21910 31328 21916 31340
rect 20487 31300 21916 31328
rect 20487 31297 20499 31300
rect 20441 31291 20499 31297
rect 21910 31288 21916 31300
rect 21968 31288 21974 31340
rect 22278 31288 22284 31340
rect 22336 31328 22342 31340
rect 22465 31331 22523 31337
rect 22465 31328 22477 31331
rect 22336 31300 22477 31328
rect 22336 31288 22342 31300
rect 22465 31297 22477 31300
rect 22511 31297 22523 31331
rect 22465 31291 22523 31297
rect 25317 31331 25375 31337
rect 25317 31297 25329 31331
rect 25363 31328 25375 31331
rect 25498 31328 25504 31340
rect 25363 31300 25504 31328
rect 25363 31297 25375 31300
rect 25317 31291 25375 31297
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 13354 31220 13360 31272
rect 13412 31220 13418 31272
rect 13633 31263 13691 31269
rect 13633 31229 13645 31263
rect 13679 31260 13691 31263
rect 15473 31263 15531 31269
rect 15473 31260 15485 31263
rect 13679 31232 15485 31260
rect 13679 31229 13691 31232
rect 13633 31223 13691 31229
rect 15473 31229 15485 31232
rect 15519 31260 15531 31263
rect 16114 31260 16120 31272
rect 15519 31232 16120 31260
rect 15519 31229 15531 31232
rect 15473 31223 15531 31229
rect 16114 31220 16120 31232
rect 16172 31260 16178 31272
rect 16393 31263 16451 31269
rect 16393 31260 16405 31263
rect 16172 31232 16405 31260
rect 16172 31220 16178 31232
rect 16393 31229 16405 31232
rect 16439 31229 16451 31263
rect 16393 31223 16451 31229
rect 17678 31220 17684 31272
rect 17736 31220 17742 31272
rect 18690 31220 18696 31272
rect 18748 31260 18754 31272
rect 20625 31263 20683 31269
rect 20625 31260 20637 31263
rect 18748 31232 20637 31260
rect 18748 31220 18754 31232
rect 20625 31229 20637 31232
rect 20671 31229 20683 31263
rect 20625 31223 20683 31229
rect 22189 31263 22247 31269
rect 22189 31229 22201 31263
rect 22235 31260 22247 31263
rect 22370 31260 22376 31272
rect 22235 31232 22376 31260
rect 22235 31229 22247 31232
rect 22189 31223 22247 31229
rect 22370 31220 22376 31232
rect 22428 31220 22434 31272
rect 15010 31152 15016 31204
rect 15068 31192 15074 31204
rect 21545 31195 21603 31201
rect 15068 31164 15792 31192
rect 15068 31152 15074 31164
rect 13814 31084 13820 31136
rect 13872 31124 13878 31136
rect 15764 31133 15792 31164
rect 21545 31161 21557 31195
rect 21591 31192 21603 31195
rect 22002 31192 22008 31204
rect 21591 31164 22008 31192
rect 21591 31161 21603 31164
rect 21545 31155 21603 31161
rect 22002 31152 22008 31164
rect 22060 31192 22066 31204
rect 22278 31192 22284 31204
rect 22060 31164 22284 31192
rect 22060 31152 22066 31164
rect 22278 31152 22284 31164
rect 22336 31152 22342 31204
rect 15105 31127 15163 31133
rect 15105 31124 15117 31127
rect 13872 31096 15117 31124
rect 13872 31084 13878 31096
rect 15105 31093 15117 31096
rect 15151 31093 15163 31127
rect 15105 31087 15163 31093
rect 15749 31127 15807 31133
rect 15749 31093 15761 31127
rect 15795 31124 15807 31127
rect 18414 31124 18420 31136
rect 15795 31096 18420 31124
rect 15795 31093 15807 31096
rect 15749 31087 15807 31093
rect 18414 31084 18420 31096
rect 18472 31084 18478 31136
rect 19886 31084 19892 31136
rect 19944 31124 19950 31136
rect 20073 31127 20131 31133
rect 20073 31124 20085 31127
rect 19944 31096 20085 31124
rect 19944 31084 19950 31096
rect 20073 31093 20085 31096
rect 20119 31093 20131 31127
rect 20073 31087 20131 31093
rect 21910 31084 21916 31136
rect 21968 31124 21974 31136
rect 22186 31124 22192 31136
rect 21968 31096 22192 31124
rect 21968 31084 21974 31096
rect 22186 31084 22192 31096
rect 22244 31084 22250 31136
rect 23474 31084 23480 31136
rect 23532 31124 23538 31136
rect 24213 31127 24271 31133
rect 24213 31124 24225 31127
rect 23532 31096 24225 31124
rect 23532 31084 23538 31096
rect 24213 31093 24225 31096
rect 24259 31093 24271 31127
rect 24213 31087 24271 31093
rect 25130 31084 25136 31136
rect 25188 31084 25194 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 9125 30923 9183 30929
rect 9125 30889 9137 30923
rect 9171 30920 9183 30923
rect 10226 30920 10232 30932
rect 9171 30892 10232 30920
rect 9171 30889 9183 30892
rect 9125 30883 9183 30889
rect 10226 30880 10232 30892
rect 10284 30880 10290 30932
rect 15378 30880 15384 30932
rect 15436 30920 15442 30932
rect 15565 30923 15623 30929
rect 15565 30920 15577 30923
rect 15436 30892 15577 30920
rect 15436 30880 15442 30892
rect 15565 30889 15577 30892
rect 15611 30920 15623 30923
rect 15749 30923 15807 30929
rect 15749 30920 15761 30923
rect 15611 30892 15761 30920
rect 15611 30889 15623 30892
rect 15565 30883 15623 30889
rect 15749 30889 15761 30892
rect 15795 30889 15807 30923
rect 15749 30883 15807 30889
rect 18506 30880 18512 30932
rect 18564 30920 18570 30932
rect 18690 30920 18696 30932
rect 18564 30892 18696 30920
rect 18564 30880 18570 30892
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 18877 30923 18935 30929
rect 18877 30889 18889 30923
rect 18923 30920 18935 30923
rect 19242 30920 19248 30932
rect 18923 30892 19248 30920
rect 18923 30889 18935 30892
rect 18877 30883 18935 30889
rect 19242 30880 19248 30892
rect 19300 30920 19306 30932
rect 19705 30923 19763 30929
rect 19705 30920 19717 30923
rect 19300 30892 19717 30920
rect 19300 30880 19306 30892
rect 19705 30889 19717 30892
rect 19751 30889 19763 30923
rect 19705 30883 19763 30889
rect 22465 30923 22523 30929
rect 22465 30889 22477 30923
rect 22511 30920 22523 30923
rect 22646 30920 22652 30932
rect 22511 30892 22652 30920
rect 22511 30889 22523 30892
rect 22465 30883 22523 30889
rect 22646 30880 22652 30892
rect 22704 30880 22710 30932
rect 25498 30880 25504 30932
rect 25556 30880 25562 30932
rect 16761 30787 16819 30793
rect 16761 30753 16773 30787
rect 16807 30784 16819 30787
rect 19426 30784 19432 30796
rect 16807 30756 19432 30784
rect 16807 30753 16819 30756
rect 16761 30747 16819 30753
rect 19426 30744 19432 30756
rect 19484 30784 19490 30796
rect 20717 30787 20775 30793
rect 20717 30784 20729 30787
rect 19484 30756 20729 30784
rect 19484 30744 19490 30756
rect 20717 30753 20729 30756
rect 20763 30753 20775 30787
rect 20717 30747 20775 30753
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9309 30719 9367 30725
rect 9309 30716 9321 30719
rect 8812 30688 9321 30716
rect 8812 30676 8818 30688
rect 9309 30685 9321 30688
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 14090 30676 14096 30728
rect 14148 30716 14154 30728
rect 14369 30719 14427 30725
rect 14369 30716 14381 30719
rect 14148 30688 14381 30716
rect 14148 30676 14154 30688
rect 14369 30685 14381 30688
rect 14415 30716 14427 30719
rect 15378 30716 15384 30728
rect 14415 30688 15384 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 15378 30676 15384 30688
rect 15436 30676 15442 30728
rect 15102 30608 15108 30660
rect 15160 30608 15166 30660
rect 17037 30651 17095 30657
rect 17037 30617 17049 30651
rect 17083 30617 17095 30651
rect 18414 30648 18420 30660
rect 18262 30620 18420 30648
rect 17037 30611 17095 30617
rect 17052 30580 17080 30611
rect 18414 30608 18420 30620
rect 18472 30648 18478 30660
rect 19242 30648 19248 30660
rect 18472 30620 19248 30648
rect 18472 30608 18478 30620
rect 19242 30608 19248 30620
rect 19300 30608 19306 30660
rect 20990 30608 20996 30660
rect 21048 30608 21054 30660
rect 22370 30648 22376 30660
rect 22218 30620 22376 30648
rect 22370 30608 22376 30620
rect 22428 30648 22434 30660
rect 22428 30620 22600 30648
rect 22428 30608 22434 30620
rect 18690 30580 18696 30592
rect 17052 30552 18696 30580
rect 18690 30540 18696 30552
rect 18748 30540 18754 30592
rect 20070 30540 20076 30592
rect 20128 30540 20134 30592
rect 22572 30580 22600 30620
rect 22646 30608 22652 30660
rect 22704 30648 22710 30660
rect 24581 30651 24639 30657
rect 24581 30648 24593 30651
rect 22704 30620 24593 30648
rect 22704 30608 22710 30620
rect 24581 30617 24593 30620
rect 24627 30617 24639 30651
rect 24581 30611 24639 30617
rect 23201 30583 23259 30589
rect 23201 30580 23213 30583
rect 22572 30552 23213 30580
rect 23201 30549 23213 30552
rect 23247 30580 23259 30583
rect 24026 30580 24032 30592
rect 23247 30552 24032 30580
rect 23247 30549 23259 30552
rect 23201 30543 23259 30549
rect 24026 30540 24032 30552
rect 24084 30540 24090 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 13354 30376 13360 30388
rect 12406 30348 13360 30376
rect 12406 30308 12434 30348
rect 13354 30336 13360 30348
rect 13412 30336 13418 30388
rect 18969 30379 19027 30385
rect 18969 30345 18981 30379
rect 19015 30376 19027 30379
rect 19242 30376 19248 30388
rect 19015 30348 19248 30376
rect 19015 30345 19027 30348
rect 18969 30339 19027 30345
rect 19242 30336 19248 30348
rect 19300 30336 19306 30388
rect 20070 30336 20076 30388
rect 20128 30376 20134 30388
rect 20257 30379 20315 30385
rect 20257 30376 20269 30379
rect 20128 30348 20269 30376
rect 20128 30336 20134 30348
rect 20257 30345 20269 30348
rect 20303 30345 20315 30379
rect 20257 30339 20315 30345
rect 11808 30280 12434 30308
rect 7650 30200 7656 30252
rect 7708 30240 7714 30252
rect 11808 30249 11836 30280
rect 12710 30268 12716 30320
rect 12768 30268 12774 30320
rect 14090 30268 14096 30320
rect 14148 30268 14154 30320
rect 20349 30311 20407 30317
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 20622 30308 20628 30320
rect 20395 30280 20628 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 20622 30268 20628 30280
rect 20680 30268 20686 30320
rect 22462 30268 22468 30320
rect 22520 30268 22526 30320
rect 23474 30268 23480 30320
rect 23532 30308 23538 30320
rect 23569 30311 23627 30317
rect 23569 30308 23581 30311
rect 23532 30280 23581 30308
rect 23532 30268 23538 30280
rect 23569 30277 23581 30280
rect 23615 30277 23627 30311
rect 23569 30271 23627 30277
rect 24026 30268 24032 30320
rect 24084 30268 24090 30320
rect 9125 30243 9183 30249
rect 9125 30240 9137 30243
rect 7708 30212 9137 30240
rect 7708 30200 7714 30212
rect 9125 30209 9137 30212
rect 9171 30209 9183 30243
rect 9125 30203 9183 30209
rect 11793 30243 11851 30249
rect 11793 30209 11805 30243
rect 11839 30209 11851 30243
rect 11793 30203 11851 30209
rect 15841 30243 15899 30249
rect 15841 30209 15853 30243
rect 15887 30240 15899 30243
rect 16758 30240 16764 30252
rect 15887 30212 16764 30240
rect 15887 30209 15899 30212
rect 15841 30203 15899 30209
rect 16758 30200 16764 30212
rect 16816 30200 16822 30252
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 21315 30212 22385 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 12066 30132 12072 30184
rect 12124 30132 12130 30184
rect 12434 30132 12440 30184
rect 12492 30172 12498 30184
rect 12710 30172 12716 30184
rect 12492 30144 12716 30172
rect 12492 30132 12498 30144
rect 12710 30132 12716 30144
rect 12768 30132 12774 30184
rect 13354 30132 13360 30184
rect 13412 30172 13418 30184
rect 14829 30175 14887 30181
rect 14829 30172 14841 30175
rect 13412 30144 14841 30172
rect 13412 30132 13418 30144
rect 14829 30141 14841 30144
rect 14875 30141 14887 30175
rect 14829 30135 14887 30141
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30141 15991 30175
rect 15933 30135 15991 30141
rect 8938 30064 8944 30116
rect 8996 30064 9002 30116
rect 15948 30104 15976 30135
rect 16022 30132 16028 30184
rect 16080 30132 16086 30184
rect 16482 30132 16488 30184
rect 16540 30172 16546 30184
rect 16540 30144 17356 30172
rect 16540 30132 16546 30144
rect 17034 30104 17040 30116
rect 15948 30076 17040 30104
rect 16684 30048 16712 30076
rect 17034 30064 17040 30076
rect 17092 30064 17098 30116
rect 17328 30104 17356 30144
rect 20530 30132 20536 30184
rect 20588 30132 20594 30184
rect 22649 30175 22707 30181
rect 22649 30141 22661 30175
rect 22695 30172 22707 30175
rect 22830 30172 22836 30184
rect 22695 30144 22836 30172
rect 22695 30141 22707 30144
rect 22649 30135 22707 30141
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 23290 30132 23296 30184
rect 23348 30132 23354 30184
rect 23934 30172 23940 30184
rect 23400 30144 23940 30172
rect 23400 30104 23428 30144
rect 23934 30132 23940 30144
rect 23992 30132 23998 30184
rect 25041 30175 25099 30181
rect 25041 30141 25053 30175
rect 25087 30172 25099 30175
rect 25222 30172 25228 30184
rect 25087 30144 25228 30172
rect 25087 30141 25099 30144
rect 25041 30135 25099 30141
rect 25222 30132 25228 30144
rect 25280 30132 25286 30184
rect 17328 30076 23428 30104
rect 11514 29996 11520 30048
rect 11572 30036 11578 30048
rect 13541 30039 13599 30045
rect 13541 30036 13553 30039
rect 11572 30008 13553 30036
rect 11572 29996 11578 30008
rect 13541 30005 13553 30008
rect 13587 30036 13599 30039
rect 13630 30036 13636 30048
rect 13587 30008 13636 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 13630 29996 13636 30008
rect 13688 29996 13694 30048
rect 15473 30039 15531 30045
rect 15473 30005 15485 30039
rect 15519 30036 15531 30039
rect 15930 30036 15936 30048
rect 15519 30008 15936 30036
rect 15519 30005 15531 30008
rect 15473 29999 15531 30005
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 16666 29996 16672 30048
rect 16724 29996 16730 30048
rect 16758 29996 16764 30048
rect 16816 30036 16822 30048
rect 16853 30039 16911 30045
rect 16853 30036 16865 30039
rect 16816 30008 16865 30036
rect 16816 29996 16822 30008
rect 16853 30005 16865 30008
rect 16899 30005 16911 30039
rect 16853 29999 16911 30005
rect 19242 29996 19248 30048
rect 19300 30036 19306 30048
rect 19889 30039 19947 30045
rect 19889 30036 19901 30039
rect 19300 30008 19901 30036
rect 19300 29996 19306 30008
rect 19889 30005 19901 30008
rect 19935 30005 19947 30039
rect 19889 29999 19947 30005
rect 20346 29996 20352 30048
rect 20404 30036 20410 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 20404 30008 22017 30036
rect 20404 29996 20410 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 22005 29999 22063 30005
rect 23750 29996 23756 30048
rect 23808 30036 23814 30048
rect 25774 30036 25780 30048
rect 23808 30008 25780 30036
rect 23808 29996 23814 30008
rect 25774 29996 25780 30008
rect 25832 29996 25838 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 12066 29792 12072 29844
rect 12124 29832 12130 29844
rect 13449 29835 13507 29841
rect 12124 29804 12940 29832
rect 12124 29792 12130 29804
rect 12912 29773 12940 29804
rect 13449 29801 13461 29835
rect 13495 29832 13507 29835
rect 13814 29832 13820 29844
rect 13495 29804 13820 29832
rect 13495 29801 13507 29804
rect 13449 29795 13507 29801
rect 13814 29792 13820 29804
rect 13872 29792 13878 29844
rect 16301 29835 16359 29841
rect 16301 29801 16313 29835
rect 16347 29832 16359 29835
rect 16347 29804 18368 29832
rect 16347 29801 16359 29804
rect 16301 29795 16359 29801
rect 12897 29767 12955 29773
rect 12897 29733 12909 29767
rect 12943 29764 12955 29767
rect 12943 29736 15884 29764
rect 12943 29733 12955 29736
rect 12897 29727 12955 29733
rect 11149 29699 11207 29705
rect 11149 29665 11161 29699
rect 11195 29696 11207 29699
rect 11422 29696 11428 29708
rect 11195 29668 11428 29696
rect 11195 29665 11207 29668
rect 11149 29659 11207 29665
rect 11422 29656 11428 29668
rect 11480 29696 11486 29708
rect 13354 29696 13360 29708
rect 11480 29668 13360 29696
rect 11480 29656 11486 29668
rect 13354 29656 13360 29668
rect 13412 29656 13418 29708
rect 15856 29705 15884 29736
rect 15841 29699 15899 29705
rect 15841 29665 15853 29699
rect 15887 29696 15899 29699
rect 16022 29696 16028 29708
rect 15887 29668 16028 29696
rect 15887 29665 15899 29668
rect 15841 29659 15899 29665
rect 16022 29656 16028 29668
rect 16080 29656 16086 29708
rect 15286 29588 15292 29640
rect 15344 29628 15350 29640
rect 15565 29631 15623 29637
rect 15565 29628 15577 29631
rect 15344 29600 15577 29628
rect 15344 29588 15350 29600
rect 15565 29597 15577 29600
rect 15611 29628 15623 29631
rect 16316 29628 16344 29795
rect 16482 29724 16488 29776
rect 16540 29724 16546 29776
rect 18340 29764 18368 29804
rect 18690 29792 18696 29844
rect 18748 29832 18754 29844
rect 18785 29835 18843 29841
rect 18785 29832 18797 29835
rect 18748 29804 18797 29832
rect 18748 29792 18754 29804
rect 18785 29801 18797 29804
rect 18831 29801 18843 29835
rect 18785 29795 18843 29801
rect 22830 29792 22836 29844
rect 22888 29832 22894 29844
rect 25133 29835 25191 29841
rect 25133 29832 25145 29835
rect 22888 29804 25145 29832
rect 22888 29792 22894 29804
rect 25133 29801 25145 29804
rect 25179 29801 25191 29835
rect 25133 29795 25191 29801
rect 23750 29764 23756 29776
rect 18340 29736 23756 29764
rect 23750 29724 23756 29736
rect 23808 29724 23814 29776
rect 23845 29767 23903 29773
rect 23845 29733 23857 29767
rect 23891 29764 23903 29767
rect 25682 29764 25688 29776
rect 23891 29736 25688 29764
rect 23891 29733 23903 29736
rect 23845 29727 23903 29733
rect 25682 29724 25688 29736
rect 25740 29724 25746 29776
rect 17037 29699 17095 29705
rect 17037 29665 17049 29699
rect 17083 29696 17095 29699
rect 19334 29696 19340 29708
rect 17083 29668 19340 29696
rect 17083 29665 17095 29668
rect 17037 29659 17095 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 20717 29699 20775 29705
rect 20717 29696 20729 29699
rect 19444 29668 20729 29696
rect 15611 29600 16344 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 18414 29588 18420 29640
rect 18472 29588 18478 29640
rect 18874 29628 18880 29640
rect 18616 29600 18880 29628
rect 11146 29520 11152 29572
rect 11204 29560 11210 29572
rect 11425 29563 11483 29569
rect 11425 29560 11437 29563
rect 11204 29532 11437 29560
rect 11204 29520 11210 29532
rect 11425 29529 11437 29532
rect 11471 29529 11483 29563
rect 12710 29560 12716 29572
rect 12650 29532 12716 29560
rect 11425 29523 11483 29529
rect 12710 29520 12716 29532
rect 12768 29520 12774 29572
rect 15657 29563 15715 29569
rect 15657 29529 15669 29563
rect 15703 29560 15715 29563
rect 16482 29560 16488 29572
rect 15703 29532 16488 29560
rect 15703 29529 15715 29532
rect 15657 29523 15715 29529
rect 16482 29520 16488 29532
rect 16540 29520 16546 29572
rect 17313 29563 17371 29569
rect 17313 29529 17325 29563
rect 17359 29529 17371 29563
rect 17313 29523 17371 29529
rect 12728 29492 12756 29520
rect 13265 29495 13323 29501
rect 13265 29492 13277 29495
rect 12728 29464 13277 29492
rect 13265 29461 13277 29464
rect 13311 29492 13323 29495
rect 13725 29495 13783 29501
rect 13725 29492 13737 29495
rect 13311 29464 13737 29492
rect 13311 29461 13323 29464
rect 13265 29455 13323 29461
rect 13725 29461 13737 29464
rect 13771 29492 13783 29495
rect 15010 29492 15016 29504
rect 13771 29464 15016 29492
rect 13771 29461 13783 29464
rect 13725 29455 13783 29461
rect 15010 29452 15016 29464
rect 15068 29452 15074 29504
rect 15194 29452 15200 29504
rect 15252 29452 15258 29504
rect 17328 29492 17356 29523
rect 18616 29492 18644 29600
rect 18874 29588 18880 29600
rect 18932 29628 18938 29640
rect 19444 29628 19472 29668
rect 20717 29665 20729 29668
rect 20763 29665 20775 29699
rect 24854 29696 24860 29708
rect 20717 29659 20775 29665
rect 22066 29668 24860 29696
rect 18932 29600 19472 29628
rect 20625 29631 20683 29637
rect 18932 29588 18938 29600
rect 20625 29597 20637 29631
rect 20671 29628 20683 29631
rect 22066 29628 22094 29668
rect 24854 29656 24860 29668
rect 24912 29656 24918 29708
rect 20671 29600 22094 29628
rect 23385 29631 23443 29637
rect 20671 29597 20683 29600
rect 20625 29591 20683 29597
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29628 24087 29631
rect 24578 29628 24584 29640
rect 24075 29600 24584 29628
rect 24075 29597 24087 29600
rect 24029 29591 24087 29597
rect 22925 29563 22983 29569
rect 22925 29529 22937 29563
rect 22971 29560 22983 29563
rect 23400 29560 23428 29591
rect 24578 29588 24584 29600
rect 24636 29588 24642 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 24854 29560 24860 29572
rect 22971 29532 24860 29560
rect 22971 29529 22983 29532
rect 22925 29523 22983 29529
rect 24854 29520 24860 29532
rect 24912 29520 24918 29572
rect 17328 29464 18644 29492
rect 19150 29452 19156 29504
rect 19208 29492 19214 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 19208 29464 19441 29492
rect 19208 29452 19214 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19429 29455 19487 29461
rect 19610 29452 19616 29504
rect 19668 29492 19674 29504
rect 20165 29495 20223 29501
rect 20165 29492 20177 29495
rect 19668 29464 20177 29492
rect 19668 29452 19674 29464
rect 20165 29461 20177 29464
rect 20211 29461 20223 29495
rect 20165 29455 20223 29461
rect 20530 29452 20536 29504
rect 20588 29452 20594 29504
rect 22462 29452 22468 29504
rect 22520 29492 22526 29504
rect 23201 29495 23259 29501
rect 23201 29492 23213 29495
rect 22520 29464 23213 29492
rect 22520 29452 22526 29464
rect 23201 29461 23213 29464
rect 23247 29461 23259 29495
rect 23201 29455 23259 29461
rect 24489 29495 24547 29501
rect 24489 29461 24501 29495
rect 24535 29492 24547 29495
rect 24578 29492 24584 29504
rect 24535 29464 24584 29492
rect 24535 29461 24547 29464
rect 24489 29455 24547 29461
rect 24578 29452 24584 29464
rect 24636 29452 24642 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 8846 29248 8852 29300
rect 8904 29288 8910 29300
rect 9493 29291 9551 29297
rect 9493 29288 9505 29291
rect 8904 29260 9505 29288
rect 8904 29248 8910 29260
rect 9493 29257 9505 29260
rect 9539 29257 9551 29291
rect 9493 29251 9551 29257
rect 12434 29248 12440 29300
rect 12492 29288 12498 29300
rect 12529 29291 12587 29297
rect 12529 29288 12541 29291
rect 12492 29260 12541 29288
rect 12492 29248 12498 29260
rect 12529 29257 12541 29260
rect 12575 29257 12587 29291
rect 12529 29251 12587 29257
rect 12618 29248 12624 29300
rect 12676 29248 12682 29300
rect 13814 29248 13820 29300
rect 13872 29248 13878 29300
rect 13906 29248 13912 29300
rect 13964 29288 13970 29300
rect 15105 29291 15163 29297
rect 15105 29288 15117 29291
rect 13964 29260 15117 29288
rect 13964 29248 13970 29260
rect 15105 29257 15117 29260
rect 15151 29257 15163 29291
rect 15105 29251 15163 29257
rect 9861 29223 9919 29229
rect 9861 29189 9873 29223
rect 9907 29220 9919 29223
rect 10410 29220 10416 29232
rect 9907 29192 10416 29220
rect 9907 29189 9919 29192
rect 9861 29183 9919 29189
rect 10410 29180 10416 29192
rect 10468 29180 10474 29232
rect 13832 29220 13860 29248
rect 15010 29220 15016 29232
rect 13280 29192 13860 29220
rect 14858 29192 15016 29220
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29152 10011 29155
rect 10226 29152 10232 29164
rect 9999 29124 10232 29152
rect 9999 29121 10011 29124
rect 9953 29115 10011 29121
rect 10226 29112 10232 29124
rect 10284 29112 10290 29164
rect 10042 29044 10048 29096
rect 10100 29044 10106 29096
rect 11606 29044 11612 29096
rect 11664 29084 11670 29096
rect 12805 29087 12863 29093
rect 12805 29084 12817 29087
rect 11664 29056 12817 29084
rect 11664 29044 11670 29056
rect 12805 29053 12817 29056
rect 12851 29084 12863 29087
rect 13280 29084 13308 29192
rect 15010 29180 15016 29192
rect 15068 29180 15074 29232
rect 13354 29112 13360 29164
rect 13412 29112 13418 29164
rect 15120 29152 15148 29251
rect 15194 29248 15200 29300
rect 15252 29288 15258 29300
rect 16025 29291 16083 29297
rect 16025 29288 16037 29291
rect 15252 29260 16037 29288
rect 15252 29248 15258 29260
rect 16025 29257 16037 29260
rect 16071 29257 16083 29291
rect 16025 29251 16083 29257
rect 16206 29248 16212 29300
rect 16264 29288 16270 29300
rect 18785 29291 18843 29297
rect 18785 29288 18797 29291
rect 16264 29260 18797 29288
rect 16264 29248 16270 29260
rect 18785 29257 18797 29260
rect 18831 29257 18843 29291
rect 18785 29251 18843 29257
rect 19150 29248 19156 29300
rect 19208 29248 19214 29300
rect 20530 29248 20536 29300
rect 20588 29288 20594 29300
rect 23842 29288 23848 29300
rect 20588 29260 23848 29288
rect 20588 29248 20594 29260
rect 23842 29248 23848 29260
rect 23900 29288 23906 29300
rect 23937 29291 23995 29297
rect 23937 29288 23949 29291
rect 23900 29260 23949 29288
rect 23900 29248 23906 29260
rect 23937 29257 23949 29260
rect 23983 29257 23995 29291
rect 23937 29251 23995 29257
rect 25314 29248 25320 29300
rect 25372 29288 25378 29300
rect 25409 29291 25467 29297
rect 25409 29288 25421 29291
rect 25372 29260 25421 29288
rect 25372 29248 25378 29260
rect 25409 29257 25421 29260
rect 25455 29257 25467 29291
rect 25409 29251 25467 29257
rect 15930 29180 15936 29232
rect 15988 29180 15994 29232
rect 17144 29192 17448 29220
rect 17144 29152 17172 29192
rect 15120 29124 17172 29152
rect 17218 29112 17224 29164
rect 17276 29112 17282 29164
rect 17310 29112 17316 29164
rect 17368 29112 17374 29164
rect 12851 29056 13308 29084
rect 12851 29053 12863 29056
rect 12805 29047 12863 29053
rect 13630 29044 13636 29096
rect 13688 29084 13694 29096
rect 16117 29087 16175 29093
rect 16117 29084 16129 29087
rect 13688 29056 16129 29084
rect 13688 29044 13694 29056
rect 16117 29053 16129 29056
rect 16163 29053 16175 29087
rect 16117 29047 16175 29053
rect 12161 29019 12219 29025
rect 12161 28985 12173 29019
rect 12207 29016 12219 29019
rect 12250 29016 12256 29028
rect 12207 28988 12256 29016
rect 12207 28985 12219 28988
rect 12161 28979 12219 28985
rect 12250 28976 12256 28988
rect 12308 28976 12314 29028
rect 15194 28976 15200 29028
rect 15252 29016 15258 29028
rect 15565 29019 15623 29025
rect 15565 29016 15577 29019
rect 15252 28988 15577 29016
rect 15252 28976 15258 28988
rect 15565 28985 15577 28988
rect 15611 28985 15623 29019
rect 15565 28979 15623 28985
rect 16574 28976 16580 29028
rect 16632 29016 16638 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 16632 28988 16865 29016
rect 16632 28976 16638 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 17236 29016 17264 29112
rect 17420 29096 17448 29192
rect 19058 29180 19064 29232
rect 19116 29220 19122 29232
rect 19245 29223 19303 29229
rect 19245 29220 19257 29223
rect 19116 29192 19257 29220
rect 19116 29180 19122 29192
rect 19245 29189 19257 29192
rect 19291 29189 19303 29223
rect 19245 29183 19303 29189
rect 17494 29112 17500 29164
rect 17552 29152 17558 29164
rect 17865 29155 17923 29161
rect 17865 29152 17877 29155
rect 17552 29124 17877 29152
rect 17552 29112 17558 29124
rect 17865 29121 17877 29124
rect 17911 29121 17923 29155
rect 17865 29115 17923 29121
rect 18414 29112 18420 29164
rect 18472 29152 18478 29164
rect 20441 29155 20499 29161
rect 20441 29152 20453 29155
rect 18472 29124 20453 29152
rect 18472 29112 18478 29124
rect 20441 29121 20453 29124
rect 20487 29121 20499 29155
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 20441 29115 20499 29121
rect 22066 29124 22201 29152
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 19429 29087 19487 29093
rect 19429 29053 19441 29087
rect 19475 29084 19487 29087
rect 20898 29084 20904 29096
rect 19475 29056 20904 29084
rect 19475 29053 19487 29056
rect 19429 29047 19487 29053
rect 20898 29044 20904 29056
rect 20956 29044 20962 29096
rect 17494 29016 17500 29028
rect 17236 28988 17500 29016
rect 16853 28979 16911 28985
rect 17494 28976 17500 28988
rect 17552 29016 17558 29028
rect 18049 29019 18107 29025
rect 18049 29016 18061 29019
rect 17552 28988 18061 29016
rect 17552 28976 17558 28988
rect 18049 28985 18061 28988
rect 18095 28985 18107 29019
rect 18049 28979 18107 28985
rect 19518 28976 19524 29028
rect 19576 29016 19582 29028
rect 19981 29019 20039 29025
rect 19981 29016 19993 29019
rect 19576 28988 19993 29016
rect 19576 28976 19582 28988
rect 19981 28985 19993 28988
rect 20027 29016 20039 29019
rect 20530 29016 20536 29028
rect 20027 28988 20536 29016
rect 20027 28985 20039 28988
rect 19981 28979 20039 28985
rect 20530 28976 20536 28988
rect 20588 28976 20594 29028
rect 21818 28976 21824 29028
rect 21876 29016 21882 29028
rect 22066 29016 22094 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 24029 29155 24087 29161
rect 24029 29121 24041 29155
rect 24075 29152 24087 29155
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 24075 29124 25329 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 25317 29121 25329 29124
rect 25363 29152 25375 29155
rect 26510 29152 26516 29164
rect 25363 29124 26516 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 26510 29112 26516 29124
rect 26568 29112 26574 29164
rect 23017 29087 23075 29093
rect 23017 29053 23029 29087
rect 23063 29084 23075 29087
rect 23382 29084 23388 29096
rect 23063 29056 23388 29084
rect 23063 29053 23075 29056
rect 23017 29047 23075 29053
rect 23382 29044 23388 29056
rect 23440 29044 23446 29096
rect 23750 29044 23756 29096
rect 23808 29084 23814 29096
rect 24121 29087 24179 29093
rect 24121 29084 24133 29087
rect 23808 29056 24133 29084
rect 23808 29044 23814 29056
rect 24121 29053 24133 29056
rect 24167 29053 24179 29087
rect 24121 29047 24179 29053
rect 24765 29087 24823 29093
rect 24765 29053 24777 29087
rect 24811 29084 24823 29087
rect 24946 29084 24952 29096
rect 24811 29056 24952 29084
rect 24811 29053 24823 29056
rect 24765 29047 24823 29053
rect 24946 29044 24952 29056
rect 25004 29044 25010 29096
rect 21876 28988 22094 29016
rect 23569 29019 23627 29025
rect 21876 28976 21882 28988
rect 23569 28985 23581 29019
rect 23615 29016 23627 29019
rect 23615 28988 24164 29016
rect 23615 28985 23627 28988
rect 23569 28979 23627 28985
rect 24136 28960 24164 28988
rect 13620 28951 13678 28957
rect 13620 28917 13632 28951
rect 13666 28948 13678 28951
rect 14090 28948 14096 28960
rect 13666 28920 14096 28948
rect 13666 28917 13678 28920
rect 13620 28911 13678 28917
rect 14090 28908 14096 28920
rect 14148 28908 14154 28960
rect 15010 28908 15016 28960
rect 15068 28948 15074 28960
rect 15930 28948 15936 28960
rect 15068 28920 15936 28948
rect 15068 28908 15074 28920
rect 15930 28908 15936 28920
rect 15988 28948 15994 28960
rect 18414 28948 18420 28960
rect 15988 28920 18420 28948
rect 15988 28908 15994 28920
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 24118 28908 24124 28960
rect 24176 28908 24182 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 10042 28704 10048 28756
rect 10100 28744 10106 28756
rect 10873 28747 10931 28753
rect 10873 28744 10885 28747
rect 10100 28716 10885 28744
rect 10100 28704 10106 28716
rect 10873 28713 10885 28716
rect 10919 28713 10931 28747
rect 10873 28707 10931 28713
rect 12066 28704 12072 28756
rect 12124 28744 12130 28756
rect 14550 28744 14556 28756
rect 12124 28716 14556 28744
rect 12124 28704 12130 28716
rect 14550 28704 14556 28716
rect 14608 28704 14614 28756
rect 16301 28747 16359 28753
rect 16301 28744 16313 28747
rect 15304 28716 16313 28744
rect 9125 28611 9183 28617
rect 9125 28577 9137 28611
rect 9171 28608 9183 28611
rect 11422 28608 11428 28620
rect 9171 28580 11428 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 13173 28611 13231 28617
rect 13173 28577 13185 28611
rect 13219 28608 13231 28611
rect 14090 28608 14096 28620
rect 13219 28580 14096 28608
rect 13219 28577 13231 28580
rect 13173 28571 13231 28577
rect 14090 28568 14096 28580
rect 14148 28568 14154 28620
rect 15304 28617 15332 28716
rect 16301 28713 16313 28716
rect 16347 28744 16359 28747
rect 16482 28744 16488 28756
rect 16347 28716 16488 28744
rect 16347 28713 16359 28716
rect 16301 28707 16359 28713
rect 16482 28704 16488 28716
rect 16540 28744 16546 28756
rect 18598 28744 18604 28756
rect 16540 28716 18604 28744
rect 16540 28704 16546 28716
rect 18598 28704 18604 28716
rect 18656 28704 18662 28756
rect 18874 28704 18880 28756
rect 18932 28704 18938 28756
rect 22373 28747 22431 28753
rect 22373 28713 22385 28747
rect 22419 28744 22431 28747
rect 23750 28744 23756 28756
rect 22419 28716 23756 28744
rect 22419 28713 22431 28716
rect 22373 28707 22431 28713
rect 23750 28704 23756 28716
rect 23808 28704 23814 28756
rect 15930 28636 15936 28688
rect 15988 28636 15994 28688
rect 21910 28636 21916 28688
rect 21968 28676 21974 28688
rect 22833 28679 22891 28685
rect 22833 28676 22845 28679
rect 21968 28648 22845 28676
rect 21968 28636 21974 28648
rect 22833 28645 22845 28648
rect 22879 28645 22891 28679
rect 22833 28639 22891 28645
rect 23198 28636 23204 28688
rect 23256 28676 23262 28688
rect 24029 28679 24087 28685
rect 24029 28676 24041 28679
rect 23256 28648 24041 28676
rect 23256 28636 23262 28648
rect 24029 28645 24041 28648
rect 24075 28645 24087 28679
rect 24029 28639 24087 28645
rect 15289 28611 15347 28617
rect 15289 28577 15301 28611
rect 15335 28577 15347 28611
rect 15289 28571 15347 28577
rect 15378 28568 15384 28620
rect 15436 28568 15442 28620
rect 17405 28611 17463 28617
rect 17405 28577 17417 28611
rect 17451 28608 17463 28611
rect 18966 28608 18972 28620
rect 17451 28580 18972 28608
rect 17451 28577 17463 28580
rect 17405 28571 17463 28577
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 20073 28611 20131 28617
rect 20073 28577 20085 28611
rect 20119 28608 20131 28611
rect 20990 28608 20996 28620
rect 20119 28580 20996 28608
rect 20119 28577 20131 28580
rect 20073 28571 20131 28577
rect 20990 28568 20996 28580
rect 21048 28568 21054 28620
rect 23385 28611 23443 28617
rect 23385 28577 23397 28611
rect 23431 28608 23443 28611
rect 23658 28608 23664 28620
rect 23431 28580 23664 28608
rect 23431 28577 23443 28580
rect 23385 28571 23443 28577
rect 23658 28568 23664 28580
rect 23716 28568 23722 28620
rect 24854 28568 24860 28620
rect 24912 28608 24918 28620
rect 25041 28611 25099 28617
rect 25041 28608 25053 28611
rect 24912 28580 25053 28608
rect 24912 28568 24918 28580
rect 25041 28577 25053 28580
rect 25087 28577 25099 28611
rect 25041 28571 25099 28577
rect 25225 28611 25283 28617
rect 25225 28577 25237 28611
rect 25271 28608 25283 28611
rect 25406 28608 25412 28620
rect 25271 28580 25412 28608
rect 25271 28577 25283 28580
rect 25225 28571 25283 28577
rect 25406 28568 25412 28580
rect 25464 28568 25470 28620
rect 15102 28500 15108 28552
rect 15160 28540 15166 28552
rect 17129 28543 17187 28549
rect 17129 28540 17141 28543
rect 15160 28512 17141 28540
rect 15160 28500 15166 28512
rect 17129 28509 17141 28512
rect 17175 28509 17187 28543
rect 17129 28503 17187 28509
rect 18414 28500 18420 28552
rect 18472 28540 18478 28552
rect 18472 28512 18538 28540
rect 18472 28500 18478 28512
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 20622 28540 20628 28552
rect 19392 28512 20628 28540
rect 19392 28500 19398 28512
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 23293 28543 23351 28549
rect 23293 28509 23305 28543
rect 23339 28540 23351 28543
rect 23566 28540 23572 28552
rect 23339 28512 23572 28540
rect 23339 28509 23351 28512
rect 23293 28503 23351 28509
rect 23566 28500 23572 28512
rect 23624 28500 23630 28552
rect 24946 28500 24952 28552
rect 25004 28500 25010 28552
rect 9401 28475 9459 28481
rect 9401 28441 9413 28475
rect 9447 28472 9459 28475
rect 9674 28472 9680 28484
rect 9447 28444 9680 28472
rect 9447 28441 9459 28444
rect 9401 28435 9459 28441
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 10962 28472 10968 28484
rect 10626 28444 10968 28472
rect 10962 28432 10968 28444
rect 11020 28432 11026 28484
rect 11701 28475 11759 28481
rect 11701 28472 11713 28475
rect 11532 28444 11713 28472
rect 11532 28416 11560 28444
rect 11701 28441 11713 28444
rect 11747 28441 11759 28475
rect 15197 28475 15255 28481
rect 12926 28444 13584 28472
rect 11701 28435 11759 28441
rect 13556 28416 13584 28444
rect 15197 28441 15209 28475
rect 15243 28441 15255 28475
rect 15197 28435 15255 28441
rect 19889 28475 19947 28481
rect 19889 28441 19901 28475
rect 19935 28472 19947 28475
rect 20806 28472 20812 28484
rect 19935 28444 20812 28472
rect 19935 28441 19947 28444
rect 19889 28435 19947 28441
rect 11514 28364 11520 28416
rect 11572 28364 11578 28416
rect 13538 28364 13544 28416
rect 13596 28364 13602 28416
rect 14826 28364 14832 28416
rect 14884 28364 14890 28416
rect 15212 28404 15240 28435
rect 20806 28432 20812 28444
rect 20864 28432 20870 28484
rect 20898 28432 20904 28484
rect 20956 28432 20962 28484
rect 22126 28444 23980 28472
rect 23952 28416 23980 28444
rect 16022 28404 16028 28416
rect 15212 28376 16028 28404
rect 16022 28364 16028 28376
rect 16080 28364 16086 28416
rect 19429 28407 19487 28413
rect 19429 28373 19441 28407
rect 19475 28404 19487 28407
rect 19518 28404 19524 28416
rect 19475 28376 19524 28404
rect 19475 28373 19487 28376
rect 19429 28367 19487 28373
rect 19518 28364 19524 28376
rect 19576 28364 19582 28416
rect 19702 28364 19708 28416
rect 19760 28404 19766 28416
rect 19797 28407 19855 28413
rect 19797 28404 19809 28407
rect 19760 28376 19809 28404
rect 19760 28364 19766 28376
rect 19797 28373 19809 28376
rect 19843 28373 19855 28407
rect 19797 28367 19855 28373
rect 22278 28364 22284 28416
rect 22336 28404 22342 28416
rect 23198 28404 23204 28416
rect 22336 28376 23204 28404
rect 22336 28364 22342 28376
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 23934 28364 23940 28416
rect 23992 28364 23998 28416
rect 24394 28364 24400 28416
rect 24452 28404 24458 28416
rect 24581 28407 24639 28413
rect 24581 28404 24593 28407
rect 24452 28376 24593 28404
rect 24452 28364 24458 28376
rect 24581 28373 24593 28376
rect 24627 28373 24639 28407
rect 24581 28367 24639 28373
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 13538 28160 13544 28212
rect 13596 28200 13602 28212
rect 13817 28203 13875 28209
rect 13817 28200 13829 28203
rect 13596 28172 13829 28200
rect 13596 28160 13602 28172
rect 13817 28169 13829 28172
rect 13863 28200 13875 28203
rect 15010 28200 15016 28212
rect 13863 28172 15016 28200
rect 13863 28169 13875 28172
rect 13817 28163 13875 28169
rect 15010 28160 15016 28172
rect 15068 28160 15074 28212
rect 15565 28203 15623 28209
rect 15565 28169 15577 28203
rect 15611 28200 15623 28203
rect 15838 28200 15844 28212
rect 15611 28172 15844 28200
rect 15611 28169 15623 28172
rect 15565 28163 15623 28169
rect 15838 28160 15844 28172
rect 15896 28200 15902 28212
rect 16393 28203 16451 28209
rect 16393 28200 16405 28203
rect 15896 28172 16405 28200
rect 15896 28160 15902 28172
rect 16393 28169 16405 28172
rect 16439 28169 16451 28203
rect 16393 28163 16451 28169
rect 17126 28160 17132 28212
rect 17184 28200 17190 28212
rect 17221 28203 17279 28209
rect 17221 28200 17233 28203
rect 17184 28172 17233 28200
rect 17184 28160 17190 28172
rect 17221 28169 17233 28172
rect 17267 28169 17279 28203
rect 17221 28163 17279 28169
rect 11054 28092 11060 28144
rect 11112 28132 11118 28144
rect 11977 28135 12035 28141
rect 11977 28132 11989 28135
rect 11112 28104 11989 28132
rect 11112 28092 11118 28104
rect 11977 28101 11989 28104
rect 12023 28101 12035 28135
rect 13556 28132 13584 28160
rect 13202 28118 13584 28132
rect 11977 28095 12035 28101
rect 13188 28104 13584 28118
rect 17236 28132 17264 28163
rect 18506 28160 18512 28212
rect 18564 28200 18570 28212
rect 18782 28200 18788 28212
rect 18564 28172 18788 28200
rect 18564 28160 18570 28172
rect 18782 28160 18788 28172
rect 18840 28200 18846 28212
rect 18969 28203 19027 28209
rect 18969 28200 18981 28203
rect 18840 28172 18981 28200
rect 18840 28160 18846 28172
rect 18969 28169 18981 28172
rect 19015 28169 19027 28203
rect 18969 28163 19027 28169
rect 19702 28160 19708 28212
rect 19760 28160 19766 28212
rect 22465 28203 22523 28209
rect 22465 28169 22477 28203
rect 22511 28200 22523 28203
rect 24210 28200 24216 28212
rect 22511 28172 24216 28200
rect 22511 28169 22523 28172
rect 22465 28163 22523 28169
rect 24210 28160 24216 28172
rect 24268 28160 24274 28212
rect 18693 28135 18751 28141
rect 18693 28132 18705 28135
rect 17236 28104 18705 28132
rect 11698 27956 11704 28008
rect 11756 27956 11762 28008
rect 12618 27956 12624 28008
rect 12676 27996 12682 28008
rect 13188 27996 13216 28104
rect 18432 28076 18460 28104
rect 18693 28101 18705 28104
rect 18739 28101 18751 28135
rect 18693 28095 18751 28101
rect 20622 28092 20628 28144
rect 20680 28132 20686 28144
rect 21085 28135 21143 28141
rect 21085 28132 21097 28135
rect 20680 28104 21097 28132
rect 20680 28092 20686 28104
rect 21085 28101 21097 28104
rect 21131 28101 21143 28135
rect 21085 28095 21143 28101
rect 22554 28092 22560 28144
rect 22612 28092 22618 28144
rect 23382 28132 23388 28144
rect 23216 28104 23388 28132
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28064 15715 28067
rect 16298 28064 16304 28076
rect 15703 28036 16304 28064
rect 15703 28033 15715 28036
rect 15657 28027 15715 28033
rect 16298 28024 16304 28036
rect 16356 28024 16362 28076
rect 18414 28024 18420 28076
rect 18472 28024 18478 28076
rect 20349 28067 20407 28073
rect 20349 28033 20361 28067
rect 20395 28064 20407 28067
rect 21818 28064 21824 28076
rect 20395 28036 21824 28064
rect 20395 28033 20407 28036
rect 20349 28027 20407 28033
rect 12676 27968 13216 27996
rect 15749 27999 15807 28005
rect 12676 27956 12682 27968
rect 15749 27965 15761 27999
rect 15795 27965 15807 27999
rect 15749 27959 15807 27965
rect 17313 27999 17371 28005
rect 17313 27965 17325 27999
rect 17359 27965 17371 27999
rect 17313 27959 17371 27965
rect 10778 27888 10784 27940
rect 10836 27928 10842 27940
rect 15378 27928 15384 27940
rect 10836 27900 11652 27928
rect 10836 27888 10842 27900
rect 10962 27820 10968 27872
rect 11020 27820 11026 27872
rect 11624 27860 11652 27900
rect 13464 27900 15384 27928
rect 13464 27869 13492 27900
rect 15378 27888 15384 27900
rect 15436 27928 15442 27940
rect 15764 27928 15792 27959
rect 15436 27900 15792 27928
rect 15436 27888 15442 27900
rect 13449 27863 13507 27869
rect 13449 27860 13461 27863
rect 11624 27832 13461 27860
rect 13449 27829 13461 27832
rect 13495 27829 13507 27863
rect 13449 27823 13507 27829
rect 13814 27820 13820 27872
rect 13872 27860 13878 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 13872 27832 15209 27860
rect 13872 27820 13878 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 16298 27820 16304 27872
rect 16356 27820 16362 27872
rect 16850 27820 16856 27872
rect 16908 27820 16914 27872
rect 17328 27860 17356 27959
rect 17402 27956 17408 28008
rect 17460 27956 17466 28008
rect 18049 27999 18107 28005
rect 18049 27965 18061 27999
rect 18095 27996 18107 27999
rect 18138 27996 18144 28008
rect 18095 27968 18144 27996
rect 18095 27965 18107 27968
rect 18049 27959 18107 27965
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 17678 27888 17684 27940
rect 17736 27928 17742 27940
rect 19337 27931 19395 27937
rect 19337 27928 19349 27931
rect 17736 27900 19349 27928
rect 17736 27888 17742 27900
rect 19337 27897 19349 27900
rect 19383 27928 19395 27931
rect 20364 27928 20392 28027
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28064 22431 28067
rect 22572 28064 22600 28092
rect 23216 28073 23244 28104
rect 23382 28092 23388 28104
rect 23440 28092 23446 28144
rect 23474 28092 23480 28144
rect 23532 28092 23538 28144
rect 23934 28092 23940 28144
rect 23992 28092 23998 28144
rect 23201 28067 23259 28073
rect 22419 28036 23152 28064
rect 22419 28033 22431 28036
rect 22373 28027 22431 28033
rect 19383 27900 20392 27928
rect 19383 27897 19395 27900
rect 19337 27891 19395 27897
rect 20530 27888 20536 27940
rect 20588 27928 20594 27940
rect 22005 27931 22063 27937
rect 22005 27928 22017 27931
rect 20588 27900 22017 27928
rect 20588 27888 20594 27900
rect 22005 27897 22017 27900
rect 22051 27897 22063 27931
rect 22388 27928 22416 28027
rect 22554 27956 22560 28008
rect 22612 27956 22618 28008
rect 23124 27996 23152 28036
rect 23201 28033 23213 28067
rect 23247 28033 23259 28067
rect 23201 28027 23259 28033
rect 23124 27968 25544 27996
rect 22005 27891 22063 27897
rect 22296 27900 22416 27928
rect 17586 27860 17592 27872
rect 17328 27832 17592 27860
rect 17586 27820 17592 27832
rect 17644 27860 17650 27872
rect 18506 27860 18512 27872
rect 17644 27832 18512 27860
rect 17644 27820 17650 27832
rect 18506 27820 18512 27832
rect 18564 27820 18570 27872
rect 20990 27820 20996 27872
rect 21048 27860 21054 27872
rect 21545 27863 21603 27869
rect 21545 27860 21557 27863
rect 21048 27832 21557 27860
rect 21048 27820 21054 27832
rect 21545 27829 21557 27832
rect 21591 27860 21603 27863
rect 22296 27860 22324 27900
rect 21591 27832 22324 27860
rect 21591 27829 21603 27832
rect 21545 27823 21603 27829
rect 22370 27820 22376 27872
rect 22428 27860 22434 27872
rect 23290 27860 23296 27872
rect 22428 27832 23296 27860
rect 22428 27820 22434 27832
rect 23290 27820 23296 27832
rect 23348 27860 23354 27872
rect 24949 27863 25007 27869
rect 24949 27860 24961 27863
rect 23348 27832 24961 27860
rect 23348 27820 23354 27832
rect 24949 27829 24961 27832
rect 24995 27829 25007 27863
rect 24949 27823 25007 27829
rect 25222 27820 25228 27872
rect 25280 27820 25286 27872
rect 25516 27869 25544 27968
rect 25501 27863 25559 27869
rect 25501 27829 25513 27863
rect 25547 27860 25559 27863
rect 25958 27860 25964 27872
rect 25547 27832 25964 27860
rect 25547 27829 25559 27832
rect 25501 27823 25559 27829
rect 25958 27820 25964 27832
rect 26016 27820 26022 27872
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 11422 27656 11428 27668
rect 10612 27628 11428 27656
rect 9030 27548 9036 27600
rect 9088 27588 9094 27600
rect 9125 27591 9183 27597
rect 9125 27588 9137 27591
rect 9088 27560 9137 27588
rect 9088 27548 9094 27560
rect 9125 27557 9137 27560
rect 9171 27557 9183 27591
rect 9125 27551 9183 27557
rect 3418 27480 3424 27532
rect 3476 27520 3482 27532
rect 7653 27523 7711 27529
rect 7653 27520 7665 27523
rect 3476 27492 7665 27520
rect 3476 27480 3482 27492
rect 7653 27489 7665 27492
rect 7699 27520 7711 27523
rect 10505 27523 10563 27529
rect 7699 27492 10456 27520
rect 7699 27489 7711 27492
rect 7653 27483 7711 27489
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27452 7435 27455
rect 7423 27424 9076 27452
rect 7423 27421 7435 27424
rect 7377 27415 7435 27421
rect 9048 27393 9076 27424
rect 9033 27387 9091 27393
rect 9033 27353 9045 27387
rect 9079 27384 9091 27387
rect 10428 27384 10456 27492
rect 10505 27489 10517 27523
rect 10551 27520 10563 27523
rect 10612 27520 10640 27628
rect 11422 27616 11428 27628
rect 11480 27616 11486 27668
rect 12618 27616 12624 27668
rect 12676 27616 12682 27668
rect 15102 27656 15108 27668
rect 13188 27628 15108 27656
rect 11790 27548 11796 27600
rect 11848 27588 11854 27600
rect 13078 27588 13084 27600
rect 11848 27560 13084 27588
rect 11848 27548 11854 27560
rect 13078 27548 13084 27560
rect 13136 27588 13142 27600
rect 13188 27588 13216 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 16482 27616 16488 27668
rect 16540 27616 16546 27668
rect 19978 27616 19984 27668
rect 20036 27616 20042 27668
rect 20152 27659 20210 27665
rect 20152 27625 20164 27659
rect 20198 27656 20210 27659
rect 23658 27656 23664 27668
rect 20198 27628 23664 27656
rect 20198 27625 20210 27628
rect 20152 27619 20210 27625
rect 23658 27616 23664 27628
rect 23716 27656 23722 27668
rect 23845 27659 23903 27665
rect 23845 27656 23857 27659
rect 23716 27628 23857 27656
rect 23716 27616 23722 27628
rect 23845 27625 23857 27628
rect 23891 27625 23903 27659
rect 23845 27619 23903 27625
rect 13136 27560 13216 27588
rect 13136 27548 13142 27560
rect 19426 27548 19432 27600
rect 19484 27588 19490 27600
rect 19996 27588 20024 27616
rect 19484 27560 20024 27588
rect 19484 27548 19490 27560
rect 23474 27548 23480 27600
rect 23532 27588 23538 27600
rect 24762 27588 24768 27600
rect 23532 27560 24768 27588
rect 23532 27548 23538 27560
rect 24762 27548 24768 27560
rect 24820 27588 24826 27600
rect 24820 27560 25176 27588
rect 24820 27548 24826 27560
rect 10551 27492 10640 27520
rect 10551 27489 10563 27492
rect 10505 27483 10563 27489
rect 10778 27480 10784 27532
rect 10836 27480 10842 27532
rect 10870 27480 10876 27532
rect 10928 27520 10934 27532
rect 11974 27520 11980 27532
rect 10928 27492 11980 27520
rect 10928 27480 10934 27492
rect 11974 27480 11980 27492
rect 12032 27480 12038 27532
rect 13354 27480 13360 27532
rect 13412 27520 13418 27532
rect 13541 27523 13599 27529
rect 13541 27520 13553 27523
rect 13412 27492 13553 27520
rect 13412 27480 13418 27492
rect 13541 27489 13553 27492
rect 13587 27489 13599 27523
rect 13541 27483 13599 27489
rect 14734 27480 14740 27532
rect 14792 27520 14798 27532
rect 15749 27523 15807 27529
rect 15749 27520 15761 27523
rect 14792 27492 15761 27520
rect 14792 27480 14798 27492
rect 15749 27489 15761 27492
rect 15795 27489 15807 27523
rect 15749 27483 15807 27489
rect 17770 27480 17776 27532
rect 17828 27520 17834 27532
rect 18049 27523 18107 27529
rect 18049 27520 18061 27523
rect 17828 27492 18061 27520
rect 17828 27480 17834 27492
rect 18049 27489 18061 27492
rect 18095 27489 18107 27523
rect 18049 27483 18107 27489
rect 19889 27523 19947 27529
rect 19889 27489 19901 27523
rect 19935 27520 19947 27523
rect 22097 27523 22155 27529
rect 22097 27520 22109 27523
rect 19935 27492 22109 27520
rect 19935 27489 19947 27492
rect 19889 27483 19947 27489
rect 22097 27489 22109 27492
rect 22143 27520 22155 27523
rect 23382 27520 23388 27532
rect 22143 27492 23388 27520
rect 22143 27489 22155 27492
rect 22097 27483 22155 27489
rect 23382 27480 23388 27492
rect 23440 27480 23446 27532
rect 23842 27480 23848 27532
rect 23900 27520 23906 27532
rect 24121 27523 24179 27529
rect 24121 27520 24133 27523
rect 23900 27492 24133 27520
rect 23900 27480 23906 27492
rect 24121 27489 24133 27492
rect 24167 27489 24179 27523
rect 24121 27483 24179 27489
rect 25038 27480 25044 27532
rect 25096 27480 25102 27532
rect 25148 27529 25176 27560
rect 25133 27523 25191 27529
rect 25133 27489 25145 27523
rect 25179 27489 25191 27523
rect 25133 27483 25191 27489
rect 11882 27412 11888 27464
rect 11940 27452 11946 27464
rect 12618 27452 12624 27464
rect 11940 27424 12624 27452
rect 11940 27412 11946 27424
rect 12618 27412 12624 27424
rect 12676 27412 12682 27464
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 14826 27452 14832 27464
rect 13495 27424 14832 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 15657 27455 15715 27461
rect 15657 27421 15669 27455
rect 15703 27452 15715 27455
rect 16482 27452 16488 27464
rect 15703 27424 16488 27452
rect 15703 27421 15715 27424
rect 15657 27415 15715 27421
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 18138 27452 18144 27464
rect 17911 27424 18144 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 18138 27412 18144 27424
rect 18196 27412 18202 27464
rect 23934 27452 23940 27464
rect 23506 27424 23940 27452
rect 23934 27412 23940 27424
rect 23992 27412 23998 27464
rect 10870 27384 10876 27396
rect 9079 27356 9536 27384
rect 10428 27356 10876 27384
rect 9079 27353 9091 27356
rect 9033 27347 9091 27353
rect 9508 27316 9536 27356
rect 10870 27344 10876 27356
rect 10928 27344 10934 27396
rect 13357 27387 13415 27393
rect 13357 27353 13369 27387
rect 13403 27384 13415 27387
rect 13814 27384 13820 27396
rect 13403 27356 13820 27384
rect 13403 27353 13415 27356
rect 13357 27347 13415 27353
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 16022 27384 16028 27396
rect 15580 27356 16028 27384
rect 15580 27328 15608 27356
rect 16022 27344 16028 27356
rect 16080 27384 16086 27396
rect 16209 27387 16267 27393
rect 16209 27384 16221 27387
rect 16080 27356 16221 27384
rect 16080 27344 16086 27356
rect 16209 27353 16221 27356
rect 16255 27353 16267 27387
rect 17957 27387 18015 27393
rect 16209 27347 16267 27353
rect 16408 27356 17908 27384
rect 12066 27316 12072 27328
rect 9508 27288 12072 27316
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 12158 27276 12164 27328
rect 12216 27316 12222 27328
rect 12253 27319 12311 27325
rect 12253 27316 12265 27319
rect 12216 27288 12265 27316
rect 12216 27276 12222 27288
rect 12253 27285 12265 27288
rect 12299 27285 12311 27319
rect 12253 27279 12311 27285
rect 12618 27276 12624 27328
rect 12676 27316 12682 27328
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 12676 27288 13001 27316
rect 12676 27276 12682 27288
rect 12989 27285 13001 27288
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13722 27276 13728 27328
rect 13780 27316 13786 27328
rect 15197 27319 15255 27325
rect 15197 27316 15209 27319
rect 13780 27288 15209 27316
rect 13780 27276 13786 27288
rect 15197 27285 15209 27288
rect 15243 27285 15255 27319
rect 15197 27279 15255 27285
rect 15562 27276 15568 27328
rect 15620 27276 15626 27328
rect 15654 27276 15660 27328
rect 15712 27316 15718 27328
rect 16408 27316 16436 27356
rect 15712 27288 16436 27316
rect 15712 27276 15718 27288
rect 16482 27276 16488 27328
rect 16540 27316 16546 27328
rect 17497 27319 17555 27325
rect 17497 27316 17509 27319
rect 16540 27288 17509 27316
rect 16540 27276 16546 27288
rect 17497 27285 17509 27288
rect 17543 27285 17555 27319
rect 17880 27316 17908 27356
rect 17957 27353 17969 27387
rect 18003 27384 18015 27387
rect 19886 27384 19892 27396
rect 18003 27356 19892 27384
rect 18003 27353 18015 27356
rect 17957 27347 18015 27353
rect 19886 27344 19892 27356
rect 19944 27344 19950 27396
rect 20088 27356 20654 27384
rect 20088 27328 20116 27356
rect 22370 27344 22376 27396
rect 22428 27344 22434 27396
rect 23658 27344 23664 27396
rect 23716 27384 23722 27396
rect 23716 27356 24624 27384
rect 23716 27344 23722 27356
rect 19426 27316 19432 27328
rect 17880 27288 19432 27316
rect 17497 27279 17555 27285
rect 19426 27276 19432 27288
rect 19484 27276 19490 27328
rect 19613 27319 19671 27325
rect 19613 27285 19625 27319
rect 19659 27316 19671 27319
rect 20070 27316 20076 27328
rect 19659 27288 20076 27316
rect 19659 27285 19671 27288
rect 19613 27279 19671 27285
rect 20070 27276 20076 27288
rect 20128 27276 20134 27328
rect 21634 27276 21640 27328
rect 21692 27276 21698 27328
rect 24596 27325 24624 27356
rect 24581 27319 24639 27325
rect 24581 27285 24593 27319
rect 24627 27285 24639 27319
rect 24581 27279 24639 27285
rect 24949 27319 25007 27325
rect 24949 27285 24961 27319
rect 24995 27316 25007 27319
rect 25038 27316 25044 27328
rect 24995 27288 25044 27316
rect 24995 27285 25007 27288
rect 24949 27279 25007 27285
rect 25038 27276 25044 27288
rect 25096 27316 25102 27328
rect 25222 27316 25228 27328
rect 25096 27288 25228 27316
rect 25096 27276 25102 27288
rect 25222 27276 25228 27288
rect 25280 27276 25286 27328
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 9766 27112 9772 27124
rect 9324 27084 9772 27112
rect 7653 26979 7711 26985
rect 7653 26945 7665 26979
rect 7699 26976 7711 26979
rect 9030 26976 9036 26988
rect 7699 26948 9036 26976
rect 7699 26945 7711 26948
rect 7653 26939 7711 26945
rect 9030 26936 9036 26948
rect 9088 26936 9094 26988
rect 9324 26985 9352 27084
rect 9766 27072 9772 27084
rect 9824 27112 9830 27124
rect 10870 27112 10876 27124
rect 9824 27084 10876 27112
rect 9824 27072 9830 27084
rect 10870 27072 10876 27084
rect 10928 27112 10934 27124
rect 11790 27112 11796 27124
rect 10928 27084 11796 27112
rect 10928 27072 10934 27084
rect 11790 27072 11796 27084
rect 11848 27072 11854 27124
rect 11974 27072 11980 27124
rect 12032 27112 12038 27124
rect 15562 27112 15568 27124
rect 12032 27084 15568 27112
rect 12032 27072 12038 27084
rect 15562 27072 15568 27084
rect 15620 27072 15626 27124
rect 15657 27115 15715 27121
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16850 27112 16856 27124
rect 15703 27084 16856 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 19242 27112 19248 27124
rect 18064 27084 19248 27112
rect 10962 27044 10968 27056
rect 10810 27016 10968 27044
rect 10962 27004 10968 27016
rect 11020 27044 11026 27056
rect 11609 27047 11667 27053
rect 11609 27044 11621 27047
rect 11020 27016 11621 27044
rect 11020 27004 11026 27016
rect 11609 27013 11621 27016
rect 11655 27044 11667 27047
rect 11882 27044 11888 27056
rect 11655 27016 11888 27044
rect 11655 27013 11667 27016
rect 11609 27007 11667 27013
rect 11882 27004 11888 27016
rect 11940 27004 11946 27056
rect 13262 27044 13268 27056
rect 12176 27016 13268 27044
rect 12176 26988 12204 27016
rect 13262 27004 13268 27016
rect 13320 27004 13326 27056
rect 13357 27047 13415 27053
rect 13357 27013 13369 27047
rect 13403 27044 13415 27047
rect 13630 27044 13636 27056
rect 13403 27016 13636 27044
rect 13403 27013 13415 27016
rect 13357 27007 13415 27013
rect 13630 27004 13636 27016
rect 13688 27004 13694 27056
rect 15749 27047 15807 27053
rect 15749 27013 15761 27047
rect 15795 27044 15807 27047
rect 16574 27044 16580 27056
rect 15795 27016 16580 27044
rect 15795 27013 15807 27016
rect 15749 27007 15807 27013
rect 16574 27004 16580 27016
rect 16632 27004 16638 27056
rect 18064 27044 18092 27084
rect 19242 27072 19248 27084
rect 19300 27072 19306 27124
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 22833 27115 22891 27121
rect 22833 27112 22845 27115
rect 22796 27084 22845 27112
rect 22796 27072 22802 27084
rect 22833 27081 22845 27084
rect 22879 27081 22891 27115
rect 22833 27075 22891 27081
rect 24762 27072 24768 27124
rect 24820 27112 24826 27124
rect 25317 27115 25375 27121
rect 25317 27112 25329 27115
rect 24820 27084 25329 27112
rect 24820 27072 24826 27084
rect 25317 27081 25329 27084
rect 25363 27081 25375 27115
rect 25317 27075 25375 27081
rect 17972 27016 18092 27044
rect 9309 26979 9367 26985
rect 9309 26945 9321 26979
rect 9355 26945 9367 26979
rect 12158 26976 12164 26988
rect 9309 26939 9367 26945
rect 10980 26948 12164 26976
rect 7558 26868 7564 26920
rect 7616 26908 7622 26920
rect 7929 26911 7987 26917
rect 7929 26908 7941 26911
rect 7616 26880 7941 26908
rect 7616 26868 7622 26880
rect 7929 26877 7941 26880
rect 7975 26877 7987 26911
rect 9585 26911 9643 26917
rect 9585 26908 9597 26911
rect 7929 26871 7987 26877
rect 9324 26880 9597 26908
rect 7944 26772 7972 26871
rect 9324 26852 9352 26880
rect 9585 26877 9597 26880
rect 9631 26908 9643 26911
rect 10980 26908 11008 26948
rect 12158 26936 12164 26948
rect 12216 26936 12222 26988
rect 12802 26936 12808 26988
rect 12860 26976 12866 26988
rect 13078 26976 13084 26988
rect 12860 26948 13084 26976
rect 12860 26936 12866 26948
rect 13078 26936 13084 26948
rect 13136 26936 13142 26988
rect 15930 26976 15936 26988
rect 14490 26948 15936 26976
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 17972 26985 18000 27016
rect 18782 27004 18788 27056
rect 18840 27004 18846 27056
rect 23566 27044 23572 27056
rect 23032 27016 23572 27044
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 22646 26936 22652 26988
rect 22704 26976 22710 26988
rect 22741 26979 22799 26985
rect 22741 26976 22753 26979
rect 22704 26948 22753 26976
rect 22704 26936 22710 26948
rect 22741 26945 22753 26948
rect 22787 26945 22799 26979
rect 22741 26939 22799 26945
rect 9631 26880 11008 26908
rect 11057 26911 11115 26917
rect 9631 26877 9643 26880
rect 9585 26871 9643 26877
rect 11057 26877 11069 26911
rect 11103 26908 11115 26911
rect 11146 26908 11152 26920
rect 11103 26880 11152 26908
rect 11103 26877 11115 26880
rect 11057 26871 11115 26877
rect 11146 26868 11152 26880
rect 11204 26868 11210 26920
rect 15746 26908 15752 26920
rect 11256 26880 15752 26908
rect 9306 26800 9312 26852
rect 9364 26800 9370 26852
rect 11256 26772 11284 26880
rect 15746 26868 15752 26880
rect 15804 26868 15810 26920
rect 15841 26911 15899 26917
rect 15841 26877 15853 26911
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 22094 26908 22100 26920
rect 18279 26880 22100 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 15856 26840 15884 26871
rect 22094 26868 22100 26880
rect 22152 26908 22158 26920
rect 22554 26908 22560 26920
rect 22152 26880 22560 26908
rect 22152 26868 22158 26880
rect 22554 26868 22560 26880
rect 22612 26868 22618 26920
rect 23032 26917 23060 27016
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 23934 27004 23940 27056
rect 23992 27044 23998 27056
rect 23992 27016 24334 27044
rect 23992 27004 23998 27016
rect 23017 26911 23075 26917
rect 23017 26877 23029 26911
rect 23063 26877 23075 26911
rect 23017 26871 23075 26877
rect 23382 26868 23388 26920
rect 23440 26908 23446 26920
rect 23569 26911 23627 26917
rect 23569 26908 23581 26911
rect 23440 26880 23581 26908
rect 23440 26868 23446 26880
rect 23569 26877 23581 26880
rect 23615 26877 23627 26911
rect 23569 26871 23627 26877
rect 23845 26911 23903 26917
rect 23845 26877 23857 26911
rect 23891 26908 23903 26911
rect 25222 26908 25228 26920
rect 23891 26880 25228 26908
rect 23891 26877 23903 26880
rect 23845 26871 23903 26877
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 14844 26812 15884 26840
rect 7944 26744 11284 26772
rect 11974 26732 11980 26784
rect 12032 26772 12038 26784
rect 14844 26781 14872 26812
rect 14829 26775 14887 26781
rect 14829 26772 14841 26775
rect 12032 26744 14841 26772
rect 12032 26732 12038 26744
rect 14829 26741 14841 26744
rect 14875 26741 14887 26775
rect 14829 26735 14887 26741
rect 14918 26732 14924 26784
rect 14976 26772 14982 26784
rect 15289 26775 15347 26781
rect 15289 26772 15301 26775
rect 14976 26744 15301 26772
rect 14976 26732 14982 26744
rect 15289 26741 15301 26744
rect 15335 26741 15347 26775
rect 15289 26735 15347 26741
rect 18966 26732 18972 26784
rect 19024 26772 19030 26784
rect 19705 26775 19763 26781
rect 19705 26772 19717 26775
rect 19024 26744 19717 26772
rect 19024 26732 19030 26744
rect 19705 26741 19717 26744
rect 19751 26741 19763 26775
rect 19705 26735 19763 26741
rect 20070 26732 20076 26784
rect 20128 26772 20134 26784
rect 21082 26772 21088 26784
rect 20128 26744 21088 26772
rect 20128 26732 20134 26744
rect 21082 26732 21088 26744
rect 21140 26772 21146 26784
rect 21545 26775 21603 26781
rect 21545 26772 21557 26775
rect 21140 26744 21557 26772
rect 21140 26732 21146 26744
rect 21545 26741 21557 26744
rect 21591 26772 21603 26775
rect 21913 26775 21971 26781
rect 21913 26772 21925 26775
rect 21591 26744 21925 26772
rect 21591 26741 21603 26744
rect 21545 26735 21603 26741
rect 21913 26741 21925 26744
rect 21959 26741 21971 26775
rect 21913 26735 21971 26741
rect 22370 26732 22376 26784
rect 22428 26732 22434 26784
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 9398 26528 9404 26580
rect 9456 26568 9462 26580
rect 11333 26571 11391 26577
rect 11333 26568 11345 26571
rect 9456 26540 11345 26568
rect 9456 26528 9462 26540
rect 11333 26537 11345 26540
rect 11379 26568 11391 26571
rect 11606 26568 11612 26580
rect 11379 26540 11612 26568
rect 11379 26537 11391 26540
rect 11333 26531 11391 26537
rect 11606 26528 11612 26540
rect 11664 26528 11670 26580
rect 15746 26528 15752 26580
rect 15804 26568 15810 26580
rect 20990 26568 20996 26580
rect 15804 26540 20996 26568
rect 15804 26528 15810 26540
rect 20990 26528 20996 26540
rect 21048 26528 21054 26580
rect 21177 26571 21235 26577
rect 21177 26537 21189 26571
rect 21223 26568 21235 26571
rect 22094 26568 22100 26580
rect 21223 26540 22100 26568
rect 21223 26537 21235 26540
rect 21177 26531 21235 26537
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 25038 26568 25044 26580
rect 22480 26540 25044 26568
rect 11241 26503 11299 26509
rect 11241 26469 11253 26503
rect 11287 26500 11299 26503
rect 11882 26500 11888 26512
rect 11287 26472 11888 26500
rect 11287 26469 11299 26472
rect 11241 26463 11299 26469
rect 9125 26435 9183 26441
rect 9125 26401 9137 26435
rect 9171 26432 9183 26435
rect 9766 26432 9772 26444
rect 9171 26404 9772 26432
rect 9171 26401 9183 26404
rect 9125 26395 9183 26401
rect 9766 26392 9772 26404
rect 9824 26392 9830 26444
rect 10873 26435 10931 26441
rect 10873 26401 10885 26435
rect 10919 26432 10931 26435
rect 11054 26432 11060 26444
rect 10919 26404 11060 26432
rect 10919 26401 10931 26404
rect 10873 26395 10931 26401
rect 11054 26392 11060 26404
rect 11112 26392 11118 26444
rect 11256 26364 11284 26463
rect 11882 26460 11888 26472
rect 11940 26500 11946 26512
rect 12710 26500 12716 26512
rect 11940 26472 12716 26500
rect 11940 26460 11946 26472
rect 12710 26460 12716 26472
rect 12768 26460 12774 26512
rect 14274 26460 14280 26512
rect 14332 26500 14338 26512
rect 15657 26503 15715 26509
rect 15657 26500 15669 26503
rect 14332 26472 15669 26500
rect 14332 26460 14338 26472
rect 15657 26469 15669 26472
rect 15703 26469 15715 26503
rect 15657 26463 15715 26469
rect 16022 26460 16028 26512
rect 16080 26500 16086 26512
rect 16758 26500 16764 26512
rect 16080 26472 16764 26500
rect 16080 26460 16086 26472
rect 16758 26460 16764 26472
rect 16816 26500 16822 26512
rect 16816 26472 16896 26500
rect 16816 26460 16822 26472
rect 14826 26392 14832 26444
rect 14884 26392 14890 26444
rect 15381 26435 15439 26441
rect 15381 26401 15393 26435
rect 15427 26432 15439 26435
rect 15470 26432 15476 26444
rect 15427 26404 15476 26432
rect 15427 26401 15439 26404
rect 15381 26395 15439 26401
rect 15470 26392 15476 26404
rect 15528 26432 15534 26444
rect 15930 26432 15936 26444
rect 15528 26404 15936 26432
rect 15528 26392 15534 26404
rect 15930 26392 15936 26404
rect 15988 26392 15994 26444
rect 16209 26435 16267 26441
rect 16209 26401 16221 26435
rect 16255 26401 16267 26435
rect 16209 26395 16267 26401
rect 11330 26364 11336 26376
rect 10534 26336 11336 26364
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 14734 26324 14740 26376
rect 14792 26364 14798 26376
rect 16224 26364 16252 26395
rect 14792 26336 16252 26364
rect 14792 26324 14798 26336
rect 16666 26324 16672 26376
rect 16724 26324 16730 26376
rect 16868 26373 16896 26472
rect 18782 26460 18788 26512
rect 18840 26500 18846 26512
rect 18969 26503 19027 26509
rect 18969 26500 18981 26503
rect 18840 26472 18981 26500
rect 18840 26460 18846 26472
rect 18969 26469 18981 26472
rect 19015 26469 19027 26503
rect 18969 26463 19027 26469
rect 22002 26460 22008 26512
rect 22060 26500 22066 26512
rect 22480 26500 22508 26540
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 22060 26472 22508 26500
rect 22060 26460 22066 26472
rect 22554 26460 22560 26512
rect 22612 26500 22618 26512
rect 22649 26503 22707 26509
rect 22649 26500 22661 26503
rect 22612 26472 22661 26500
rect 22612 26460 22618 26472
rect 22649 26469 22661 26472
rect 22695 26469 22707 26503
rect 22649 26463 22707 26469
rect 23845 26503 23903 26509
rect 23845 26469 23857 26503
rect 23891 26469 23903 26503
rect 23845 26463 23903 26469
rect 24581 26503 24639 26509
rect 24581 26469 24593 26503
rect 24627 26500 24639 26503
rect 24854 26500 24860 26512
rect 24627 26472 24860 26500
rect 24627 26469 24639 26472
rect 24581 26463 24639 26469
rect 19426 26392 19432 26444
rect 19484 26392 19490 26444
rect 19705 26435 19763 26441
rect 19705 26401 19717 26435
rect 19751 26432 19763 26435
rect 20990 26432 20996 26444
rect 19751 26404 20996 26432
rect 19751 26401 19763 26404
rect 19705 26395 19763 26401
rect 20990 26392 20996 26404
rect 21048 26432 21054 26444
rect 21634 26432 21640 26444
rect 21048 26404 21640 26432
rect 21048 26392 21054 26404
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 22186 26392 22192 26444
rect 22244 26432 22250 26444
rect 23201 26435 23259 26441
rect 23201 26432 23213 26435
rect 22244 26404 23213 26432
rect 22244 26392 22250 26404
rect 23201 26401 23213 26404
rect 23247 26401 23259 26435
rect 23860 26432 23888 26463
rect 24854 26460 24860 26472
rect 24912 26460 24918 26512
rect 23860 26404 24992 26432
rect 23201 26395 23259 26401
rect 16853 26367 16911 26373
rect 16853 26333 16865 26367
rect 16899 26364 16911 26367
rect 17862 26364 17868 26376
rect 16899 26336 17868 26364
rect 16899 26333 16911 26336
rect 16853 26327 16911 26333
rect 17862 26324 17868 26336
rect 17920 26324 17926 26376
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26364 22155 26367
rect 24026 26364 24032 26376
rect 22143 26336 24032 26364
rect 22143 26333 22155 26336
rect 22097 26327 22155 26333
rect 24026 26324 24032 26336
rect 24084 26324 24090 26376
rect 24964 26364 24992 26404
rect 25038 26392 25044 26444
rect 25096 26432 25102 26444
rect 25133 26435 25191 26441
rect 25133 26432 25145 26435
rect 25096 26404 25145 26432
rect 25096 26392 25102 26404
rect 25133 26401 25145 26404
rect 25179 26401 25191 26435
rect 25133 26395 25191 26401
rect 25498 26364 25504 26376
rect 24964 26336 25504 26364
rect 25498 26324 25504 26336
rect 25556 26324 25562 26376
rect 8938 26256 8944 26308
rect 8996 26296 9002 26308
rect 9398 26296 9404 26308
rect 8996 26268 9404 26296
rect 8996 26256 9002 26268
rect 9398 26256 9404 26268
rect 9456 26256 9462 26308
rect 14645 26299 14703 26305
rect 14645 26265 14657 26299
rect 14691 26296 14703 26299
rect 15930 26296 15936 26308
rect 14691 26268 15936 26296
rect 14691 26265 14703 26268
rect 14645 26259 14703 26265
rect 15930 26256 15936 26268
rect 15988 26256 15994 26308
rect 16117 26299 16175 26305
rect 16117 26265 16129 26299
rect 16163 26296 16175 26299
rect 16298 26296 16304 26308
rect 16163 26268 16304 26296
rect 16163 26265 16175 26268
rect 16117 26259 16175 26265
rect 16298 26256 16304 26268
rect 16356 26296 16362 26308
rect 16942 26296 16948 26308
rect 16356 26268 16948 26296
rect 16356 26256 16362 26268
rect 16942 26256 16948 26268
rect 17000 26296 17006 26308
rect 17037 26299 17095 26305
rect 17037 26296 17049 26299
rect 17000 26268 17049 26296
rect 17000 26256 17006 26268
rect 17037 26265 17049 26268
rect 17083 26265 17095 26299
rect 21082 26296 21088 26308
rect 20930 26268 21088 26296
rect 17037 26259 17095 26265
rect 21082 26256 21088 26268
rect 21140 26256 21146 26308
rect 22373 26299 22431 26305
rect 22373 26265 22385 26299
rect 22419 26265 22431 26299
rect 22373 26259 22431 26265
rect 14277 26231 14335 26237
rect 14277 26197 14289 26231
rect 14323 26228 14335 26231
rect 14458 26228 14464 26240
rect 14323 26200 14464 26228
rect 14323 26197 14335 26200
rect 14277 26191 14335 26197
rect 14458 26188 14464 26200
rect 14516 26188 14522 26240
rect 14737 26231 14795 26237
rect 14737 26197 14749 26231
rect 14783 26228 14795 26231
rect 15010 26228 15016 26240
rect 14783 26200 15016 26228
rect 14783 26197 14795 26200
rect 14737 26191 14795 26197
rect 15010 26188 15016 26200
rect 15068 26188 15074 26240
rect 15838 26188 15844 26240
rect 15896 26228 15902 26240
rect 16025 26231 16083 26237
rect 16025 26228 16037 26231
rect 15896 26200 16037 26228
rect 15896 26188 15902 26200
rect 16025 26197 16037 26200
rect 16071 26228 16083 26231
rect 17218 26228 17224 26240
rect 16071 26200 17224 26228
rect 16071 26197 16083 26200
rect 16025 26191 16083 26197
rect 17218 26188 17224 26200
rect 17276 26188 17282 26240
rect 18233 26231 18291 26237
rect 18233 26197 18245 26231
rect 18279 26228 18291 26231
rect 18322 26228 18328 26240
rect 18279 26200 18328 26228
rect 18279 26197 18291 26200
rect 18233 26191 18291 26197
rect 18322 26188 18328 26200
rect 18380 26188 18386 26240
rect 22278 26188 22284 26240
rect 22336 26228 22342 26240
rect 22388 26228 22416 26259
rect 22830 26256 22836 26308
rect 22888 26296 22894 26308
rect 23109 26299 23167 26305
rect 23109 26296 23121 26299
rect 22888 26268 23121 26296
rect 22888 26256 22894 26268
rect 23109 26265 23121 26268
rect 23155 26265 23167 26299
rect 23109 26259 23167 26265
rect 24949 26299 25007 26305
rect 24949 26265 24961 26299
rect 24995 26265 25007 26299
rect 24949 26259 25007 26265
rect 25041 26299 25099 26305
rect 25041 26265 25053 26299
rect 25087 26296 25099 26299
rect 25130 26296 25136 26308
rect 25087 26268 25136 26296
rect 25087 26265 25099 26268
rect 25041 26259 25099 26265
rect 23014 26228 23020 26240
rect 22336 26200 23020 26228
rect 22336 26188 22342 26200
rect 23014 26188 23020 26200
rect 23072 26188 23078 26240
rect 24964 26228 24992 26259
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 25958 26296 25964 26308
rect 25240 26268 25964 26296
rect 25240 26228 25268 26268
rect 25958 26256 25964 26268
rect 26016 26256 26022 26308
rect 24964 26200 25268 26228
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 9490 25984 9496 26036
rect 9548 25984 9554 26036
rect 12161 26027 12219 26033
rect 12161 25993 12173 26027
rect 12207 26024 12219 26027
rect 12207 25996 12434 26024
rect 12207 25993 12219 25996
rect 12161 25987 12219 25993
rect 8021 25891 8079 25897
rect 8021 25857 8033 25891
rect 8067 25888 8079 25891
rect 9508 25888 9536 25984
rect 12406 25956 12434 25996
rect 12618 25984 12624 26036
rect 12676 25984 12682 26036
rect 13832 25996 16252 26024
rect 13832 25956 13860 25996
rect 12406 25928 13860 25956
rect 13906 25916 13912 25968
rect 13964 25916 13970 25968
rect 14001 25959 14059 25965
rect 14001 25925 14013 25959
rect 14047 25956 14059 25959
rect 15102 25956 15108 25968
rect 14047 25928 15108 25956
rect 14047 25925 14059 25928
rect 14001 25919 14059 25925
rect 15102 25916 15108 25928
rect 15160 25916 15166 25968
rect 16224 25956 16252 25996
rect 16850 25984 16856 26036
rect 16908 25984 16914 26036
rect 17034 25984 17040 26036
rect 17092 26024 17098 26036
rect 17773 26027 17831 26033
rect 17773 26024 17785 26027
rect 17092 25996 17785 26024
rect 17092 25984 17098 25996
rect 17773 25993 17785 25996
rect 17819 25993 17831 26027
rect 17773 25987 17831 25993
rect 18141 26027 18199 26033
rect 18141 25993 18153 26027
rect 18187 26024 18199 26027
rect 18322 26024 18328 26036
rect 18187 25996 18328 26024
rect 18187 25993 18199 25996
rect 18141 25987 18199 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 18598 25984 18604 26036
rect 18656 26024 18662 26036
rect 19061 26027 19119 26033
rect 19061 26024 19073 26027
rect 18656 25996 19073 26024
rect 18656 25984 18662 25996
rect 19061 25993 19073 25996
rect 19107 25993 19119 26027
rect 22278 26024 22284 26036
rect 19061 25987 19119 25993
rect 19720 25996 22284 26024
rect 18233 25959 18291 25965
rect 16224 25928 17080 25956
rect 8067 25860 9536 25888
rect 12529 25891 12587 25897
rect 8067 25857 8079 25860
rect 8021 25851 8079 25857
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 12618 25888 12624 25900
rect 12575 25860 12624 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 12618 25848 12624 25860
rect 12676 25848 12682 25900
rect 17052 25897 17080 25928
rect 18233 25925 18245 25959
rect 18279 25956 18291 25959
rect 19610 25956 19616 25968
rect 18279 25928 19616 25956
rect 18279 25925 18291 25928
rect 18233 25919 18291 25925
rect 19610 25916 19616 25928
rect 19668 25916 19674 25968
rect 15197 25891 15255 25897
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 16025 25891 16083 25897
rect 16025 25888 16037 25891
rect 15243 25860 16037 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 16025 25857 16037 25860
rect 16071 25857 16083 25891
rect 16025 25851 16083 25857
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 17126 25848 17132 25900
rect 17184 25888 17190 25900
rect 19720 25888 19748 25996
rect 22278 25984 22284 25996
rect 22336 25984 22342 26036
rect 22462 25984 22468 26036
rect 22520 25984 22526 26036
rect 23014 25984 23020 26036
rect 23072 26024 23078 26036
rect 24946 26024 24952 26036
rect 23072 25996 24952 26024
rect 23072 25984 23078 25996
rect 24946 25984 24952 25996
rect 25004 25984 25010 26036
rect 26234 25956 26240 25968
rect 17184 25860 19748 25888
rect 19812 25928 26240 25956
rect 17184 25848 17190 25860
rect 4798 25780 4804 25832
rect 4856 25820 4862 25832
rect 8297 25823 8355 25829
rect 8297 25820 8309 25823
rect 4856 25792 8309 25820
rect 4856 25780 4862 25792
rect 8297 25789 8309 25792
rect 8343 25789 8355 25823
rect 8297 25783 8355 25789
rect 8312 25752 8340 25783
rect 11146 25780 11152 25832
rect 11204 25820 11210 25832
rect 12713 25823 12771 25829
rect 12713 25820 12725 25823
rect 11204 25792 12725 25820
rect 11204 25780 11210 25792
rect 12713 25789 12725 25792
rect 12759 25789 12771 25823
rect 12713 25783 12771 25789
rect 14090 25780 14096 25832
rect 14148 25780 14154 25832
rect 15289 25823 15347 25829
rect 15289 25820 15301 25823
rect 15212 25792 15301 25820
rect 13446 25752 13452 25764
rect 8312 25724 13452 25752
rect 13446 25712 13452 25724
rect 13504 25712 13510 25764
rect 11790 25644 11796 25696
rect 11848 25684 11854 25696
rect 12434 25684 12440 25696
rect 11848 25656 12440 25684
rect 11848 25644 11854 25656
rect 12434 25644 12440 25656
rect 12492 25644 12498 25696
rect 13538 25644 13544 25696
rect 13596 25644 13602 25696
rect 13814 25644 13820 25696
rect 13872 25684 13878 25696
rect 14829 25687 14887 25693
rect 14829 25684 14841 25687
rect 13872 25656 14841 25684
rect 13872 25644 13878 25656
rect 14829 25653 14841 25656
rect 14875 25653 14887 25687
rect 15212 25684 15240 25792
rect 15289 25789 15301 25792
rect 15335 25789 15347 25823
rect 15289 25783 15347 25789
rect 15378 25780 15384 25832
rect 15436 25780 15442 25832
rect 18417 25823 18475 25829
rect 18417 25789 18429 25823
rect 18463 25820 18475 25823
rect 18690 25820 18696 25832
rect 18463 25792 18696 25820
rect 18463 25789 18475 25792
rect 18417 25783 18475 25789
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 19812 25752 19840 25928
rect 26234 25916 26240 25928
rect 26292 25916 26298 25968
rect 22373 25891 22431 25897
rect 22373 25857 22385 25891
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 22002 25820 22008 25832
rect 17420 25724 19840 25752
rect 21560 25792 22008 25820
rect 17420 25696 17448 25724
rect 21560 25696 21588 25792
rect 22002 25780 22008 25792
rect 22060 25820 22066 25832
rect 22388 25820 22416 25851
rect 23474 25848 23480 25900
rect 23532 25848 23538 25900
rect 23937 25891 23995 25897
rect 23937 25857 23949 25891
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 22060 25792 22416 25820
rect 22649 25823 22707 25829
rect 22060 25780 22066 25792
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 22738 25820 22744 25832
rect 22695 25792 22744 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 22738 25780 22744 25792
rect 22796 25780 22802 25832
rect 22830 25780 22836 25832
rect 22888 25820 22894 25832
rect 23952 25820 23980 25851
rect 22888 25792 23980 25820
rect 22888 25780 22894 25792
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 17402 25684 17408 25696
rect 15212 25656 17408 25684
rect 14829 25647 14887 25653
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 21542 25644 21548 25696
rect 21600 25644 21606 25696
rect 21634 25644 21640 25696
rect 21692 25684 21698 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21692 25656 22017 25684
rect 21692 25644 21698 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 22094 25644 22100 25696
rect 22152 25684 22158 25696
rect 23293 25687 23351 25693
rect 23293 25684 23305 25687
rect 22152 25656 23305 25684
rect 22152 25644 22158 25656
rect 23293 25653 23305 25656
rect 23339 25653 23351 25687
rect 23293 25647 23351 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 11698 25440 11704 25492
rect 11756 25480 11762 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 11756 25452 14289 25480
rect 11756 25440 11762 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 17589 25483 17647 25489
rect 17589 25449 17601 25483
rect 17635 25480 17647 25483
rect 17954 25480 17960 25492
rect 17635 25452 17960 25480
rect 17635 25449 17647 25452
rect 17589 25443 17647 25449
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 18325 25483 18383 25489
rect 18325 25449 18337 25483
rect 18371 25480 18383 25483
rect 18598 25480 18604 25492
rect 18371 25452 18604 25480
rect 18371 25449 18383 25452
rect 18325 25443 18383 25449
rect 18598 25440 18604 25452
rect 18656 25440 18662 25492
rect 20349 25483 20407 25489
rect 20349 25449 20361 25483
rect 20395 25480 20407 25483
rect 21082 25480 21088 25492
rect 20395 25452 21088 25480
rect 20395 25449 20407 25452
rect 20349 25443 20407 25449
rect 21082 25440 21088 25452
rect 21140 25440 21146 25492
rect 21545 25483 21603 25489
rect 21545 25449 21557 25483
rect 21591 25480 21603 25483
rect 22830 25480 22836 25492
rect 21591 25452 22836 25480
rect 21591 25449 21603 25452
rect 21545 25443 21603 25449
rect 22830 25440 22836 25452
rect 22888 25440 22894 25492
rect 23474 25440 23480 25492
rect 23532 25480 23538 25492
rect 25317 25483 25375 25489
rect 25317 25480 25329 25483
rect 23532 25452 25329 25480
rect 23532 25440 23538 25452
rect 25317 25449 25329 25452
rect 25363 25449 25375 25483
rect 25317 25443 25375 25449
rect 12434 25372 12440 25424
rect 12492 25412 12498 25424
rect 15289 25415 15347 25421
rect 15289 25412 15301 25415
rect 12492 25384 15301 25412
rect 12492 25372 12498 25384
rect 15289 25381 15301 25384
rect 15335 25412 15347 25415
rect 15378 25412 15384 25424
rect 15335 25384 15384 25412
rect 15335 25381 15347 25384
rect 15289 25375 15347 25381
rect 15378 25372 15384 25384
rect 15436 25372 15442 25424
rect 16945 25415 17003 25421
rect 16945 25381 16957 25415
rect 16991 25412 17003 25415
rect 16991 25384 21772 25412
rect 16991 25381 17003 25384
rect 16945 25375 17003 25381
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 11149 25347 11207 25353
rect 11149 25313 11161 25347
rect 11195 25344 11207 25347
rect 14734 25344 14740 25356
rect 11195 25316 14740 25344
rect 11195 25313 11207 25316
rect 11149 25307 11207 25313
rect 14734 25304 14740 25316
rect 14792 25304 14798 25356
rect 14826 25304 14832 25356
rect 14884 25304 14890 25356
rect 16301 25347 16359 25353
rect 16301 25344 16313 25347
rect 14936 25316 16313 25344
rect 12710 25276 12716 25288
rect 12282 25248 12716 25276
rect 12710 25236 12716 25248
rect 12768 25276 12774 25288
rect 12897 25279 12955 25285
rect 12897 25276 12909 25279
rect 12768 25248 12909 25276
rect 12768 25236 12774 25248
rect 12897 25245 12909 25248
rect 12943 25245 12955 25279
rect 12897 25239 12955 25245
rect 13354 25236 13360 25288
rect 13412 25276 13418 25288
rect 14936 25276 14964 25316
rect 16301 25313 16313 25316
rect 16347 25313 16359 25347
rect 16301 25307 16359 25313
rect 16850 25304 16856 25356
rect 16908 25344 16914 25356
rect 16908 25316 21036 25344
rect 16908 25304 16914 25316
rect 13412 25248 14964 25276
rect 13412 25236 13418 25248
rect 15194 25236 15200 25288
rect 15252 25276 15258 25288
rect 17129 25279 17187 25285
rect 17129 25276 17141 25279
rect 15252 25248 17141 25276
rect 15252 25236 15258 25248
rect 17129 25245 17141 25248
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 17586 25236 17592 25288
rect 17644 25276 17650 25288
rect 17773 25279 17831 25285
rect 17773 25276 17785 25279
rect 17644 25248 17785 25276
rect 17644 25236 17650 25248
rect 17773 25245 17785 25248
rect 17819 25245 17831 25279
rect 17773 25239 17831 25245
rect 18141 25279 18199 25285
rect 18141 25245 18153 25279
rect 18187 25276 18199 25279
rect 18414 25276 18420 25288
rect 18187 25248 18420 25276
rect 18187 25245 18199 25248
rect 18141 25239 18199 25245
rect 18414 25236 18420 25248
rect 18472 25276 18478 25288
rect 18472 25248 19380 25276
rect 18472 25236 18478 25248
rect 14645 25211 14703 25217
rect 14645 25177 14657 25211
rect 14691 25208 14703 25211
rect 15286 25208 15292 25220
rect 14691 25180 15292 25208
rect 14691 25177 14703 25180
rect 14645 25171 14703 25177
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 16209 25211 16267 25217
rect 16209 25177 16221 25211
rect 16255 25208 16267 25211
rect 18598 25208 18604 25220
rect 16255 25180 18604 25208
rect 16255 25177 16267 25180
rect 16209 25171 16267 25177
rect 18598 25168 18604 25180
rect 18656 25168 18662 25220
rect 19352 25217 19380 25248
rect 19794 25236 19800 25288
rect 19852 25276 19858 25288
rect 21008 25285 21036 25316
rect 21744 25285 21772 25384
rect 20441 25279 20499 25285
rect 20441 25276 20453 25279
rect 19852 25248 20453 25276
rect 19852 25236 19858 25248
rect 20441 25245 20453 25248
rect 20487 25245 20499 25279
rect 20441 25239 20499 25245
rect 20993 25279 21051 25285
rect 20993 25245 21005 25279
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25245 21787 25279
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 21729 25239 21787 25245
rect 22066 25248 22661 25276
rect 19337 25211 19395 25217
rect 19337 25177 19349 25211
rect 19383 25208 19395 25211
rect 20070 25208 20076 25220
rect 19383 25180 20076 25208
rect 19383 25177 19395 25180
rect 19337 25171 19395 25177
rect 20070 25168 20076 25180
rect 20128 25168 20134 25220
rect 22066 25208 22094 25248
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25276 24731 25279
rect 25314 25276 25320 25288
rect 24719 25248 25320 25276
rect 24719 25245 24731 25248
rect 24673 25239 24731 25245
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 20824 25180 22094 25208
rect 12621 25143 12679 25149
rect 12621 25109 12633 25143
rect 12667 25140 12679 25143
rect 12710 25140 12716 25152
rect 12667 25112 12716 25140
rect 12667 25109 12679 25112
rect 12621 25103 12679 25109
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 14737 25143 14795 25149
rect 14737 25109 14749 25143
rect 14783 25140 14795 25143
rect 15378 25140 15384 25152
rect 14783 25112 15384 25140
rect 14783 25109 14795 25112
rect 14737 25103 14795 25109
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 15562 25100 15568 25152
rect 15620 25140 15626 25152
rect 15749 25143 15807 25149
rect 15749 25140 15761 25143
rect 15620 25112 15761 25140
rect 15620 25100 15626 25112
rect 15749 25109 15761 25112
rect 15795 25109 15807 25143
rect 15749 25103 15807 25109
rect 16117 25143 16175 25149
rect 16117 25109 16129 25143
rect 16163 25140 16175 25143
rect 16298 25140 16304 25152
rect 16163 25112 16304 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 16298 25100 16304 25112
rect 16356 25100 16362 25152
rect 18506 25100 18512 25152
rect 18564 25140 18570 25152
rect 18693 25143 18751 25149
rect 18693 25140 18705 25143
rect 18564 25112 18705 25140
rect 18564 25100 18570 25112
rect 18693 25109 18705 25112
rect 18739 25109 18751 25143
rect 18693 25103 18751 25109
rect 19886 25100 19892 25152
rect 19944 25100 19950 25152
rect 20824 25149 20852 25180
rect 23842 25168 23848 25220
rect 23900 25168 23906 25220
rect 20809 25143 20867 25149
rect 20809 25109 20821 25143
rect 20855 25109 20867 25143
rect 20809 25103 20867 25109
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 8312 24908 11008 24936
rect 7282 24760 7288 24812
rect 7340 24800 7346 24812
rect 8312 24800 8340 24908
rect 10134 24828 10140 24880
rect 10192 24828 10198 24880
rect 10980 24868 11008 24908
rect 11238 24896 11244 24948
rect 11296 24936 11302 24948
rect 14826 24936 14832 24948
rect 11296 24908 14832 24936
rect 11296 24896 11302 24908
rect 14826 24896 14832 24908
rect 14884 24896 14890 24948
rect 15105 24939 15163 24945
rect 15105 24905 15117 24939
rect 15151 24936 15163 24939
rect 15286 24936 15292 24948
rect 15151 24908 15292 24936
rect 15151 24905 15163 24908
rect 15105 24899 15163 24905
rect 15286 24896 15292 24908
rect 15344 24896 15350 24948
rect 15470 24896 15476 24948
rect 15528 24896 15534 24948
rect 17218 24896 17224 24948
rect 17276 24896 17282 24948
rect 17862 24896 17868 24948
rect 17920 24936 17926 24948
rect 22278 24936 22284 24948
rect 17920 24908 22284 24936
rect 17920 24896 17926 24908
rect 22278 24896 22284 24908
rect 22336 24896 22342 24948
rect 12069 24871 12127 24877
rect 12069 24868 12081 24871
rect 10980 24840 12081 24868
rect 12069 24837 12081 24840
rect 12115 24837 12127 24871
rect 12069 24831 12127 24837
rect 13538 24828 13544 24880
rect 13596 24868 13602 24880
rect 17236 24868 17264 24896
rect 18322 24868 18328 24880
rect 13596 24840 13754 24868
rect 17236 24840 18328 24868
rect 13596 24828 13602 24840
rect 18322 24828 18328 24840
rect 18380 24868 18386 24880
rect 18380 24840 19104 24868
rect 18380 24828 18386 24840
rect 11146 24800 11152 24812
rect 7340 24772 8340 24800
rect 10980 24772 11152 24800
rect 7340 24760 7346 24772
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24701 9459 24735
rect 9401 24695 9459 24701
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24732 9735 24735
rect 10980 24732 11008 24772
rect 11146 24760 11152 24772
rect 11204 24760 11210 24812
rect 12158 24760 12164 24812
rect 12216 24760 12222 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12860 24772 13001 24800
rect 12860 24760 12866 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 16390 24760 16396 24812
rect 16448 24800 16454 24812
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 16448 24772 17325 24800
rect 16448 24760 16454 24772
rect 17313 24769 17325 24772
rect 17359 24800 17371 24803
rect 17359 24772 18000 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 9723 24704 11008 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 9416 24596 9444 24695
rect 11054 24692 11060 24744
rect 11112 24732 11118 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 11112 24704 12265 24732
rect 11112 24692 11118 24704
rect 12253 24701 12265 24704
rect 12299 24701 12311 24735
rect 12253 24695 12311 24701
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 13906 24732 13912 24744
rect 13311 24704 13912 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 14734 24692 14740 24744
rect 14792 24692 14798 24744
rect 15102 24692 15108 24744
rect 15160 24732 15166 24744
rect 15160 24704 15332 24732
rect 15160 24692 15166 24704
rect 15194 24664 15200 24676
rect 14660 24636 15200 24664
rect 11054 24596 11060 24608
rect 9416 24568 11060 24596
rect 11054 24556 11060 24568
rect 11112 24556 11118 24608
rect 11149 24599 11207 24605
rect 11149 24565 11161 24599
rect 11195 24596 11207 24599
rect 11238 24596 11244 24608
rect 11195 24568 11244 24596
rect 11195 24565 11207 24568
rect 11149 24559 11207 24565
rect 11238 24556 11244 24568
rect 11296 24556 11302 24608
rect 11701 24599 11759 24605
rect 11701 24565 11713 24599
rect 11747 24596 11759 24599
rect 14660 24596 14688 24636
rect 15194 24624 15200 24636
rect 15252 24624 15258 24676
rect 15304 24664 15332 24704
rect 15378 24692 15384 24744
rect 15436 24732 15442 24744
rect 16408 24732 16436 24760
rect 15436 24704 16436 24732
rect 17405 24735 17463 24741
rect 15436 24692 15442 24704
rect 17405 24701 17417 24735
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 17420 24664 17448 24695
rect 15304 24636 17448 24664
rect 17972 24664 18000 24772
rect 18414 24760 18420 24812
rect 18472 24760 18478 24812
rect 18509 24803 18567 24809
rect 18509 24769 18521 24803
rect 18555 24800 18567 24803
rect 18690 24800 18696 24812
rect 18555 24772 18696 24800
rect 18555 24769 18567 24772
rect 18509 24763 18567 24769
rect 18690 24760 18696 24772
rect 18748 24760 18754 24812
rect 19076 24809 19104 24840
rect 22462 24828 22468 24880
rect 22520 24828 22526 24880
rect 23934 24828 23940 24880
rect 23992 24868 23998 24880
rect 23992 24840 24334 24868
rect 23992 24828 23998 24840
rect 19061 24803 19119 24809
rect 19061 24769 19073 24803
rect 19107 24769 19119 24803
rect 19061 24763 19119 24769
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 19484 24772 19717 24800
rect 19484 24760 19490 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 19705 24763 19763 24769
rect 21082 24760 21088 24812
rect 21140 24760 21146 24812
rect 22186 24760 22192 24812
rect 22244 24760 22250 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 23474 24800 23480 24812
rect 22603 24772 23480 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 18598 24692 18604 24744
rect 18656 24692 18662 24744
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 20438 24732 20444 24744
rect 20027 24704 20444 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 20438 24692 20444 24704
rect 20496 24692 20502 24744
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24732 21511 24735
rect 22204 24732 22232 24760
rect 21499 24704 22232 24732
rect 21499 24701 21511 24704
rect 21453 24695 21511 24701
rect 19058 24664 19064 24676
rect 17972 24636 19064 24664
rect 19058 24624 19064 24636
rect 19116 24664 19122 24676
rect 19245 24667 19303 24673
rect 19245 24664 19257 24667
rect 19116 24636 19257 24664
rect 19116 24624 19122 24636
rect 19245 24633 19257 24636
rect 19291 24633 19303 24667
rect 19245 24627 19303 24633
rect 11747 24568 14688 24596
rect 11747 24565 11759 24568
rect 11701 24559 11759 24565
rect 15930 24556 15936 24608
rect 15988 24596 15994 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 15988 24568 16865 24596
rect 15988 24556 15994 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 16853 24559 16911 24565
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17920 24568 18061 24596
rect 17920 24556 17926 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 22097 24599 22155 24605
rect 22097 24596 22109 24599
rect 19392 24568 22109 24596
rect 19392 24556 19398 24568
rect 22097 24565 22109 24568
rect 22143 24565 22155 24599
rect 22204 24596 22232 24704
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24732 22799 24735
rect 23290 24732 23296 24744
rect 22787 24704 23296 24732
rect 22787 24701 22799 24704
rect 22741 24695 22799 24701
rect 23290 24692 23296 24704
rect 23348 24692 23354 24744
rect 23569 24735 23627 24741
rect 23569 24701 23581 24735
rect 23615 24701 23627 24735
rect 23569 24695 23627 24701
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 25038 24732 25044 24744
rect 23891 24704 25044 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 22830 24624 22836 24676
rect 22888 24664 22894 24676
rect 23382 24664 23388 24676
rect 22888 24636 23388 24664
rect 22888 24624 22894 24636
rect 23382 24624 23388 24636
rect 23440 24664 23446 24676
rect 23584 24664 23612 24695
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 25222 24692 25228 24744
rect 25280 24732 25286 24744
rect 25317 24735 25375 24741
rect 25317 24732 25329 24735
rect 25280 24704 25329 24732
rect 25280 24692 25286 24704
rect 25317 24701 25329 24704
rect 25363 24701 25375 24735
rect 25317 24695 25375 24701
rect 23440 24636 23612 24664
rect 23440 24624 23446 24636
rect 22646 24596 22652 24608
rect 22204 24568 22652 24596
rect 22097 24559 22155 24565
rect 22646 24556 22652 24568
rect 22704 24556 22710 24608
rect 23293 24599 23351 24605
rect 23293 24565 23305 24599
rect 23339 24596 23351 24599
rect 23934 24596 23940 24608
rect 23339 24568 23940 24596
rect 23339 24565 23351 24568
rect 23293 24559 23351 24565
rect 23934 24556 23940 24568
rect 23992 24556 23998 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 12710 24392 12716 24404
rect 10428 24364 12716 24392
rect 9401 24259 9459 24265
rect 9401 24225 9413 24259
rect 9447 24256 9459 24259
rect 9490 24256 9496 24268
rect 9447 24228 9496 24256
rect 9447 24225 9459 24228
rect 9401 24219 9459 24225
rect 9490 24216 9496 24228
rect 9548 24256 9554 24268
rect 10428 24256 10456 24364
rect 12710 24352 12716 24364
rect 12768 24392 12774 24404
rect 12894 24392 12900 24404
rect 12768 24364 12900 24392
rect 12768 24352 12774 24364
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 20438 24352 20444 24404
rect 20496 24392 20502 24404
rect 21177 24395 21235 24401
rect 21177 24392 21189 24395
rect 20496 24364 21189 24392
rect 20496 24352 20502 24364
rect 21177 24361 21189 24364
rect 21223 24361 21235 24395
rect 21177 24355 21235 24361
rect 22176 24395 22234 24401
rect 22176 24361 22188 24395
rect 22222 24392 22234 24395
rect 22646 24392 22652 24404
rect 22222 24364 22652 24392
rect 22222 24361 22234 24364
rect 22176 24355 22234 24361
rect 22646 24352 22652 24364
rect 22704 24352 22710 24404
rect 11330 24284 11336 24336
rect 11388 24324 11394 24336
rect 11425 24327 11483 24333
rect 11425 24324 11437 24327
rect 11388 24296 11437 24324
rect 11388 24284 11394 24296
rect 11425 24293 11437 24296
rect 11471 24293 11483 24327
rect 11425 24287 11483 24293
rect 23382 24284 23388 24336
rect 23440 24324 23446 24336
rect 25133 24327 25191 24333
rect 25133 24324 25145 24327
rect 23440 24296 25145 24324
rect 23440 24284 23446 24296
rect 25133 24293 25145 24296
rect 25179 24293 25191 24327
rect 25133 24287 25191 24293
rect 9548 24228 10456 24256
rect 9548 24216 9554 24228
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11977 24259 12035 24265
rect 11977 24256 11989 24259
rect 11112 24228 11989 24256
rect 11112 24216 11118 24228
rect 11977 24225 11989 24228
rect 12023 24256 12035 24259
rect 12342 24256 12348 24268
rect 12023 24228 12348 24256
rect 12023 24225 12035 24228
rect 11977 24219 12035 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 18966 24256 18972 24268
rect 18831 24228 18972 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 19426 24216 19432 24268
rect 19484 24216 19490 24268
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 22186 24256 22192 24268
rect 21959 24228 22192 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 22186 24216 22192 24228
rect 22244 24216 22250 24268
rect 22278 24216 22284 24268
rect 22336 24256 22342 24268
rect 22646 24256 22652 24268
rect 22336 24228 22652 24256
rect 22336 24216 22342 24228
rect 22646 24216 22652 24228
rect 22704 24216 22710 24268
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 7892 24160 9137 24188
rect 7892 24148 7898 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 17678 24148 17684 24200
rect 17736 24148 17742 24200
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 24857 24191 24915 24197
rect 24857 24157 24869 24191
rect 24903 24188 24915 24191
rect 25317 24191 25375 24197
rect 25317 24188 25329 24191
rect 24903 24160 25329 24188
rect 24903 24157 24915 24160
rect 24857 24151 24915 24157
rect 25317 24157 25329 24160
rect 25363 24188 25375 24191
rect 25406 24188 25412 24200
rect 25363 24160 25412 24188
rect 25363 24157 25375 24160
rect 25317 24151 25375 24157
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 9858 24120 9864 24132
rect 9600 24092 9864 24120
rect 9600 24064 9628 24092
rect 9858 24080 9864 24092
rect 9916 24080 9922 24132
rect 11330 24120 11336 24132
rect 10796 24092 11336 24120
rect 9582 24012 9588 24064
rect 9640 24052 9646 24064
rect 10796 24052 10824 24092
rect 11330 24080 11336 24092
rect 11388 24080 11394 24132
rect 11974 24080 11980 24132
rect 12032 24120 12038 24132
rect 12253 24123 12311 24129
rect 12253 24120 12265 24123
rect 12032 24092 12265 24120
rect 12032 24080 12038 24092
rect 12253 24089 12265 24092
rect 12299 24089 12311 24123
rect 13538 24120 13544 24132
rect 13478 24092 13544 24120
rect 12253 24083 12311 24089
rect 13538 24080 13544 24092
rect 13596 24120 13602 24132
rect 15933 24123 15991 24129
rect 13596 24092 14136 24120
rect 13596 24080 13602 24092
rect 14108 24064 14136 24092
rect 15933 24089 15945 24123
rect 15979 24120 15991 24123
rect 18874 24120 18880 24132
rect 15979 24092 18880 24120
rect 15979 24089 15991 24092
rect 15933 24083 15991 24089
rect 18874 24080 18880 24092
rect 18932 24080 18938 24132
rect 19702 24080 19708 24132
rect 19760 24080 19766 24132
rect 21082 24120 21088 24132
rect 20930 24092 21088 24120
rect 21082 24080 21088 24092
rect 21140 24120 21146 24132
rect 21140 24092 21588 24120
rect 21140 24080 21146 24092
rect 9640 24024 10824 24052
rect 10873 24055 10931 24061
rect 9640 24012 9646 24024
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11054 24052 11060 24064
rect 10919 24024 11060 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 13725 24055 13783 24061
rect 13725 24021 13737 24055
rect 13771 24052 13783 24055
rect 13906 24052 13912 24064
rect 13771 24024 13912 24052
rect 13771 24021 13783 24024
rect 13725 24015 13783 24021
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 14090 24012 14096 24064
rect 14148 24012 14154 24064
rect 18141 24055 18199 24061
rect 18141 24021 18153 24055
rect 18187 24052 18199 24055
rect 18506 24052 18512 24064
rect 18187 24024 18512 24052
rect 18187 24021 18199 24024
rect 18141 24015 18199 24021
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 20530 24052 20536 24064
rect 18647 24024 20536 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 20530 24012 20536 24024
rect 20588 24012 20594 24064
rect 21560 24061 21588 24092
rect 22296 24092 22678 24120
rect 22296 24064 22324 24092
rect 21545 24055 21603 24061
rect 21545 24021 21557 24055
rect 21591 24052 21603 24055
rect 22278 24052 22284 24064
rect 21591 24024 22284 24052
rect 21591 24021 21603 24024
rect 21545 24015 21603 24021
rect 22278 24012 22284 24024
rect 22336 24012 22342 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23624 24024 23673 24052
rect 23624 24012 23630 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 9769 23851 9827 23857
rect 9769 23848 9781 23851
rect 9732 23820 9781 23848
rect 9732 23808 9738 23820
rect 9769 23817 9781 23820
rect 9815 23817 9827 23851
rect 9769 23811 9827 23817
rect 9582 23780 9588 23792
rect 9522 23752 9588 23780
rect 9582 23740 9588 23752
rect 9640 23740 9646 23792
rect 7834 23672 7840 23724
rect 7892 23712 7898 23724
rect 8021 23715 8079 23721
rect 8021 23712 8033 23715
rect 7892 23684 8033 23712
rect 7892 23672 7898 23684
rect 8021 23681 8033 23684
rect 8067 23681 8079 23715
rect 9784 23712 9812 23811
rect 10410 23808 10416 23860
rect 10468 23808 10474 23860
rect 10781 23851 10839 23857
rect 10781 23817 10793 23851
rect 10827 23848 10839 23851
rect 13814 23848 13820 23860
rect 10827 23820 13820 23848
rect 10827 23817 10839 23820
rect 10781 23811 10839 23817
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23817 14519 23851
rect 14461 23811 14519 23817
rect 11146 23740 11152 23792
rect 11204 23780 11210 23792
rect 11609 23783 11667 23789
rect 11609 23780 11621 23783
rect 11204 23752 11621 23780
rect 11204 23740 11210 23752
rect 11609 23749 11621 23752
rect 11655 23780 11667 23783
rect 11790 23780 11796 23792
rect 11655 23752 11796 23780
rect 11655 23749 11667 23752
rect 11609 23743 11667 23749
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 13633 23783 13691 23789
rect 13633 23749 13645 23783
rect 13679 23780 13691 23783
rect 14274 23780 14280 23792
rect 13679 23752 14280 23780
rect 13679 23749 13691 23752
rect 13633 23743 13691 23749
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 14476 23780 14504 23811
rect 14918 23808 14924 23860
rect 14976 23808 14982 23860
rect 16574 23808 16580 23860
rect 16632 23848 16638 23860
rect 17310 23848 17316 23860
rect 16632 23820 17316 23848
rect 16632 23808 16638 23820
rect 17310 23808 17316 23820
rect 17368 23848 17374 23860
rect 18693 23851 18751 23857
rect 18693 23848 18705 23851
rect 17368 23820 18705 23848
rect 17368 23808 17374 23820
rect 18693 23817 18705 23820
rect 18739 23817 18751 23851
rect 18693 23811 18751 23817
rect 18708 23780 18736 23811
rect 18874 23808 18880 23860
rect 18932 23808 18938 23860
rect 19794 23848 19800 23860
rect 19352 23820 19800 23848
rect 19242 23780 19248 23792
rect 14476 23752 18276 23780
rect 18708 23752 19248 23780
rect 10686 23712 10692 23724
rect 9784 23684 10692 23712
rect 8021 23675 8079 23681
rect 10686 23672 10692 23684
rect 10744 23712 10750 23724
rect 10744 23684 11008 23712
rect 10744 23672 10750 23684
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23644 8355 23647
rect 8343 23616 9996 23644
rect 8343 23613 8355 23616
rect 8297 23607 8355 23613
rect 9968 23576 9996 23616
rect 10042 23604 10048 23656
rect 10100 23644 10106 23656
rect 10980 23653 11008 23684
rect 13722 23672 13728 23724
rect 13780 23672 13786 23724
rect 14182 23672 14188 23724
rect 14240 23712 14246 23724
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 14240 23684 14841 23712
rect 14240 23672 14246 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 14918 23672 14924 23724
rect 14976 23712 14982 23724
rect 16666 23712 16672 23724
rect 14976 23684 16672 23712
rect 14976 23672 14982 23684
rect 16666 23672 16672 23684
rect 16724 23712 16730 23724
rect 18248 23721 18276 23752
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 17221 23715 17279 23721
rect 17221 23712 17233 23715
rect 16724 23684 17233 23712
rect 16724 23672 16730 23684
rect 17221 23681 17233 23684
rect 17267 23712 17279 23715
rect 18233 23715 18291 23721
rect 17267 23684 17540 23712
rect 17267 23681 17279 23684
rect 17221 23675 17279 23681
rect 10873 23647 10931 23653
rect 10873 23644 10885 23647
rect 10100 23616 10885 23644
rect 10100 23604 10106 23616
rect 10873 23613 10885 23616
rect 10919 23613 10931 23647
rect 10873 23607 10931 23613
rect 10965 23647 11023 23653
rect 10965 23613 10977 23647
rect 11011 23613 11023 23647
rect 10965 23607 11023 23613
rect 13817 23647 13875 23653
rect 13817 23613 13829 23647
rect 13863 23613 13875 23647
rect 13817 23607 13875 23613
rect 11146 23576 11152 23588
rect 9968 23548 11152 23576
rect 11146 23536 11152 23548
rect 11204 23536 11210 23588
rect 12894 23536 12900 23588
rect 12952 23576 12958 23588
rect 13832 23576 13860 23607
rect 13906 23604 13912 23656
rect 13964 23644 13970 23656
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 13964 23616 15025 23644
rect 13964 23604 13970 23616
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 15654 23604 15660 23656
rect 15712 23604 15718 23656
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23613 17463 23647
rect 17512 23644 17540 23684
rect 18233 23681 18245 23715
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 18601 23715 18659 23721
rect 18601 23681 18613 23715
rect 18647 23712 18659 23715
rect 19352 23712 19380 23820
rect 19794 23808 19800 23820
rect 19852 23808 19858 23860
rect 20901 23851 20959 23857
rect 20901 23817 20913 23851
rect 20947 23848 20959 23851
rect 21910 23848 21916 23860
rect 20947 23820 21916 23848
rect 20947 23817 20959 23820
rect 20901 23811 20959 23817
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23848 22247 23851
rect 23842 23848 23848 23860
rect 22235 23820 23848 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24949 23851 25007 23857
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 25038 23848 25044 23860
rect 24995 23820 25044 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 25038 23808 25044 23820
rect 25096 23808 25102 23860
rect 25314 23808 25320 23860
rect 25372 23848 25378 23860
rect 25409 23851 25467 23857
rect 25409 23848 25421 23851
rect 25372 23820 25421 23848
rect 25372 23808 25378 23820
rect 25409 23817 25421 23820
rect 25455 23817 25467 23851
rect 25409 23811 25467 23817
rect 19702 23740 19708 23792
rect 19760 23780 19766 23792
rect 22738 23780 22744 23792
rect 19760 23752 20116 23780
rect 19760 23740 19766 23752
rect 18647 23684 19380 23712
rect 18647 23681 18659 23684
rect 18601 23675 18659 23681
rect 18616 23644 18644 23675
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 19978 23716 19984 23724
rect 19904 23712 19984 23716
rect 19720 23688 19984 23712
rect 19720 23684 19932 23688
rect 19720 23656 19748 23684
rect 19978 23672 19984 23688
rect 20036 23672 20042 23724
rect 17512 23616 18644 23644
rect 17405 23607 17463 23613
rect 12952 23548 13860 23576
rect 12952 23536 12958 23548
rect 15470 23536 15476 23588
rect 15528 23576 15534 23588
rect 17420 23576 17448 23607
rect 19702 23604 19708 23656
rect 19760 23604 19766 23656
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23644 19947 23647
rect 20088 23644 20116 23752
rect 20548 23752 22744 23780
rect 20548 23644 20576 23752
rect 22738 23740 22744 23752
rect 22796 23780 22802 23792
rect 23198 23780 23204 23792
rect 22796 23752 23204 23780
rect 22796 23740 22802 23752
rect 23198 23740 23204 23752
rect 23256 23740 23262 23792
rect 23934 23740 23940 23792
rect 23992 23740 23998 23792
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 22186 23672 22192 23724
rect 22244 23712 22250 23724
rect 22373 23715 22431 23721
rect 22244 23684 22324 23712
rect 22244 23672 22250 23684
rect 19935 23616 20576 23644
rect 19935 23613 19947 23616
rect 19889 23607 19947 23613
rect 20990 23604 20996 23656
rect 21048 23604 21054 23656
rect 22296 23644 22324 23684
rect 22373 23681 22385 23715
rect 22419 23712 22431 23715
rect 22646 23712 22652 23724
rect 22419 23684 22652 23712
rect 22419 23681 22431 23684
rect 22373 23675 22431 23681
rect 22646 23672 22652 23684
rect 22704 23672 22710 23724
rect 22830 23644 22836 23656
rect 22296 23616 22836 23644
rect 22830 23604 22836 23616
rect 22888 23644 22894 23656
rect 23201 23647 23259 23653
rect 23201 23644 23213 23647
rect 22888 23616 23213 23644
rect 22888 23604 22894 23616
rect 23201 23613 23213 23616
rect 23247 23613 23259 23647
rect 23201 23607 23259 23613
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 23566 23644 23572 23656
rect 23523 23616 23572 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 23566 23604 23572 23616
rect 23624 23604 23630 23656
rect 15528 23548 17448 23576
rect 18049 23579 18107 23585
rect 15528 23536 15534 23548
rect 18049 23545 18061 23579
rect 18095 23576 18107 23579
rect 21174 23576 21180 23588
rect 18095 23548 21180 23576
rect 18095 23545 18107 23548
rect 18049 23539 18107 23545
rect 21174 23536 21180 23548
rect 21232 23536 21238 23588
rect 9582 23468 9588 23520
rect 9640 23508 9646 23520
rect 10045 23511 10103 23517
rect 10045 23508 10057 23511
rect 9640 23480 10057 23508
rect 9640 23468 9646 23480
rect 10045 23477 10057 23480
rect 10091 23508 10103 23511
rect 10134 23508 10140 23520
rect 10091 23480 10140 23508
rect 10091 23477 10103 23480
rect 10045 23471 10103 23477
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 12802 23468 12808 23520
rect 12860 23508 12866 23520
rect 13265 23511 13323 23517
rect 13265 23508 13277 23511
rect 12860 23480 13277 23508
rect 12860 23468 12866 23480
rect 13265 23477 13277 23480
rect 13311 23477 13323 23511
rect 13265 23471 13323 23477
rect 16853 23511 16911 23517
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 17310 23508 17316 23520
rect 16899 23480 17316 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 19245 23511 19303 23517
rect 19245 23477 19257 23511
rect 19291 23508 19303 23511
rect 19886 23508 19892 23520
rect 19291 23480 19892 23508
rect 19291 23477 19303 23480
rect 19245 23471 19303 23477
rect 19886 23468 19892 23480
rect 19944 23468 19950 23520
rect 20254 23468 20260 23520
rect 20312 23508 20318 23520
rect 20441 23511 20499 23517
rect 20441 23508 20453 23511
rect 20312 23480 20453 23508
rect 20312 23468 20318 23480
rect 20441 23477 20453 23480
rect 20487 23477 20499 23511
rect 20441 23471 20499 23477
rect 21913 23511 21971 23517
rect 21913 23477 21925 23511
rect 21959 23508 21971 23511
rect 22278 23508 22284 23520
rect 21959 23480 22284 23508
rect 21959 23477 21971 23480
rect 21913 23471 21971 23477
rect 22278 23468 22284 23480
rect 22336 23508 22342 23520
rect 22833 23511 22891 23517
rect 22833 23508 22845 23511
rect 22336 23480 22845 23508
rect 22336 23468 22342 23480
rect 22833 23477 22845 23480
rect 22879 23508 22891 23511
rect 23934 23508 23940 23520
rect 22879 23480 23940 23508
rect 22879 23477 22891 23480
rect 22833 23471 22891 23477
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 25314 23468 25320 23520
rect 25372 23508 25378 23520
rect 25958 23508 25964 23520
rect 25372 23480 25964 23508
rect 25372 23468 25378 23480
rect 25958 23468 25964 23480
rect 26016 23468 26022 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 10594 23264 10600 23316
rect 10652 23304 10658 23316
rect 10781 23307 10839 23313
rect 10781 23304 10793 23307
rect 10652 23276 10793 23304
rect 10652 23264 10658 23276
rect 10781 23273 10793 23276
rect 10827 23273 10839 23307
rect 10781 23267 10839 23273
rect 15841 23307 15899 23313
rect 15841 23273 15853 23307
rect 15887 23304 15899 23307
rect 17218 23304 17224 23316
rect 15887 23276 17224 23304
rect 15887 23273 15899 23276
rect 15841 23267 15899 23273
rect 9582 23196 9588 23248
rect 9640 23236 9646 23248
rect 9640 23208 12434 23236
rect 9640 23196 9646 23208
rect 6178 23128 6184 23180
rect 6236 23168 6242 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 6236 23140 9689 23168
rect 6236 23128 6242 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 9309 23103 9367 23109
rect 9309 23069 9321 23103
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 9324 22964 9352 23063
rect 9692 23032 9720 23131
rect 11698 23128 11704 23180
rect 11756 23128 11762 23180
rect 11790 23128 11796 23180
rect 11848 23128 11854 23180
rect 12406 23168 12434 23208
rect 12526 23196 12532 23248
rect 12584 23236 12590 23248
rect 14737 23239 14795 23245
rect 14737 23236 14749 23239
rect 12584 23208 14749 23236
rect 12584 23196 12590 23208
rect 14737 23205 14749 23208
rect 14783 23205 14795 23239
rect 14737 23199 14795 23205
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 12406 23140 13553 23168
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 13541 23131 13599 23137
rect 14384 23140 15301 23168
rect 14384 23112 14412 23140
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 11609 23103 11667 23109
rect 11609 23069 11621 23103
rect 11655 23100 11667 23103
rect 14274 23100 14280 23112
rect 11655 23072 14280 23100
rect 11655 23069 11667 23072
rect 11609 23063 11667 23069
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 14366 23060 14372 23112
rect 14424 23060 14430 23112
rect 15105 23103 15163 23109
rect 15105 23069 15117 23103
rect 15151 23100 15163 23103
rect 15654 23100 15660 23112
rect 15151 23072 15660 23100
rect 15151 23069 15163 23072
rect 15105 23063 15163 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 13262 23032 13268 23044
rect 9692 23004 13268 23032
rect 13262 22992 13268 23004
rect 13320 22992 13326 23044
rect 13357 23035 13415 23041
rect 13357 23001 13369 23035
rect 13403 23032 13415 23035
rect 14918 23032 14924 23044
rect 13403 23004 14924 23032
rect 13403 23001 13415 23004
rect 13357 22995 13415 23001
rect 14918 22992 14924 23004
rect 14976 22992 14982 23044
rect 15197 23035 15255 23041
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 15856 23032 15884 23267
rect 17218 23264 17224 23276
rect 17276 23304 17282 23316
rect 25774 23304 25780 23316
rect 17276 23276 25780 23304
rect 17276 23264 17282 23276
rect 25774 23264 25780 23276
rect 25832 23264 25838 23316
rect 17865 23239 17923 23245
rect 17865 23205 17877 23239
rect 17911 23236 17923 23239
rect 18322 23236 18328 23248
rect 17911 23208 18328 23236
rect 17911 23205 17923 23208
rect 17865 23199 17923 23205
rect 18322 23196 18328 23208
rect 18380 23196 18386 23248
rect 18414 23196 18420 23248
rect 18472 23236 18478 23248
rect 19521 23239 19579 23245
rect 19521 23236 19533 23239
rect 18472 23208 19533 23236
rect 18472 23196 18478 23208
rect 19521 23205 19533 23208
rect 19567 23205 19579 23239
rect 19521 23199 19579 23205
rect 18509 23171 18567 23177
rect 18509 23137 18521 23171
rect 18555 23168 18567 23171
rect 18690 23168 18696 23180
rect 18555 23140 18696 23168
rect 18555 23137 18567 23140
rect 18509 23131 18567 23137
rect 18690 23128 18696 23140
rect 18748 23128 18754 23180
rect 18969 23171 19027 23177
rect 18969 23137 18981 23171
rect 19015 23168 19027 23171
rect 19702 23168 19708 23180
rect 19015 23140 19708 23168
rect 19015 23137 19027 23140
rect 18969 23131 19027 23137
rect 19702 23128 19708 23140
rect 19760 23128 19766 23180
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23168 20223 23171
rect 20438 23168 20444 23180
rect 20211 23140 20444 23168
rect 20211 23137 20223 23140
rect 20165 23131 20223 23137
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23168 20775 23171
rect 20806 23168 20812 23180
rect 20763 23140 20812 23168
rect 20763 23137 20775 23140
rect 20717 23131 20775 23137
rect 20806 23128 20812 23140
rect 20864 23128 20870 23180
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25406 23168 25412 23180
rect 25271 23140 25412 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25406 23128 25412 23140
rect 25464 23128 25470 23180
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 18782 23100 18788 23112
rect 18288 23072 18788 23100
rect 18288 23060 18294 23072
rect 18782 23060 18788 23072
rect 18840 23060 18846 23112
rect 19886 23060 19892 23112
rect 19944 23060 19950 23112
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23100 20039 23103
rect 21634 23100 21640 23112
rect 20027 23072 21640 23100
rect 20027 23069 20039 23072
rect 19981 23063 20039 23069
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 15243 23004 15884 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 16850 22992 16856 23044
rect 16908 23032 16914 23044
rect 21836 23032 21864 23063
rect 22830 23060 22836 23112
rect 22888 23060 22894 23112
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23100 25099 23103
rect 25682 23100 25688 23112
rect 25087 23072 25688 23100
rect 25087 23069 25099 23072
rect 25041 23063 25099 23069
rect 25682 23060 25688 23072
rect 25740 23060 25746 23112
rect 16908 23004 21864 23032
rect 23845 23035 23903 23041
rect 16908 22992 16914 23004
rect 23845 23001 23857 23035
rect 23891 23032 23903 23035
rect 24854 23032 24860 23044
rect 23891 23004 24860 23032
rect 23891 23001 23903 23004
rect 23845 22995 23903 23001
rect 24854 22992 24860 23004
rect 24912 22992 24918 23044
rect 24949 23035 25007 23041
rect 24949 23001 24961 23035
rect 24995 23032 25007 23035
rect 25314 23032 25320 23044
rect 24995 23004 25320 23032
rect 24995 23001 25007 23004
rect 24949 22995 25007 23001
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 10594 22964 10600 22976
rect 9324 22936 10600 22964
rect 10594 22924 10600 22936
rect 10652 22924 10658 22976
rect 10870 22924 10876 22976
rect 10928 22964 10934 22976
rect 11241 22967 11299 22973
rect 11241 22964 11253 22967
rect 10928 22936 11253 22964
rect 10928 22924 10934 22936
rect 11241 22933 11253 22936
rect 11287 22933 11299 22967
rect 11241 22927 11299 22933
rect 12066 22924 12072 22976
rect 12124 22964 12130 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12124 22936 13001 22964
rect 12124 22924 12130 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 13449 22967 13507 22973
rect 13449 22933 13461 22967
rect 13495 22964 13507 22967
rect 14185 22967 14243 22973
rect 14185 22964 14197 22967
rect 13495 22936 14197 22964
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 14185 22933 14197 22936
rect 14231 22964 14243 22967
rect 16574 22964 16580 22976
rect 14231 22936 16580 22964
rect 14231 22933 14243 22936
rect 14185 22927 14243 22933
rect 16574 22924 16580 22936
rect 16632 22924 16638 22976
rect 18325 22967 18383 22973
rect 18325 22933 18337 22967
rect 18371 22964 18383 22967
rect 19058 22964 19064 22976
rect 18371 22936 19064 22964
rect 18371 22933 18383 22936
rect 18325 22927 18383 22933
rect 19058 22924 19064 22936
rect 19116 22924 19122 22976
rect 21637 22967 21695 22973
rect 21637 22933 21649 22967
rect 21683 22964 21695 22967
rect 22094 22964 22100 22976
rect 21683 22936 22100 22964
rect 21683 22933 21695 22936
rect 21637 22927 21695 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 23532 22936 24593 22964
rect 23532 22924 23538 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 10134 22720 10140 22772
rect 10192 22720 10198 22772
rect 11330 22720 11336 22772
rect 11388 22760 11394 22772
rect 14366 22760 14372 22772
rect 11388 22732 14372 22760
rect 11388 22720 11394 22732
rect 14366 22720 14372 22732
rect 14424 22720 14430 22772
rect 14461 22763 14519 22769
rect 14461 22729 14473 22763
rect 14507 22760 14519 22763
rect 14918 22760 14924 22772
rect 14507 22732 14924 22760
rect 14507 22729 14519 22732
rect 14461 22723 14519 22729
rect 14918 22720 14924 22732
rect 14976 22720 14982 22772
rect 16850 22720 16856 22772
rect 16908 22720 16914 22772
rect 18782 22720 18788 22772
rect 18840 22720 18846 22772
rect 18877 22763 18935 22769
rect 18877 22729 18889 22763
rect 18923 22760 18935 22763
rect 19058 22760 19064 22772
rect 18923 22732 19064 22760
rect 18923 22729 18935 22732
rect 18877 22723 18935 22729
rect 19058 22720 19064 22732
rect 19116 22720 19122 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19668 22732 19717 22760
rect 19668 22720 19674 22732
rect 19705 22729 19717 22732
rect 19751 22729 19763 22763
rect 19705 22723 19763 22729
rect 21177 22763 21235 22769
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 23382 22760 23388 22772
rect 21223 22732 23388 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7892 22596 8125 22624
rect 7892 22584 7898 22596
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 9490 22584 9496 22636
rect 9548 22624 9554 22636
rect 10152 22624 10180 22720
rect 14090 22692 14096 22704
rect 13846 22664 14096 22692
rect 14090 22652 14096 22664
rect 14148 22692 14154 22704
rect 14642 22692 14648 22704
rect 14148 22664 14648 22692
rect 14148 22652 14154 22664
rect 14642 22652 14648 22664
rect 14700 22652 14706 22704
rect 19076 22692 19104 22720
rect 21450 22692 21456 22704
rect 19076 22664 21456 22692
rect 21450 22652 21456 22664
rect 21508 22652 21514 22704
rect 25130 22652 25136 22704
rect 25188 22652 25194 22704
rect 9548 22596 10180 22624
rect 9548 22584 9554 22596
rect 12342 22584 12348 22636
rect 12400 22584 12406 22636
rect 15286 22584 15292 22636
rect 15344 22624 15350 22636
rect 17037 22627 17095 22633
rect 17037 22624 17049 22627
rect 15344 22596 17049 22624
rect 15344 22584 15350 22596
rect 17037 22593 17049 22596
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 19058 22584 19064 22636
rect 19116 22624 19122 22636
rect 19702 22624 19708 22636
rect 19116 22596 19708 22624
rect 19116 22584 19122 22596
rect 19702 22584 19708 22596
rect 19760 22584 19766 22636
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 19904 22596 21097 22624
rect 8389 22559 8447 22565
rect 8389 22525 8401 22559
rect 8435 22556 8447 22559
rect 11238 22556 11244 22568
rect 8435 22528 11244 22556
rect 8435 22525 8447 22528
rect 8389 22519 8447 22525
rect 11238 22516 11244 22528
rect 11296 22516 11302 22568
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 13354 22556 13360 22568
rect 12667 22528 13360 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 18782 22516 18788 22568
rect 18840 22556 18846 22568
rect 18966 22556 18972 22568
rect 18840 22528 18972 22556
rect 18840 22516 18846 22528
rect 18966 22516 18972 22528
rect 19024 22516 19030 22568
rect 11790 22488 11796 22500
rect 9876 22460 11796 22488
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 9876 22429 9904 22460
rect 11790 22448 11796 22460
rect 11848 22448 11854 22500
rect 19904 22488 19932 22596
rect 21085 22593 21097 22596
rect 21131 22624 21143 22627
rect 21542 22624 21548 22636
rect 21131 22596 21548 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 23842 22584 23848 22636
rect 23900 22624 23906 22636
rect 23937 22627 23995 22633
rect 23937 22624 23949 22627
rect 23900 22596 23949 22624
rect 23900 22584 23906 22596
rect 23937 22593 23949 22596
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 19978 22516 19984 22568
rect 20036 22556 20042 22568
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 20036 22528 21281 22556
rect 20036 22516 20042 22528
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 23290 22516 23296 22568
rect 23348 22516 23354 22568
rect 20349 22491 20407 22497
rect 20349 22488 20361 22491
rect 14016 22460 20361 22488
rect 9861 22423 9919 22429
rect 9861 22420 9873 22423
rect 6972 22392 9873 22420
rect 6972 22380 6978 22392
rect 9861 22389 9873 22392
rect 9907 22389 9919 22423
rect 9861 22383 9919 22389
rect 13262 22380 13268 22432
rect 13320 22420 13326 22432
rect 14016 22420 14044 22460
rect 20349 22457 20361 22460
rect 20395 22457 20407 22491
rect 20349 22451 20407 22457
rect 13320 22392 14044 22420
rect 13320 22380 13326 22392
rect 14090 22380 14096 22432
rect 14148 22380 14154 22432
rect 14642 22380 14648 22432
rect 14700 22380 14706 22432
rect 16114 22380 16120 22432
rect 16172 22420 16178 22432
rect 17034 22420 17040 22432
rect 16172 22392 17040 22420
rect 16172 22380 16178 22392
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 11054 22176 11060 22228
rect 11112 22216 11118 22228
rect 11112 22188 12388 22216
rect 11112 22176 11118 22188
rect 11514 22148 11520 22160
rect 11348 22120 11520 22148
rect 8662 22040 8668 22092
rect 8720 22080 8726 22092
rect 11348 22089 11376 22120
rect 11514 22108 11520 22120
rect 11572 22108 11578 22160
rect 9677 22083 9735 22089
rect 9677 22080 9689 22083
rect 8720 22052 9689 22080
rect 8720 22040 8726 22052
rect 9677 22049 9689 22052
rect 9723 22049 9735 22083
rect 9677 22043 9735 22049
rect 11333 22083 11391 22089
rect 11333 22049 11345 22083
rect 11379 22080 11391 22083
rect 11379 22052 11413 22080
rect 11992 22052 12296 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 10410 21972 10416 22024
rect 10468 22012 10474 22024
rect 11149 22015 11207 22021
rect 11149 22012 11161 22015
rect 10468 21984 11161 22012
rect 10468 21972 10474 21984
rect 11149 21981 11161 21984
rect 11195 21981 11207 22015
rect 11149 21975 11207 21981
rect 9585 21947 9643 21953
rect 9585 21913 9597 21947
rect 9631 21944 9643 21947
rect 11790 21944 11796 21956
rect 9631 21916 11796 21944
rect 9631 21913 9643 21916
rect 9585 21907 9643 21913
rect 11790 21904 11796 21916
rect 11848 21904 11854 21956
rect 9125 21879 9183 21885
rect 9125 21845 9137 21879
rect 9171 21876 9183 21879
rect 9214 21876 9220 21888
rect 9171 21848 9220 21876
rect 9171 21845 9183 21848
rect 9125 21839 9183 21845
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 9493 21879 9551 21885
rect 9493 21845 9505 21879
rect 9539 21876 9551 21879
rect 10134 21876 10140 21888
rect 9539 21848 10140 21876
rect 9539 21845 9551 21848
rect 9493 21839 9551 21845
rect 10134 21836 10140 21848
rect 10192 21836 10198 21888
rect 10410 21836 10416 21888
rect 10468 21836 10474 21888
rect 10689 21879 10747 21885
rect 10689 21845 10701 21879
rect 10735 21876 10747 21879
rect 10778 21876 10784 21888
rect 10735 21848 10784 21876
rect 10735 21845 10747 21848
rect 10689 21839 10747 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 11054 21836 11060 21888
rect 11112 21836 11118 21888
rect 11992 21885 12020 22052
rect 12268 21944 12296 22052
rect 12360 22012 12388 22188
rect 16206 22176 16212 22228
rect 16264 22216 16270 22228
rect 21808 22219 21866 22225
rect 16264 22188 17448 22216
rect 16264 22176 16270 22188
rect 12802 22148 12808 22160
rect 12452 22120 12808 22148
rect 12452 22089 12480 22120
rect 12802 22108 12808 22120
rect 12860 22108 12866 22160
rect 15562 22148 15568 22160
rect 15304 22120 15568 22148
rect 15304 22089 15332 22120
rect 15562 22108 15568 22120
rect 15620 22108 15626 22160
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 12529 22083 12587 22089
rect 12529 22049 12541 22083
rect 12575 22049 12587 22083
rect 12529 22043 12587 22049
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 15381 22083 15439 22089
rect 15381 22049 15393 22083
rect 15427 22049 15439 22083
rect 15381 22043 15439 22049
rect 16117 22083 16175 22089
rect 16117 22049 16129 22083
rect 16163 22080 16175 22083
rect 16758 22080 16764 22092
rect 16163 22052 16764 22080
rect 16163 22049 16175 22052
rect 16117 22043 16175 22049
rect 12544 22012 12572 22043
rect 12360 21984 12572 22012
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 15396 22012 15424 22043
rect 16758 22040 16764 22052
rect 16816 22040 16822 22092
rect 17420 22080 17448 22188
rect 21808 22185 21820 22219
rect 21854 22216 21866 22219
rect 23106 22216 23112 22228
rect 21854 22188 23112 22216
rect 21854 22185 21866 22188
rect 21808 22179 21866 22185
rect 23106 22176 23112 22188
rect 23164 22176 23170 22228
rect 23293 22219 23351 22225
rect 23293 22185 23305 22219
rect 23339 22216 23351 22219
rect 23382 22216 23388 22228
rect 23339 22188 23388 22216
rect 23339 22185 23351 22188
rect 23293 22179 23351 22185
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 25222 22216 25228 22228
rect 25148 22188 25228 22216
rect 20530 22148 20536 22160
rect 20364 22120 20536 22148
rect 18598 22080 18604 22092
rect 17420 22052 18604 22080
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 20364 22089 20392 22120
rect 20530 22108 20536 22120
rect 20588 22108 20594 22160
rect 25148 22094 25176 22188
rect 25222 22176 25228 22188
rect 25280 22176 25286 22228
rect 20349 22083 20407 22089
rect 20349 22049 20361 22083
rect 20395 22049 20407 22083
rect 20349 22043 20407 22049
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22080 21603 22083
rect 22186 22080 22192 22092
rect 21591 22052 22192 22080
rect 21591 22049 21603 22052
rect 21545 22043 21603 22049
rect 22186 22040 22192 22052
rect 22244 22080 22250 22092
rect 23014 22080 23020 22092
rect 22244 22052 23020 22080
rect 22244 22040 22250 22052
rect 23014 22040 23020 22052
rect 23072 22040 23078 22092
rect 24854 22040 24860 22092
rect 24912 22080 24918 22092
rect 25148 22089 25268 22094
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 24912 22052 25053 22080
rect 24912 22040 24918 22052
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25148 22083 25283 22089
rect 25148 22066 25237 22083
rect 25041 22043 25099 22049
rect 25225 22049 25237 22066
rect 25271 22049 25283 22083
rect 25225 22043 25283 22049
rect 14148 21984 15424 22012
rect 14148 21972 14154 21984
rect 17494 21972 17500 22024
rect 17552 22012 17558 22024
rect 18141 22015 18199 22021
rect 18141 22012 18153 22015
rect 17552 21984 18153 22012
rect 17552 21972 17558 21984
rect 18141 21981 18153 21984
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23845 22015 23903 22021
rect 23845 22012 23857 22015
rect 23256 21984 23857 22012
rect 23256 21972 23262 21984
rect 23845 21981 23857 21984
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 15286 21944 15292 21956
rect 12268 21916 15292 21944
rect 15286 21904 15292 21916
rect 15344 21904 15350 21956
rect 16393 21947 16451 21953
rect 16393 21944 16405 21947
rect 16224 21916 16405 21944
rect 16224 21888 16252 21916
rect 16393 21913 16405 21916
rect 16439 21913 16451 21947
rect 21358 21944 21364 21956
rect 16393 21907 16451 21913
rect 19720 21916 21364 21944
rect 11977 21879 12035 21885
rect 11977 21845 11989 21879
rect 12023 21845 12035 21879
rect 11977 21839 12035 21845
rect 12342 21836 12348 21888
rect 12400 21836 12406 21888
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 16206 21836 16212 21888
rect 16264 21836 16270 21888
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 19720 21885 19748 21916
rect 21358 21904 21364 21916
rect 21416 21904 21422 21956
rect 22278 21904 22284 21956
rect 22336 21904 22342 21956
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 23216 21916 24961 21944
rect 17865 21879 17923 21885
rect 17865 21876 17877 21879
rect 17184 21848 17877 21876
rect 17184 21836 17190 21848
rect 17865 21845 17877 21848
rect 17911 21845 17923 21879
rect 17865 21839 17923 21845
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21845 19763 21879
rect 19705 21839 19763 21845
rect 20070 21836 20076 21888
rect 20128 21836 20134 21888
rect 20162 21836 20168 21888
rect 20220 21836 20226 21888
rect 20901 21879 20959 21885
rect 20901 21845 20913 21879
rect 20947 21876 20959 21879
rect 23216 21876 23244 21916
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 20947 21848 23244 21876
rect 20947 21845 20959 21848
rect 20901 21839 20959 21845
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23348 21848 24593 21876
rect 23348 21836 23354 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10284 21644 10425 21672
rect 10284 21632 10290 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 10413 21635 10471 21641
rect 10781 21675 10839 21681
rect 10781 21641 10793 21675
rect 10827 21672 10839 21675
rect 10962 21672 10968 21684
rect 10827 21644 10968 21672
rect 10827 21641 10839 21644
rect 10781 21635 10839 21641
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 11054 21632 11060 21684
rect 11112 21672 11118 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 11112 21644 11713 21672
rect 11112 21632 11118 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 11790 21632 11796 21684
rect 11848 21672 11854 21684
rect 12710 21672 12716 21684
rect 11848 21644 12716 21672
rect 11848 21632 11854 21644
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 15197 21675 15255 21681
rect 15197 21672 15209 21675
rect 14752 21644 15209 21672
rect 8570 21604 8576 21616
rect 8418 21576 8576 21604
rect 8570 21564 8576 21576
rect 8628 21604 8634 21616
rect 9490 21604 9496 21616
rect 8628 21576 9496 21604
rect 8628 21564 8634 21576
rect 9490 21564 9496 21576
rect 9548 21564 9554 21616
rect 10873 21607 10931 21613
rect 10873 21573 10885 21607
rect 10919 21604 10931 21607
rect 12158 21604 12164 21616
rect 10919 21576 12164 21604
rect 10919 21573 10931 21576
rect 10873 21567 10931 21573
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 14642 21604 14648 21616
rect 14582 21576 14648 21604
rect 14642 21564 14648 21576
rect 14700 21604 14706 21616
rect 14752 21604 14780 21644
rect 15197 21641 15209 21644
rect 15243 21672 15255 21675
rect 15654 21672 15660 21684
rect 15243 21644 15660 21672
rect 15243 21641 15255 21644
rect 15197 21635 15255 21641
rect 15654 21632 15660 21644
rect 15712 21632 15718 21684
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 19153 21675 19211 21681
rect 19153 21672 19165 21675
rect 19116 21644 19165 21672
rect 19116 21632 19122 21644
rect 19153 21641 19165 21644
rect 19199 21672 19211 21675
rect 19981 21675 20039 21681
rect 19981 21672 19993 21675
rect 19199 21644 19993 21672
rect 19199 21641 19211 21644
rect 19153 21635 19211 21641
rect 19981 21641 19993 21644
rect 20027 21641 20039 21675
rect 19981 21635 20039 21641
rect 20070 21632 20076 21684
rect 20128 21672 20134 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 20128 21644 21189 21672
rect 20128 21632 20134 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 22554 21672 22560 21684
rect 22511 21644 22560 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 23106 21672 23112 21684
rect 22796 21644 23112 21672
rect 22796 21632 22802 21644
rect 23106 21632 23112 21644
rect 23164 21672 23170 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 23164 21644 25053 21672
rect 23164 21632 23170 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 14700 21576 14780 21604
rect 14700 21564 14706 21576
rect 14826 21564 14832 21616
rect 14884 21604 14890 21616
rect 14884 21576 16574 21604
rect 14884 21564 14890 21576
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9950 21536 9956 21548
rect 9631 21508 9956 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10686 21496 10692 21548
rect 10744 21536 10750 21548
rect 10744 21508 11100 21536
rect 10744 21496 10750 21508
rect 6917 21471 6975 21477
rect 6917 21437 6929 21471
rect 6963 21468 6975 21471
rect 7193 21471 7251 21477
rect 6963 21440 7052 21468
rect 6963 21437 6975 21440
rect 6917 21431 6975 21437
rect 7024 21332 7052 21440
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 8386 21468 8392 21480
rect 7239 21440 8392 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 8386 21428 8392 21440
rect 8444 21428 8450 21480
rect 8846 21428 8852 21480
rect 8904 21468 8910 21480
rect 11072 21477 11100 21508
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 13081 21539 13139 21545
rect 13081 21536 13093 21539
rect 12492 21508 13093 21536
rect 12492 21496 12498 21508
rect 13081 21505 13093 21508
rect 13127 21505 13139 21539
rect 13081 21499 13139 21505
rect 15657 21539 15715 21545
rect 15657 21505 15669 21539
rect 15703 21536 15715 21539
rect 15746 21536 15752 21548
rect 15703 21508 15752 21536
rect 15703 21505 15715 21508
rect 15657 21499 15715 21505
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 16546 21536 16574 21576
rect 18782 21564 18788 21616
rect 18840 21604 18846 21616
rect 20162 21604 20168 21616
rect 18840 21576 20168 21604
rect 18840 21564 18846 21576
rect 20162 21564 20168 21576
rect 20220 21604 20226 21616
rect 21361 21607 21419 21613
rect 21361 21604 21373 21607
rect 20220 21576 21373 21604
rect 20220 21564 20226 21576
rect 21361 21573 21373 21576
rect 21407 21573 21419 21607
rect 23198 21604 23204 21616
rect 21361 21567 21419 21573
rect 22480 21576 23204 21604
rect 22480 21548 22508 21576
rect 23198 21564 23204 21576
rect 23256 21564 23262 21616
rect 24026 21564 24032 21616
rect 24084 21564 24090 21616
rect 18877 21539 18935 21545
rect 18877 21536 18889 21539
rect 16546 21508 18889 21536
rect 18877 21505 18889 21508
rect 18923 21505 18935 21539
rect 18877 21499 18935 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 20717 21539 20775 21545
rect 20717 21536 20729 21539
rect 19935 21508 20729 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20717 21505 20729 21508
rect 20763 21505 20775 21539
rect 20717 21499 20775 21505
rect 22002 21496 22008 21548
rect 22060 21536 22066 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22060 21508 22385 21536
rect 22060 21496 22066 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22462 21496 22468 21548
rect 22520 21496 22526 21548
rect 23014 21496 23020 21548
rect 23072 21536 23078 21548
rect 23293 21539 23351 21545
rect 23293 21536 23305 21539
rect 23072 21508 23305 21536
rect 23072 21496 23078 21508
rect 23293 21505 23305 21508
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 9677 21471 9735 21477
rect 9677 21468 9689 21471
rect 8904 21440 9689 21468
rect 8904 21428 8910 21440
rect 9677 21437 9689 21440
rect 9723 21437 9735 21471
rect 9677 21431 9735 21437
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21437 9827 21471
rect 9769 21431 9827 21437
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21437 11115 21471
rect 11057 21431 11115 21437
rect 13357 21471 13415 21477
rect 13357 21437 13369 21471
rect 13403 21468 13415 21471
rect 14090 21468 14096 21480
rect 13403 21440 14096 21468
rect 13403 21437 13415 21440
rect 13357 21431 13415 21437
rect 9306 21360 9312 21412
rect 9364 21400 9370 21412
rect 9784 21400 9812 21431
rect 14090 21428 14096 21440
rect 14148 21428 14154 21480
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21468 14887 21471
rect 15102 21468 15108 21480
rect 14875 21440 15108 21468
rect 14875 21437 14887 21440
rect 14829 21431 14887 21437
rect 15102 21428 15108 21440
rect 15160 21428 15166 21480
rect 19978 21428 19984 21480
rect 20036 21468 20042 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 20036 21440 20085 21468
rect 20036 21428 20042 21440
rect 20073 21437 20085 21440
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 23569 21471 23627 21477
rect 22695 21440 23060 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 9364 21372 9812 21400
rect 9364 21360 9370 21372
rect 10778 21360 10784 21412
rect 10836 21400 10842 21412
rect 10836 21372 12434 21400
rect 10836 21360 10842 21372
rect 7742 21332 7748 21344
rect 7024 21304 7748 21332
rect 7742 21292 7748 21304
rect 7800 21292 7806 21344
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 8662 21332 8668 21344
rect 8352 21304 8668 21332
rect 8352 21292 8358 21304
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 9217 21335 9275 21341
rect 9217 21301 9229 21335
rect 9263 21332 9275 21335
rect 10962 21332 10968 21344
rect 9263 21304 10968 21332
rect 9263 21301 9275 21304
rect 9217 21295 9275 21301
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 12406 21332 12434 21372
rect 15470 21360 15476 21412
rect 15528 21400 15534 21412
rect 20990 21400 20996 21412
rect 15528 21372 20996 21400
rect 15528 21360 15534 21372
rect 20990 21360 20996 21372
rect 21048 21360 21054 21412
rect 21637 21403 21695 21409
rect 21637 21369 21649 21403
rect 21683 21400 21695 21403
rect 22278 21400 22284 21412
rect 21683 21372 22284 21400
rect 21683 21369 21695 21372
rect 21637 21363 21695 21369
rect 22278 21360 22284 21372
rect 22336 21400 22342 21412
rect 22462 21400 22468 21412
rect 22336 21372 22468 21400
rect 22336 21360 22342 21372
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 13998 21332 14004 21344
rect 12406 21304 14004 21332
rect 13998 21292 14004 21304
rect 14056 21292 14062 21344
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 15749 21335 15807 21341
rect 15749 21332 15761 21335
rect 15344 21304 15761 21332
rect 15344 21292 15350 21304
rect 15749 21301 15761 21304
rect 15795 21301 15807 21335
rect 15749 21295 15807 21301
rect 18690 21292 18696 21344
rect 18748 21292 18754 21344
rect 19518 21292 19524 21344
rect 19576 21292 19582 21344
rect 21910 21292 21916 21344
rect 21968 21332 21974 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21968 21304 22017 21332
rect 21968 21292 21974 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 23032 21332 23060 21440
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 25406 21468 25412 21480
rect 23615 21440 25412 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 25406 21428 25412 21440
rect 25464 21428 25470 21480
rect 23566 21332 23572 21344
rect 23032 21304 23572 21332
rect 22005 21295 22063 21301
rect 23566 21292 23572 21304
rect 23624 21292 23630 21344
rect 24026 21292 24032 21344
rect 24084 21332 24090 21344
rect 25317 21335 25375 21341
rect 25317 21332 25329 21335
rect 24084 21304 25329 21332
rect 24084 21292 24090 21304
rect 25317 21301 25329 21304
rect 25363 21301 25375 21335
rect 25317 21295 25375 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 8478 21088 8484 21140
rect 8536 21128 8542 21140
rect 12342 21128 12348 21140
rect 8536 21100 12348 21128
rect 8536 21088 8542 21100
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 12437 21131 12495 21137
rect 12437 21097 12449 21131
rect 12483 21128 12495 21131
rect 13354 21128 13360 21140
rect 12483 21100 13360 21128
rect 12483 21097 12495 21100
rect 12437 21091 12495 21097
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 16206 21088 16212 21140
rect 16264 21128 16270 21140
rect 16945 21131 17003 21137
rect 16945 21128 16957 21131
rect 16264 21100 16957 21128
rect 16264 21088 16270 21100
rect 16945 21097 16957 21100
rect 16991 21097 17003 21131
rect 16945 21091 17003 21097
rect 18690 21088 18696 21140
rect 18748 21128 18754 21140
rect 24762 21128 24768 21140
rect 18748 21100 24768 21128
rect 18748 21088 18754 21100
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 19429 21063 19487 21069
rect 19429 21029 19441 21063
rect 19475 21060 19487 21063
rect 20070 21060 20076 21072
rect 19475 21032 20076 21060
rect 19475 21029 19487 21032
rect 19429 21023 19487 21029
rect 20070 21020 20076 21032
rect 20128 21020 20134 21072
rect 20809 21063 20867 21069
rect 20809 21029 20821 21063
rect 20855 21060 20867 21063
rect 24581 21063 24639 21069
rect 20855 21032 22692 21060
rect 20855 21029 20867 21032
rect 20809 21023 20867 21029
rect 9950 20952 9956 21004
rect 10008 20952 10014 21004
rect 10962 20952 10968 21004
rect 11020 20992 11026 21004
rect 12618 20992 12624 21004
rect 11020 20964 12624 20992
rect 11020 20952 11026 20964
rect 12618 20952 12624 20964
rect 12676 20952 12682 21004
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20992 15255 20995
rect 16758 20992 16764 21004
rect 15243 20964 16764 20992
rect 15243 20961 15255 20964
rect 15197 20955 15255 20961
rect 16758 20952 16764 20964
rect 16816 20952 16822 21004
rect 19610 20952 19616 21004
rect 19668 20992 19674 21004
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19668 20964 19993 20992
rect 19668 20952 19674 20964
rect 19981 20961 19993 20964
rect 20027 20961 20039 20995
rect 19981 20955 20039 20961
rect 22002 20952 22008 21004
rect 22060 20952 22066 21004
rect 10686 20884 10692 20936
rect 10744 20884 10750 20936
rect 19794 20884 19800 20936
rect 19852 20924 19858 20936
rect 20441 20927 20499 20933
rect 20441 20924 20453 20927
rect 19852 20896 20453 20924
rect 19852 20884 19858 20896
rect 20441 20893 20453 20896
rect 20487 20893 20499 20927
rect 20441 20887 20499 20893
rect 20990 20884 20996 20936
rect 21048 20884 21054 20936
rect 22664 20933 22692 21032
rect 24581 21029 24593 21063
rect 24627 21060 24639 21063
rect 25038 21060 25044 21072
rect 24627 21032 25044 21060
rect 24627 21029 24639 21032
rect 24581 21023 24639 21029
rect 25038 21020 25044 21032
rect 25096 21020 25102 21072
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 24964 20964 25145 20992
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 24210 20884 24216 20936
rect 24268 20924 24274 20936
rect 24964 20924 24992 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 24268 20896 24992 20924
rect 25041 20927 25099 20933
rect 24268 20884 24274 20896
rect 25041 20893 25053 20927
rect 25087 20924 25099 20927
rect 25498 20924 25504 20936
rect 25087 20896 25504 20924
rect 25087 20893 25099 20896
rect 25041 20887 25099 20893
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 8570 20816 8576 20868
rect 8628 20856 8634 20868
rect 9217 20859 9275 20865
rect 9217 20856 9229 20859
rect 8628 20828 9229 20856
rect 8628 20816 8634 20828
rect 9217 20825 9229 20828
rect 9263 20825 9275 20859
rect 9217 20819 9275 20825
rect 10870 20816 10876 20868
rect 10928 20856 10934 20868
rect 10965 20859 11023 20865
rect 10965 20856 10977 20859
rect 10928 20828 10977 20856
rect 10928 20816 10934 20828
rect 10965 20825 10977 20828
rect 11011 20825 11023 20859
rect 15473 20859 15531 20865
rect 12190 20828 12848 20856
rect 10965 20819 11023 20825
rect 8846 20748 8852 20800
rect 8904 20788 8910 20800
rect 12820 20797 12848 20828
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 15746 20856 15752 20868
rect 15519 20828 15752 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 15746 20816 15752 20828
rect 15804 20816 15810 20868
rect 16698 20828 17264 20856
rect 9033 20791 9091 20797
rect 9033 20788 9045 20791
rect 8904 20760 9045 20788
rect 8904 20748 8910 20760
rect 9033 20757 9045 20760
rect 9079 20757 9091 20791
rect 9033 20751 9091 20757
rect 12805 20791 12863 20797
rect 12805 20757 12817 20791
rect 12851 20788 12863 20791
rect 14550 20788 14556 20800
rect 12851 20760 14556 20788
rect 12851 20757 12863 20760
rect 12805 20751 12863 20757
rect 14550 20748 14556 20760
rect 14608 20788 14614 20800
rect 14645 20791 14703 20797
rect 14645 20788 14657 20791
rect 14608 20760 14657 20788
rect 14608 20748 14614 20760
rect 14645 20757 14657 20760
rect 14691 20788 14703 20791
rect 15654 20788 15660 20800
rect 14691 20760 15660 20788
rect 14691 20757 14703 20760
rect 14645 20751 14703 20757
rect 15654 20748 15660 20760
rect 15712 20788 15718 20800
rect 16776 20788 16804 20828
rect 17236 20800 17264 20828
rect 19242 20816 19248 20868
rect 19300 20856 19306 20868
rect 19889 20859 19947 20865
rect 19889 20856 19901 20859
rect 19300 20828 19901 20856
rect 19300 20816 19306 20828
rect 19889 20825 19901 20828
rect 19935 20856 19947 20859
rect 21269 20859 21327 20865
rect 21269 20856 21281 20859
rect 19935 20828 21281 20856
rect 19935 20825 19947 20828
rect 19889 20819 19947 20825
rect 21269 20825 21281 20828
rect 21315 20825 21327 20859
rect 21269 20819 21327 20825
rect 24946 20816 24952 20868
rect 25004 20856 25010 20868
rect 25314 20856 25320 20868
rect 25004 20828 25320 20856
rect 25004 20816 25010 20828
rect 25314 20816 25320 20828
rect 25372 20816 25378 20868
rect 15712 20760 16804 20788
rect 15712 20748 15718 20760
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 17313 20791 17371 20797
rect 17313 20788 17325 20791
rect 17276 20760 17325 20788
rect 17276 20748 17282 20760
rect 17313 20757 17325 20760
rect 17359 20788 17371 20791
rect 17494 20788 17500 20800
rect 17359 20760 17500 20788
rect 17359 20757 17371 20760
rect 17313 20751 17371 20757
rect 17494 20748 17500 20760
rect 17552 20788 17558 20800
rect 18782 20788 18788 20800
rect 17552 20760 18788 20788
rect 17552 20748 17558 20760
rect 18782 20748 18788 20760
rect 18840 20748 18846 20800
rect 21450 20748 21456 20800
rect 21508 20748 21514 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10413 20587 10471 20593
rect 10413 20584 10425 20587
rect 10192 20556 10425 20584
rect 10192 20544 10198 20556
rect 10413 20553 10425 20556
rect 10459 20553 10471 20587
rect 10413 20547 10471 20553
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 12526 20584 12532 20596
rect 10827 20556 12532 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 15473 20587 15531 20593
rect 15473 20553 15485 20587
rect 15519 20584 15531 20587
rect 15930 20584 15936 20596
rect 15519 20556 15936 20584
rect 15519 20553 15531 20556
rect 15473 20547 15531 20553
rect 15930 20544 15936 20556
rect 15988 20544 15994 20596
rect 19426 20584 19432 20596
rect 16868 20556 19432 20584
rect 8021 20519 8079 20525
rect 8021 20485 8033 20519
rect 8067 20516 8079 20519
rect 8294 20516 8300 20528
rect 8067 20488 8300 20516
rect 8067 20485 8079 20488
rect 8021 20479 8079 20485
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 8570 20476 8576 20528
rect 8628 20476 8634 20528
rect 14550 20516 14556 20528
rect 14214 20488 14556 20516
rect 14550 20476 14556 20488
rect 14608 20476 14614 20528
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 12492 20420 12725 20448
rect 12492 20408 12498 20420
rect 12713 20417 12725 20420
rect 12759 20417 12771 20451
rect 12713 20411 12771 20417
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 16868 20457 16896 20556
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 20901 20587 20959 20593
rect 20901 20553 20913 20587
rect 20947 20584 20959 20587
rect 21450 20584 21456 20596
rect 20947 20556 21456 20584
rect 20947 20553 20959 20556
rect 20901 20547 20959 20553
rect 21450 20544 21456 20556
rect 21508 20544 21514 20596
rect 22830 20544 22836 20596
rect 22888 20584 22894 20596
rect 22925 20587 22983 20593
rect 22925 20584 22937 20587
rect 22888 20556 22937 20584
rect 22888 20544 22894 20556
rect 22925 20553 22937 20556
rect 22971 20553 22983 20587
rect 22925 20547 22983 20553
rect 24026 20544 24032 20596
rect 24084 20544 24090 20596
rect 25317 20587 25375 20593
rect 25317 20553 25329 20587
rect 25363 20584 25375 20587
rect 25406 20584 25412 20596
rect 25363 20556 25412 20584
rect 25363 20553 25375 20556
rect 25317 20547 25375 20553
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 17126 20476 17132 20528
rect 17184 20476 17190 20528
rect 18782 20516 18788 20528
rect 18354 20488 18788 20516
rect 18782 20476 18788 20488
rect 18840 20476 18846 20528
rect 18874 20476 18880 20528
rect 18932 20516 18938 20528
rect 18932 20488 20852 20516
rect 18932 20476 18938 20488
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 19150 20408 19156 20460
rect 19208 20448 19214 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 19208 20420 19257 20448
rect 19208 20408 19214 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 20346 20448 20352 20460
rect 19935 20420 20352 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20824 20457 20852 20488
rect 21174 20476 21180 20528
rect 21232 20516 21238 20528
rect 24044 20516 24072 20544
rect 21232 20488 22324 20516
rect 24044 20488 24334 20516
rect 21232 20476 21238 20488
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20448 20867 20451
rect 21453 20451 21511 20457
rect 21453 20448 21465 20451
rect 20855 20420 21465 20448
rect 20855 20417 20867 20420
rect 20809 20411 20867 20417
rect 21453 20417 21465 20420
rect 21499 20417 21511 20451
rect 21453 20411 21511 20417
rect 22186 20408 22192 20460
rect 22244 20408 22250 20460
rect 22296 20448 22324 20488
rect 23109 20451 23167 20457
rect 23109 20448 23121 20451
rect 22296 20420 23121 20448
rect 23109 20417 23121 20420
rect 23155 20417 23167 20451
rect 23109 20411 23167 20417
rect 7742 20340 7748 20392
rect 7800 20340 7806 20392
rect 8386 20340 8392 20392
rect 8444 20380 8450 20392
rect 9306 20380 9312 20392
rect 8444 20352 9312 20380
rect 8444 20340 8450 20352
rect 9306 20340 9312 20352
rect 9364 20380 9370 20392
rect 9364 20352 9720 20380
rect 9364 20340 9370 20352
rect 9692 20312 9720 20352
rect 9766 20340 9772 20392
rect 9824 20340 9830 20392
rect 10226 20340 10232 20392
rect 10284 20380 10290 20392
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10284 20352 10885 20380
rect 10284 20340 10290 20352
rect 10873 20349 10885 20352
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13446 20380 13452 20392
rect 13035 20352 13452 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 10980 20312 11008 20343
rect 13446 20340 13452 20352
rect 13504 20380 13510 20392
rect 15102 20380 15108 20392
rect 13504 20352 15108 20380
rect 13504 20340 13510 20352
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 15565 20383 15623 20389
rect 15565 20349 15577 20383
rect 15611 20349 15623 20383
rect 15565 20343 15623 20349
rect 15580 20312 15608 20343
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 18598 20380 18604 20392
rect 17552 20352 18604 20380
rect 17552 20340 17558 20352
rect 18598 20340 18604 20352
rect 18656 20340 18662 20392
rect 21085 20383 21143 20389
rect 21085 20349 21097 20383
rect 21131 20380 21143 20383
rect 22554 20380 22560 20392
rect 21131 20352 22560 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 23566 20340 23572 20392
rect 23624 20340 23630 20392
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 25130 20380 25136 20392
rect 23891 20352 25136 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 19150 20312 19156 20324
rect 9692 20284 11008 20312
rect 14476 20284 15608 20312
rect 18156 20284 19156 20312
rect 14476 20256 14504 20284
rect 10134 20204 10140 20256
rect 10192 20204 10198 20256
rect 14458 20204 14464 20256
rect 14516 20204 14522 20256
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 18156 20244 18184 20284
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 20441 20315 20499 20321
rect 20441 20281 20453 20315
rect 20487 20312 20499 20315
rect 21542 20312 21548 20324
rect 20487 20284 21548 20312
rect 20487 20281 20499 20284
rect 20441 20275 20499 20281
rect 21542 20272 21548 20284
rect 21600 20272 21606 20324
rect 22005 20315 22063 20321
rect 22005 20281 22017 20315
rect 22051 20312 22063 20315
rect 22051 20284 23060 20312
rect 22051 20281 22063 20284
rect 22005 20275 22063 20281
rect 15059 20216 18184 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 19058 20204 19064 20256
rect 19116 20204 19122 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19392 20216 19717 20244
rect 19392 20204 19398 20216
rect 19705 20213 19717 20216
rect 19751 20213 19763 20247
rect 19705 20207 19763 20213
rect 22462 20204 22468 20256
rect 22520 20204 22526 20256
rect 23032 20244 23060 20284
rect 23934 20244 23940 20256
rect 23032 20216 23940 20244
rect 23934 20204 23940 20216
rect 23992 20204 23998 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 8481 20043 8539 20049
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 8570 20040 8576 20052
rect 8527 20012 8576 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 8570 20000 8576 20012
rect 8628 20000 8634 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 14182 20040 14188 20052
rect 11379 20012 14188 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 14540 20043 14598 20049
rect 14540 20009 14552 20043
rect 14586 20040 14598 20043
rect 15562 20040 15568 20052
rect 14586 20012 15568 20040
rect 14586 20009 14598 20012
rect 14540 20003 14598 20009
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 15746 20000 15752 20052
rect 15804 20040 15810 20052
rect 16025 20043 16083 20049
rect 16025 20040 16037 20043
rect 15804 20012 16037 20040
rect 15804 20000 15810 20012
rect 16025 20009 16037 20012
rect 16071 20009 16083 20043
rect 16025 20003 16083 20009
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20040 17003 20043
rect 17218 20040 17224 20052
rect 16991 20012 17224 20040
rect 16991 20009 17003 20012
rect 16945 20003 17003 20009
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 22186 20040 22192 20052
rect 18156 20012 22192 20040
rect 15838 19932 15844 19984
rect 15896 19972 15902 19984
rect 17034 19972 17040 19984
rect 15896 19944 17040 19972
rect 15896 19932 15902 19944
rect 17034 19932 17040 19944
rect 17092 19932 17098 19984
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 17184 19944 18092 19972
rect 17184 19932 17190 19944
rect 10686 19904 10692 19916
rect 9140 19876 10692 19904
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 9030 19836 9036 19848
rect 7800 19808 9036 19836
rect 7800 19796 7806 19808
rect 9030 19796 9036 19808
rect 9088 19836 9094 19848
rect 9140 19845 9168 19876
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 12492 19876 14289 19904
rect 12492 19864 12498 19876
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 14277 19867 14335 19873
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 17218 19904 17224 19916
rect 14700 19876 17224 19904
rect 14700 19864 14706 19876
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 18064 19913 18092 19944
rect 17957 19907 18015 19913
rect 17957 19904 17969 19907
rect 17920 19876 17969 19904
rect 17920 19864 17926 19876
rect 17957 19873 17969 19876
rect 18003 19873 18015 19907
rect 17957 19867 18015 19873
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 9088 19808 9137 19836
rect 9088 19796 9094 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 15654 19796 15660 19848
rect 15712 19796 15718 19848
rect 16669 19839 16727 19845
rect 16669 19836 16681 19839
rect 15856 19808 16681 19836
rect 8662 19728 8668 19780
rect 8720 19768 8726 19780
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 8720 19740 9413 19768
rect 8720 19728 8726 19740
rect 9401 19737 9413 19740
rect 9447 19768 9459 19771
rect 9490 19768 9496 19780
rect 9447 19740 9496 19768
rect 9447 19737 9459 19740
rect 9401 19731 9459 19737
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 10134 19728 10140 19780
rect 10192 19728 10198 19780
rect 11606 19728 11612 19780
rect 11664 19768 11670 19780
rect 11793 19771 11851 19777
rect 11793 19768 11805 19771
rect 11664 19740 11805 19768
rect 11664 19728 11670 19740
rect 11793 19737 11805 19740
rect 11839 19737 11851 19771
rect 11793 19731 11851 19737
rect 10870 19660 10876 19712
rect 10928 19660 10934 19712
rect 11698 19660 11704 19712
rect 11756 19660 11762 19712
rect 12526 19660 12532 19712
rect 12584 19700 12590 19712
rect 15856 19700 15884 19808
rect 16669 19805 16681 19808
rect 16715 19805 16727 19839
rect 18156 19836 18184 20012
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 23845 20043 23903 20049
rect 23845 20040 23857 20043
rect 23716 20012 23857 20040
rect 23716 20000 23722 20012
rect 23845 20009 23857 20012
rect 23891 20040 23903 20043
rect 24210 20040 24216 20052
rect 23891 20012 24216 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 24210 20000 24216 20012
rect 24268 20000 24274 20052
rect 25314 20000 25320 20052
rect 25372 20000 25378 20052
rect 21634 19932 21640 19984
rect 21692 19972 21698 19984
rect 21692 19944 22219 19972
rect 21692 19932 21698 19944
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 20162 19904 20168 19916
rect 19935 19876 20168 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 20162 19864 20168 19876
rect 20220 19904 20226 19916
rect 22097 19907 22155 19913
rect 22097 19904 22109 19907
rect 20220 19876 22109 19904
rect 20220 19864 20226 19876
rect 22097 19873 22109 19876
rect 22143 19873 22155 19907
rect 22191 19904 22219 19944
rect 22373 19907 22431 19913
rect 22373 19904 22385 19907
rect 22191 19876 22385 19904
rect 22097 19867 22155 19873
rect 22373 19873 22385 19876
rect 22419 19873 22431 19907
rect 22373 19867 22431 19873
rect 16669 19799 16727 19805
rect 16960 19808 18184 19836
rect 18877 19839 18935 19845
rect 16960 19768 16988 19808
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19702 19836 19708 19848
rect 18923 19808 19708 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19702 19796 19708 19808
rect 19760 19796 19766 19848
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 16500 19740 16988 19768
rect 16500 19709 16528 19740
rect 17034 19728 17040 19780
rect 17092 19768 17098 19780
rect 17865 19771 17923 19777
rect 17865 19768 17877 19771
rect 17092 19740 17877 19768
rect 17092 19728 17098 19740
rect 17865 19737 17877 19740
rect 17911 19737 17923 19771
rect 19794 19768 19800 19780
rect 17865 19731 17923 19737
rect 18616 19740 19800 19768
rect 12584 19672 15884 19700
rect 16485 19703 16543 19709
rect 12584 19660 12590 19672
rect 16485 19669 16497 19703
rect 16531 19669 16543 19703
rect 16485 19663 16543 19669
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 18616 19700 18644 19740
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 19886 19728 19892 19780
rect 19944 19768 19950 19780
rect 20165 19771 20223 19777
rect 20165 19768 20177 19771
rect 19944 19740 20177 19768
rect 19944 19728 19950 19740
rect 20165 19737 20177 19740
rect 20211 19737 20223 19771
rect 20165 19731 20223 19737
rect 20548 19740 20654 19768
rect 17543 19672 18644 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 18782 19660 18788 19712
rect 18840 19700 18846 19712
rect 19521 19703 19579 19709
rect 19521 19700 19533 19703
rect 18840 19672 19533 19700
rect 18840 19660 18846 19672
rect 19521 19669 19533 19672
rect 19567 19700 19579 19703
rect 20548 19700 20576 19740
rect 22462 19728 22468 19780
rect 22520 19768 22526 19780
rect 22520 19740 22862 19768
rect 22520 19728 22526 19740
rect 22480 19700 22508 19728
rect 19567 19672 22508 19700
rect 22756 19700 22784 19740
rect 24121 19703 24179 19709
rect 24121 19700 24133 19703
rect 22756 19672 24133 19700
rect 19567 19669 19579 19672
rect 19521 19663 19579 19669
rect 24121 19669 24133 19672
rect 24167 19700 24179 19703
rect 24210 19700 24216 19712
rect 24167 19672 24216 19700
rect 24167 19669 24179 19672
rect 24121 19663 24179 19669
rect 24210 19660 24216 19672
rect 24268 19660 24274 19712
rect 24578 19660 24584 19712
rect 24636 19660 24642 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 10192 19468 10977 19496
rect 10192 19456 10198 19468
rect 10965 19465 10977 19468
rect 11011 19496 11023 19499
rect 11146 19496 11152 19508
rect 11011 19468 11152 19496
rect 11011 19465 11023 19468
rect 10965 19459 11023 19465
rect 11146 19456 11152 19468
rect 11204 19456 11210 19508
rect 11698 19456 11704 19508
rect 11756 19456 11762 19508
rect 11790 19456 11796 19508
rect 11848 19496 11854 19508
rect 15013 19499 15071 19505
rect 11848 19468 14136 19496
rect 11848 19456 11854 19468
rect 8570 19428 8576 19440
rect 8050 19400 8576 19428
rect 8570 19388 8576 19400
rect 8628 19388 8634 19440
rect 9125 19431 9183 19437
rect 9125 19397 9137 19431
rect 9171 19428 9183 19431
rect 9214 19428 9220 19440
rect 9171 19400 9220 19428
rect 9171 19397 9183 19400
rect 9125 19391 9183 19397
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 14108 19428 14136 19468
rect 15013 19465 15025 19499
rect 15059 19496 15071 19499
rect 15470 19496 15476 19508
rect 15059 19468 15476 19496
rect 15059 19465 15071 19468
rect 15013 19459 15071 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 14108 19400 15240 19428
rect 10134 19360 10140 19372
rect 9232 19332 10140 19360
rect 6546 19252 6552 19304
rect 6604 19252 6610 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 6914 19292 6920 19304
rect 6871 19264 6920 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 9232 19301 9260 19332
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12529 19363 12587 19369
rect 12529 19360 12541 19363
rect 12492 19332 12541 19360
rect 12492 19320 12498 19332
rect 12529 19329 12541 19332
rect 12575 19329 12587 19363
rect 14550 19360 14556 19372
rect 13938 19332 14556 19360
rect 12529 19323 12587 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 15212 19369 15240 19400
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19360 16175 19363
rect 16390 19360 16396 19372
rect 16163 19332 16396 19360
rect 16163 19329 16175 19332
rect 16117 19323 16175 19329
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 16868 19360 16896 19459
rect 17218 19456 17224 19508
rect 17276 19456 17282 19508
rect 17310 19456 17316 19508
rect 17368 19456 17374 19508
rect 17402 19456 17408 19508
rect 17460 19496 17466 19508
rect 18690 19496 18696 19508
rect 17460 19468 18696 19496
rect 17460 19456 17466 19468
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 18969 19499 19027 19505
rect 18969 19465 18981 19499
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 18984 19428 19012 19459
rect 19518 19456 19524 19508
rect 19576 19496 19582 19508
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19576 19468 20453 19496
rect 19576 19456 19582 19468
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 20714 19496 20720 19508
rect 20579 19468 20720 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 22649 19499 22707 19505
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 23474 19496 23480 19508
rect 22695 19468 23480 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 23474 19456 23480 19468
rect 23532 19456 23538 19508
rect 25130 19456 25136 19508
rect 25188 19456 25194 19508
rect 22186 19428 22192 19440
rect 18984 19400 22192 19428
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 23566 19428 23572 19440
rect 23400 19400 23572 19428
rect 16868 19332 19104 19360
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 14458 19292 14464 19304
rect 12851 19264 14464 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 8478 19184 8484 19236
rect 8536 19224 8542 19236
rect 9324 19224 9352 19255
rect 14458 19252 14464 19264
rect 14516 19252 14522 19304
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 8536 19196 9352 19224
rect 8536 19184 8542 19196
rect 9398 19184 9404 19236
rect 9456 19224 9462 19236
rect 10962 19224 10968 19236
rect 9456 19196 10968 19224
rect 9456 19184 9462 19196
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 15746 19184 15752 19236
rect 15804 19224 15810 19236
rect 17420 19224 17448 19255
rect 17770 19252 17776 19304
rect 17828 19292 17834 19304
rect 17865 19295 17923 19301
rect 17865 19292 17877 19295
rect 17828 19264 17877 19292
rect 17828 19252 17834 19264
rect 17865 19261 17877 19264
rect 17911 19261 17923 19295
rect 19076 19292 19104 19332
rect 19150 19320 19156 19372
rect 19208 19320 19214 19372
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 20346 19360 20352 19372
rect 19944 19332 20352 19360
rect 19944 19320 19950 19332
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 23400 19369 23428 19400
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 23658 19388 23664 19440
rect 23716 19388 23722 19440
rect 24210 19388 24216 19440
rect 24268 19388 24274 19440
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 21315 19332 22569 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 19978 19292 19984 19304
rect 19076 19264 19984 19292
rect 17865 19255 17923 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20625 19295 20683 19301
rect 20625 19261 20637 19295
rect 20671 19292 20683 19295
rect 21634 19292 21640 19304
rect 20671 19264 21640 19292
rect 20671 19261 20683 19264
rect 20625 19255 20683 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 22738 19252 22744 19304
rect 22796 19252 22802 19304
rect 15804 19196 17448 19224
rect 15804 19184 15810 19196
rect 17586 19184 17592 19236
rect 17644 19224 17650 19236
rect 18049 19227 18107 19233
rect 18049 19224 18061 19227
rect 17644 19196 18061 19224
rect 17644 19184 17650 19196
rect 18049 19193 18061 19196
rect 18095 19224 18107 19227
rect 21174 19224 21180 19236
rect 18095 19196 21180 19224
rect 18095 19193 18107 19196
rect 18049 19187 18107 19193
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 21450 19184 21456 19236
rect 21508 19224 21514 19236
rect 22189 19227 22247 19233
rect 22189 19224 22201 19227
rect 21508 19196 22201 19224
rect 21508 19184 21514 19196
rect 22189 19193 22201 19196
rect 22235 19193 22247 19227
rect 22189 19187 22247 19193
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 9306 19156 9312 19168
rect 8352 19128 9312 19156
rect 8352 19116 8358 19128
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 10318 19116 10324 19168
rect 10376 19156 10382 19168
rect 11149 19159 11207 19165
rect 11149 19156 11161 19159
rect 10376 19128 11161 19156
rect 10376 19116 10382 19128
rect 11149 19125 11161 19128
rect 11195 19156 11207 19159
rect 11606 19156 11612 19168
rect 11195 19128 11612 19156
rect 11195 19125 11207 19128
rect 11149 19119 11207 19125
rect 11606 19116 11612 19128
rect 11664 19116 11670 19168
rect 14090 19116 14096 19168
rect 14148 19156 14154 19168
rect 14277 19159 14335 19165
rect 14277 19156 14289 19159
rect 14148 19128 14289 19156
rect 14148 19116 14154 19128
rect 14277 19125 14289 19128
rect 14323 19125 14335 19159
rect 14277 19119 14335 19125
rect 14550 19116 14556 19168
rect 14608 19116 14614 19168
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15160 19128 15945 19156
rect 15160 19116 15166 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 18782 19116 18788 19168
rect 18840 19156 18846 19168
rect 20073 19159 20131 19165
rect 20073 19156 20085 19159
rect 18840 19128 20085 19156
rect 18840 19116 18846 19128
rect 20073 19125 20085 19128
rect 20119 19125 20131 19159
rect 20073 19119 20131 19125
rect 21818 19116 21824 19168
rect 21876 19116 21882 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 8665 18955 8723 18961
rect 8665 18952 8677 18955
rect 8628 18924 8677 18952
rect 8628 18912 8634 18924
rect 8665 18921 8677 18924
rect 8711 18921 8723 18955
rect 8665 18915 8723 18921
rect 10042 18912 10048 18964
rect 10100 18912 10106 18964
rect 11149 18955 11207 18961
rect 11149 18952 11161 18955
rect 10612 18924 11161 18952
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 8294 18816 8300 18828
rect 6963 18788 8300 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 10612 18825 10640 18924
rect 11149 18921 11161 18924
rect 11195 18952 11207 18955
rect 11238 18952 11244 18964
rect 11195 18924 11244 18952
rect 11195 18921 11207 18924
rect 11149 18915 11207 18921
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 11517 18955 11575 18961
rect 11517 18921 11529 18955
rect 11563 18952 11575 18955
rect 12526 18952 12532 18964
rect 11563 18924 12532 18952
rect 11563 18921 11575 18924
rect 11517 18915 11575 18921
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 12710 18912 12716 18964
rect 12768 18912 12774 18964
rect 17586 18952 17592 18964
rect 17328 18924 17592 18952
rect 10962 18844 10968 18896
rect 11020 18884 11026 18896
rect 11020 18856 13308 18884
rect 11020 18844 11026 18856
rect 10597 18819 10655 18825
rect 10597 18785 10609 18819
rect 10643 18785 10655 18819
rect 10597 18779 10655 18785
rect 10870 18776 10876 18828
rect 10928 18816 10934 18828
rect 13280 18825 13308 18856
rect 12069 18819 12127 18825
rect 12069 18816 12081 18819
rect 10928 18788 12081 18816
rect 10928 18776 10934 18788
rect 12069 18785 12081 18788
rect 12115 18785 12127 18819
rect 12069 18779 12127 18785
rect 13265 18819 13323 18825
rect 13265 18785 13277 18819
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 17328 18825 17356 18924
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 18141 18887 18199 18893
rect 18141 18853 18153 18887
rect 18187 18884 18199 18887
rect 21634 18884 21640 18896
rect 18187 18856 21640 18884
rect 18187 18853 18199 18856
rect 18141 18847 18199 18853
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 16724 18788 17325 18816
rect 16724 18776 16730 18788
rect 17313 18785 17325 18788
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18816 17555 18819
rect 17586 18816 17592 18828
rect 17543 18788 17592 18816
rect 17543 18785 17555 18788
rect 17497 18779 17555 18785
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 18598 18776 18604 18828
rect 18656 18816 18662 18828
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 18656 18788 18705 18816
rect 18656 18776 18662 18788
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 23382 18776 23388 18828
rect 23440 18816 23446 18828
rect 23477 18819 23535 18825
rect 23477 18816 23489 18819
rect 23440 18788 23489 18816
rect 23440 18776 23446 18788
rect 23477 18785 23489 18788
rect 23523 18785 23535 18819
rect 23477 18779 23535 18785
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 8570 18748 8576 18760
rect 8050 18720 8576 18748
rect 8570 18708 8576 18720
rect 8628 18748 8634 18760
rect 8754 18748 8760 18760
rect 8628 18720 8760 18748
rect 8628 18708 8634 18720
rect 8754 18708 8760 18720
rect 8812 18748 8818 18760
rect 9122 18748 9128 18760
rect 8812 18720 9128 18748
rect 8812 18708 8818 18720
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 13814 18748 13820 18760
rect 10551 18720 12434 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 11238 18680 11244 18692
rect 8352 18652 11244 18680
rect 8352 18640 8358 18652
rect 11238 18640 11244 18652
rect 11296 18640 11302 18692
rect 11977 18683 12035 18689
rect 11977 18649 11989 18683
rect 12023 18680 12035 18683
rect 12066 18680 12072 18692
rect 12023 18652 12072 18680
rect 12023 18649 12035 18652
rect 11977 18643 12035 18649
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 8389 18615 8447 18621
rect 8389 18581 8401 18615
rect 8435 18612 8447 18615
rect 8570 18612 8576 18624
rect 8435 18584 8576 18612
rect 8435 18581 8447 18584
rect 8389 18575 8447 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8846 18572 8852 18624
rect 8904 18612 8910 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 8904 18584 9689 18612
rect 8904 18572 8910 18584
rect 9677 18581 9689 18584
rect 9723 18612 9735 18615
rect 10413 18615 10471 18621
rect 10413 18612 10425 18615
rect 9723 18584 10425 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 10413 18581 10425 18584
rect 10459 18581 10471 18615
rect 10413 18575 10471 18581
rect 11422 18572 11428 18624
rect 11480 18612 11486 18624
rect 11885 18615 11943 18621
rect 11885 18612 11897 18615
rect 11480 18584 11897 18612
rect 11480 18572 11486 18584
rect 11885 18581 11897 18584
rect 11931 18581 11943 18615
rect 12406 18612 12434 18720
rect 12544 18720 13820 18748
rect 12544 18612 12572 18720
rect 13814 18708 13820 18720
rect 13872 18708 13878 18760
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18748 17279 18751
rect 17770 18748 17776 18760
rect 17267 18720 17776 18748
rect 17267 18717 17279 18720
rect 17221 18711 17279 18717
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 13081 18683 13139 18689
rect 13081 18680 13093 18683
rect 12676 18652 13093 18680
rect 12676 18640 12682 18652
rect 13081 18649 13093 18652
rect 13127 18649 13139 18683
rect 13081 18643 13139 18649
rect 18509 18683 18567 18689
rect 18509 18649 18521 18683
rect 18555 18680 18567 18683
rect 18966 18680 18972 18692
rect 18555 18652 18972 18680
rect 18555 18649 18567 18652
rect 18509 18643 18567 18649
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 21468 18680 21496 18711
rect 22186 18708 22192 18760
rect 22244 18708 22250 18760
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 24578 18748 24584 18760
rect 22879 18720 24584 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 24578 18708 24584 18720
rect 24636 18708 24642 18760
rect 25133 18751 25191 18757
rect 25133 18748 25145 18751
rect 24688 18720 25145 18748
rect 24394 18680 24400 18692
rect 21468 18652 24400 18680
rect 24394 18640 24400 18652
rect 24452 18640 24458 18692
rect 24486 18640 24492 18692
rect 24544 18680 24550 18692
rect 24688 18689 24716 18720
rect 25133 18717 25145 18720
rect 25179 18717 25191 18751
rect 25133 18711 25191 18717
rect 24673 18683 24731 18689
rect 24673 18680 24685 18683
rect 24544 18652 24685 18680
rect 24544 18640 24550 18652
rect 24673 18649 24685 18652
rect 24719 18649 24731 18683
rect 24673 18643 24731 18649
rect 24857 18683 24915 18689
rect 24857 18649 24869 18683
rect 24903 18680 24915 18683
rect 24946 18680 24952 18692
rect 24903 18652 24952 18680
rect 24903 18649 24915 18652
rect 24857 18643 24915 18649
rect 24946 18640 24952 18652
rect 25004 18640 25010 18692
rect 12406 18584 12572 18612
rect 11885 18575 11943 18581
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13173 18615 13231 18621
rect 13173 18612 13185 18615
rect 12860 18584 13185 18612
rect 12860 18572 12866 18584
rect 13173 18581 13185 18584
rect 13219 18581 13231 18615
rect 13173 18575 13231 18581
rect 13817 18615 13875 18621
rect 13817 18581 13829 18615
rect 13863 18612 13875 18615
rect 13906 18612 13912 18624
rect 13863 18584 13912 18612
rect 13863 18581 13875 18584
rect 13817 18575 13875 18581
rect 13906 18572 13912 18584
rect 13964 18572 13970 18624
rect 14274 18572 14280 18624
rect 14332 18572 14338 18624
rect 16853 18615 16911 18621
rect 16853 18581 16865 18615
rect 16899 18612 16911 18615
rect 17034 18612 17040 18624
rect 16899 18584 17040 18612
rect 16899 18581 16911 18584
rect 16853 18575 16911 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18380 18584 18613 18612
rect 18380 18572 18386 18584
rect 18601 18581 18613 18584
rect 18647 18581 18659 18615
rect 18601 18575 18659 18581
rect 19886 18572 19892 18624
rect 19944 18612 19950 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 19944 18584 21281 18612
rect 19944 18572 19950 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 22005 18615 22063 18621
rect 22005 18581 22017 18615
rect 22051 18612 22063 18615
rect 22094 18612 22100 18624
rect 22051 18584 22100 18612
rect 22051 18581 22063 18584
rect 22005 18575 22063 18581
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 9398 18368 9404 18420
rect 9456 18408 9462 18420
rect 9493 18411 9551 18417
rect 9493 18408 9505 18411
rect 9456 18380 9505 18408
rect 9456 18368 9462 18380
rect 9493 18377 9505 18380
rect 9539 18377 9551 18411
rect 9493 18371 9551 18377
rect 10413 18411 10471 18417
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 10778 18408 10784 18420
rect 10459 18380 10784 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 11057 18411 11115 18417
rect 11057 18377 11069 18411
rect 11103 18408 11115 18411
rect 11146 18408 11152 18420
rect 11103 18380 11152 18408
rect 11103 18377 11115 18380
rect 11057 18371 11115 18377
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 11238 18368 11244 18420
rect 11296 18408 11302 18420
rect 11514 18408 11520 18420
rect 11296 18380 11520 18408
rect 11296 18368 11302 18380
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 12492 18380 13216 18408
rect 12492 18368 12498 18380
rect 8021 18343 8079 18349
rect 8021 18309 8033 18343
rect 8067 18340 8079 18343
rect 8294 18340 8300 18352
rect 8067 18312 8300 18340
rect 8067 18309 8079 18312
rect 8021 18303 8079 18309
rect 8294 18300 8300 18312
rect 8352 18300 8358 18352
rect 8754 18300 8760 18352
rect 8812 18300 8818 18352
rect 9306 18300 9312 18352
rect 9364 18340 9370 18352
rect 13188 18349 13216 18380
rect 13814 18368 13820 18420
rect 13872 18368 13878 18420
rect 14185 18411 14243 18417
rect 14185 18377 14197 18411
rect 14231 18408 14243 18411
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14231 18380 14933 18408
rect 14231 18377 14243 18380
rect 14185 18371 14243 18377
rect 14921 18377 14933 18380
rect 14967 18408 14979 18411
rect 16850 18408 16856 18420
rect 14967 18380 16856 18408
rect 14967 18377 14979 18380
rect 14921 18371 14979 18377
rect 16850 18368 16856 18380
rect 16908 18408 16914 18420
rect 26142 18408 26148 18420
rect 16908 18380 26148 18408
rect 16908 18368 16914 18380
rect 26142 18368 26148 18380
rect 26200 18368 26206 18420
rect 13173 18343 13231 18349
rect 9364 18312 10548 18340
rect 9364 18300 9370 18312
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 6638 18164 6644 18216
rect 6696 18204 6702 18216
rect 7745 18207 7803 18213
rect 7745 18204 7757 18207
rect 6696 18176 7757 18204
rect 6696 18164 6702 18176
rect 7745 18173 7757 18176
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 7760 18068 7788 18167
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 10336 18204 10364 18235
rect 10520 18213 10548 18312
rect 13173 18309 13185 18343
rect 13219 18309 13231 18343
rect 18874 18340 18880 18352
rect 18354 18312 18880 18340
rect 13173 18303 13231 18309
rect 18874 18300 18880 18312
rect 18932 18300 18938 18352
rect 22370 18340 22376 18352
rect 21284 18312 22376 18340
rect 12434 18232 12440 18284
rect 12492 18232 12498 18284
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16816 18244 16865 18272
rect 16816 18232 16822 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 19978 18232 19984 18284
rect 20036 18232 20042 18284
rect 21284 18281 21312 18312
rect 22370 18300 22376 18312
rect 22428 18300 22434 18352
rect 23293 18343 23351 18349
rect 23293 18309 23305 18343
rect 23339 18340 23351 18343
rect 24854 18340 24860 18352
rect 23339 18312 24860 18340
rect 23339 18309 23351 18312
rect 23293 18303 23351 18309
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 8168 18176 10364 18204
rect 10505 18207 10563 18213
rect 8168 18164 8174 18176
rect 10505 18173 10517 18207
rect 10551 18173 10563 18207
rect 10505 18167 10563 18173
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 13964 18176 14289 18204
rect 13964 18164 13970 18176
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18173 14427 18207
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 14369 18167 14427 18173
rect 16868 18176 17141 18204
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 9582 18136 9588 18148
rect 9088 18108 9588 18136
rect 9088 18096 9094 18108
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 9953 18139 10011 18145
rect 9953 18105 9965 18139
rect 9999 18136 10011 18139
rect 11790 18136 11796 18148
rect 9999 18108 11796 18136
rect 9999 18105 10011 18108
rect 9953 18099 10011 18105
rect 11790 18096 11796 18108
rect 11848 18096 11854 18148
rect 9048 18068 9076 18096
rect 7760 18040 9076 18068
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 13722 18068 13728 18080
rect 9824 18040 13728 18068
rect 9824 18028 9830 18040
rect 13722 18028 13728 18040
rect 13780 18068 13786 18080
rect 14384 18068 14412 18167
rect 16868 18148 16896 18176
rect 17129 18173 17141 18176
rect 17175 18204 17187 18207
rect 17494 18204 17500 18216
rect 17175 18176 17500 18204
rect 17175 18173 17187 18176
rect 17129 18167 17187 18173
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 24670 18164 24676 18216
rect 24728 18164 24734 18216
rect 16850 18096 16856 18148
rect 16908 18096 16914 18148
rect 19797 18139 19855 18145
rect 19797 18105 19809 18139
rect 19843 18136 19855 18139
rect 25222 18136 25228 18148
rect 19843 18108 25228 18136
rect 19843 18105 19855 18108
rect 19797 18099 19855 18105
rect 25222 18096 25228 18108
rect 25280 18096 25286 18148
rect 13780 18040 14412 18068
rect 13780 18028 13786 18040
rect 18598 18028 18604 18080
rect 18656 18028 18662 18080
rect 18874 18028 18880 18080
rect 18932 18028 18938 18080
rect 21082 18028 21088 18080
rect 21140 18028 21146 18080
rect 22738 18028 22744 18080
rect 22796 18068 22802 18080
rect 24118 18068 24124 18080
rect 22796 18040 24124 18068
rect 22796 18028 22802 18040
rect 24118 18028 24124 18040
rect 24176 18028 24182 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7708 17836 7849 17864
rect 7708 17824 7714 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 13906 17864 13912 17876
rect 12124 17836 13912 17864
rect 12124 17824 12130 17836
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18417 17867 18475 17873
rect 18417 17864 18429 17867
rect 18012 17836 18429 17864
rect 18012 17824 18018 17836
rect 18417 17833 18429 17836
rect 18463 17833 18475 17867
rect 18417 17827 18475 17833
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 18874 17864 18880 17876
rect 18748 17836 18880 17864
rect 18748 17824 18754 17836
rect 18874 17824 18880 17836
rect 18932 17864 18938 17876
rect 18969 17867 19027 17873
rect 18969 17864 18981 17867
rect 18932 17836 18981 17864
rect 18932 17824 18938 17836
rect 18969 17833 18981 17836
rect 19015 17833 19027 17867
rect 18969 17827 19027 17833
rect 21637 17867 21695 17873
rect 21637 17833 21649 17867
rect 21683 17864 21695 17867
rect 26050 17864 26056 17876
rect 21683 17836 26056 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 9766 17756 9772 17808
rect 9824 17756 9830 17808
rect 12253 17799 12311 17805
rect 12253 17765 12265 17799
rect 12299 17796 12311 17799
rect 15194 17796 15200 17808
rect 12299 17768 15200 17796
rect 12299 17765 12311 17768
rect 12253 17759 12311 17765
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 16942 17756 16948 17808
rect 17000 17796 17006 17808
rect 17862 17796 17868 17808
rect 17000 17768 17868 17796
rect 17000 17756 17006 17768
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7892 17700 8401 17728
rect 7892 17688 7898 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 9784 17728 9812 17756
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9784 17700 10057 17728
rect 8389 17691 8447 17697
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17728 12955 17731
rect 13354 17728 13360 17740
rect 12943 17700 13360 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 16022 17688 16028 17740
rect 16080 17728 16086 17740
rect 16393 17731 16451 17737
rect 16393 17728 16405 17731
rect 16080 17700 16405 17728
rect 16080 17688 16086 17700
rect 16393 17697 16405 17700
rect 16439 17697 16451 17731
rect 16393 17691 16451 17697
rect 17494 17688 17500 17740
rect 17552 17728 17558 17740
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 17552 17700 17969 17728
rect 17552 17688 17558 17700
rect 17957 17697 17969 17700
rect 18003 17697 18015 17731
rect 17957 17691 18015 17697
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 19613 17731 19671 17737
rect 19613 17728 19625 17731
rect 19484 17700 19625 17728
rect 19484 17688 19490 17700
rect 19613 17697 19625 17700
rect 19659 17697 19671 17731
rect 19613 17691 19671 17697
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 19852 17700 21128 17728
rect 19852 17688 19858 17700
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9640 17632 9781 17660
rect 9640 17620 9646 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 11146 17620 11152 17672
rect 11204 17620 11210 17672
rect 11330 17620 11336 17672
rect 11388 17660 11394 17672
rect 11790 17660 11796 17672
rect 11388 17632 11796 17660
rect 11388 17620 11394 17632
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 14274 17660 14280 17672
rect 12667 17632 14280 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 16114 17620 16120 17672
rect 16172 17620 16178 17672
rect 17770 17620 17776 17672
rect 17828 17660 17834 17672
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 17828 17632 18797 17660
rect 17828 17620 17834 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 19702 17620 19708 17672
rect 19760 17660 19766 17672
rect 21100 17669 21128 17700
rect 22020 17669 22048 17836
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24854 17728 24860 17740
rect 23891 17700 24860 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19760 17632 19901 17660
rect 19760 17620 19766 17632
rect 19889 17629 19901 17632
rect 19935 17629 19947 17663
rect 19889 17623 19947 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17660 22891 17663
rect 24578 17660 24584 17672
rect 22879 17632 24584 17660
rect 22879 17629 22891 17632
rect 22833 17623 22891 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 8205 17595 8263 17601
rect 8205 17561 8217 17595
rect 8251 17592 8263 17595
rect 8754 17592 8760 17604
rect 8251 17564 8760 17592
rect 8251 17561 8263 17564
rect 8205 17555 8263 17561
rect 8754 17552 8760 17564
rect 8812 17552 8818 17604
rect 12434 17552 12440 17604
rect 12492 17592 12498 17604
rect 14185 17595 14243 17601
rect 14185 17592 14197 17595
rect 12492 17564 14197 17592
rect 12492 17552 12498 17564
rect 14185 17561 14197 17564
rect 14231 17592 14243 17595
rect 17678 17592 17684 17604
rect 14231 17564 17684 17592
rect 14231 17561 14243 17564
rect 14185 17555 14243 17561
rect 17678 17552 17684 17564
rect 17736 17552 17742 17604
rect 17862 17552 17868 17604
rect 17920 17592 17926 17604
rect 18601 17595 18659 17601
rect 18601 17592 18613 17595
rect 17920 17564 18613 17592
rect 17920 17552 17926 17564
rect 18601 17561 18613 17564
rect 18647 17592 18659 17595
rect 19242 17592 19248 17604
rect 18647 17564 19248 17592
rect 18647 17561 18659 17564
rect 18601 17555 18659 17561
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 19794 17552 19800 17604
rect 19852 17592 19858 17604
rect 20254 17592 20260 17604
rect 19852 17564 20260 17592
rect 19852 17552 19858 17564
rect 20254 17552 20260 17564
rect 20312 17552 20318 17604
rect 20916 17564 22094 17592
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 8294 17484 8300 17536
rect 8352 17484 8358 17536
rect 9125 17527 9183 17533
rect 9125 17493 9137 17527
rect 9171 17524 9183 17527
rect 9398 17524 9404 17536
rect 9171 17496 9404 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 12066 17484 12072 17536
rect 12124 17524 12130 17536
rect 12713 17527 12771 17533
rect 12713 17524 12725 17527
rect 12124 17496 12725 17524
rect 12124 17484 12130 17496
rect 12713 17493 12725 17496
rect 12759 17493 12771 17527
rect 12713 17487 12771 17493
rect 13170 17484 13176 17536
rect 13228 17524 13234 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 13228 17496 13461 17524
rect 13228 17484 13234 17496
rect 13449 17493 13461 17496
rect 13495 17493 13507 17527
rect 13449 17487 13507 17493
rect 15470 17484 15476 17536
rect 15528 17484 15534 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 15746 17524 15752 17536
rect 15620 17496 15752 17524
rect 15620 17484 15626 17496
rect 15746 17484 15752 17496
rect 15804 17524 15810 17536
rect 16298 17524 16304 17536
rect 15804 17496 16304 17524
rect 15804 17484 15810 17496
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 17402 17484 17408 17536
rect 17460 17484 17466 17536
rect 20916 17533 20944 17564
rect 20901 17527 20959 17533
rect 20901 17493 20913 17527
rect 20947 17493 20959 17527
rect 22066 17524 22094 17564
rect 22186 17552 22192 17604
rect 22244 17552 22250 17604
rect 25038 17592 25044 17604
rect 22296 17564 25044 17592
rect 22296 17524 22324 17564
rect 25038 17552 25044 17564
rect 25096 17552 25102 17604
rect 22066 17496 22324 17524
rect 20901 17487 20959 17493
rect 22830 17484 22836 17536
rect 22888 17524 22894 17536
rect 24581 17527 24639 17533
rect 24581 17524 24593 17527
rect 22888 17496 24593 17524
rect 22888 17484 22894 17496
rect 24581 17493 24593 17496
rect 24627 17493 24639 17527
rect 24581 17487 24639 17493
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24728 17496 24961 17524
rect 24728 17484 24734 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7248 17292 8033 17320
rect 7248 17280 7254 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8444 17292 9045 17320
rect 8444 17280 8450 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11388 17292 11621 17320
rect 11388 17280 11394 17292
rect 11609 17289 11621 17292
rect 11655 17320 11667 17323
rect 12434 17320 12440 17332
rect 11655 17292 12440 17320
rect 11655 17289 11667 17292
rect 11609 17283 11667 17289
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 13170 17280 13176 17332
rect 13228 17280 13234 17332
rect 16390 17320 16396 17332
rect 14568 17292 16396 17320
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 9640 17224 10977 17252
rect 9640 17212 9646 17224
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 8570 17184 8576 17196
rect 8312 17156 8576 17184
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 8312 17125 8340 17156
rect 8570 17144 8576 17156
rect 8628 17184 8634 17196
rect 8938 17184 8944 17196
rect 8628 17156 8944 17184
rect 8628 17144 8634 17156
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 11330 17184 11336 17196
rect 10275 17156 11336 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12802 17184 12808 17196
rect 12492 17156 12808 17184
rect 12492 17144 12498 17156
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 14568 17193 14596 17292
rect 16390 17280 16396 17292
rect 16448 17320 16454 17332
rect 16758 17320 16764 17332
rect 16448 17292 16764 17320
rect 16448 17280 16454 17292
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 20346 17280 20352 17332
rect 20404 17280 20410 17332
rect 22738 17280 22744 17332
rect 22796 17280 22802 17332
rect 16114 17252 16120 17264
rect 16054 17224 16120 17252
rect 16114 17212 16120 17224
rect 16172 17212 16178 17264
rect 16945 17255 17003 17261
rect 16945 17221 16957 17255
rect 16991 17252 17003 17255
rect 17126 17252 17132 17264
rect 16991 17224 17132 17252
rect 16991 17221 17003 17224
rect 16945 17215 17003 17221
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 17957 17255 18015 17261
rect 17957 17221 17969 17255
rect 18003 17252 18015 17255
rect 18414 17252 18420 17264
rect 18003 17224 18420 17252
rect 18003 17221 18015 17224
rect 17957 17215 18015 17221
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 23750 17212 23756 17264
rect 23808 17212 23814 17264
rect 24210 17212 24216 17264
rect 24268 17212 24274 17264
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 19978 17144 19984 17196
rect 20036 17144 20042 17196
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 21315 17156 22661 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 8113 17119 8171 17125
rect 7340 17088 7696 17116
rect 7340 17076 7346 17088
rect 7668 17057 7696 17088
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17085 8355 17119
rect 8297 17079 8355 17085
rect 8757 17119 8815 17125
rect 8757 17085 8769 17119
rect 8803 17116 8815 17119
rect 9398 17116 9404 17128
rect 8803 17088 9404 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 7653 17051 7711 17057
rect 7653 17017 7665 17051
rect 7699 17017 7711 17051
rect 7653 17011 7711 17017
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 7285 16983 7343 16989
rect 7285 16980 7297 16983
rect 3384 16952 7297 16980
rect 3384 16940 3390 16952
rect 7285 16949 7297 16952
rect 7331 16980 7343 16983
rect 8128 16980 8156 17079
rect 9398 17076 9404 17088
rect 9456 17116 9462 17128
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 9456 17088 9505 17116
rect 9456 17076 9462 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9582 17076 9588 17128
rect 9640 17076 9646 17128
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11885 17119 11943 17125
rect 11885 17116 11897 17119
rect 11204 17088 11897 17116
rect 11204 17076 11210 17088
rect 11885 17085 11897 17088
rect 11931 17116 11943 17119
rect 12529 17119 12587 17125
rect 11931 17088 12434 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 7331 16952 8156 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 12066 16940 12072 16992
rect 12124 16940 12130 16992
rect 12406 16980 12434 17088
rect 12529 17085 12541 17119
rect 12575 17116 12587 17119
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 12575 17088 13277 17116
rect 12575 17085 12587 17088
rect 12529 17079 12587 17085
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13280 17048 13308 17079
rect 13446 17076 13452 17128
rect 13504 17076 13510 17128
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 15562 17116 15568 17128
rect 14875 17088 15568 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 16298 17076 16304 17128
rect 16356 17076 16362 17128
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 17920 17088 18613 17116
rect 17920 17076 17926 17088
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 18874 17076 18880 17128
rect 18932 17076 18938 17128
rect 22830 17076 22836 17128
rect 22888 17116 22894 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22888 17088 22937 17116
rect 22888 17076 22894 17088
rect 22925 17085 22937 17088
rect 22971 17116 22983 17119
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 22971 17088 25237 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 25225 17085 25237 17088
rect 25271 17085 25283 17119
rect 25225 17079 25283 17085
rect 13630 17048 13636 17060
rect 13280 17020 13636 17048
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 15930 17008 15936 17060
rect 15988 17048 15994 17060
rect 17129 17051 17187 17057
rect 17129 17048 17141 17051
rect 15988 17020 17141 17048
rect 15988 17008 15994 17020
rect 17129 17017 17141 17020
rect 17175 17017 17187 17051
rect 18141 17051 18199 17057
rect 18141 17048 18153 17051
rect 17129 17011 17187 17017
rect 17236 17020 18153 17048
rect 12710 16980 12716 16992
rect 12406 16952 12716 16980
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16980 12863 16983
rect 15378 16980 15384 16992
rect 12851 16952 15384 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 16298 16940 16304 16992
rect 16356 16980 16362 16992
rect 17236 16980 17264 17020
rect 18141 17017 18153 17020
rect 18187 17017 18199 17051
rect 18141 17011 18199 17017
rect 16356 16952 17264 16980
rect 16356 16940 16362 16952
rect 17494 16940 17500 16992
rect 17552 16940 17558 16992
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 18690 16980 18696 16992
rect 18472 16952 18696 16980
rect 18472 16940 18478 16952
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 20990 16940 20996 16992
rect 21048 16980 21054 16992
rect 21818 16980 21824 16992
rect 21048 16952 21824 16980
rect 21048 16940 21054 16952
rect 21818 16940 21824 16952
rect 21876 16980 21882 16992
rect 21913 16983 21971 16989
rect 21913 16980 21925 16983
rect 21876 16952 21925 16980
rect 21876 16940 21882 16952
rect 21913 16949 21925 16952
rect 21959 16949 21971 16983
rect 21913 16943 21971 16949
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 22370 16980 22376 16992
rect 22327 16952 22376 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 8570 16736 8576 16788
rect 8628 16736 8634 16788
rect 11238 16736 11244 16788
rect 11296 16736 11302 16788
rect 13909 16779 13967 16785
rect 13909 16776 13921 16779
rect 13188 16748 13921 16776
rect 8846 16708 8852 16720
rect 2746 16680 8852 16708
rect 2406 16600 2412 16652
rect 2464 16640 2470 16652
rect 2746 16640 2774 16680
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 11606 16708 11612 16720
rect 10704 16680 11612 16708
rect 2464 16612 2774 16640
rect 2464 16600 2470 16612
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 9490 16640 9496 16652
rect 8352 16612 9496 16640
rect 8352 16600 8358 16612
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 10704 16649 10732 16680
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 11238 16640 11244 16652
rect 10919 16612 11244 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11238 16600 11244 16612
rect 11296 16640 11302 16652
rect 11698 16640 11704 16652
rect 11296 16612 11704 16640
rect 11296 16600 11302 16612
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 12526 16640 12532 16652
rect 11839 16612 12532 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 13188 16640 13216 16748
rect 13909 16745 13921 16748
rect 13955 16776 13967 16779
rect 14550 16776 14556 16788
rect 13955 16748 14556 16776
rect 13955 16745 13967 16748
rect 13909 16739 13967 16745
rect 14550 16736 14556 16748
rect 14608 16776 14614 16788
rect 15749 16779 15807 16785
rect 14608 16748 15240 16776
rect 14608 16736 14614 16748
rect 13538 16668 13544 16720
rect 13596 16708 13602 16720
rect 15212 16708 15240 16748
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 15838 16776 15844 16788
rect 15795 16748 15844 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 16114 16736 16120 16788
rect 16172 16776 16178 16788
rect 16853 16779 16911 16785
rect 16853 16776 16865 16779
rect 16172 16748 16865 16776
rect 16172 16736 16178 16748
rect 16853 16745 16865 16748
rect 16899 16776 16911 16779
rect 18414 16776 18420 16788
rect 16899 16748 18420 16776
rect 16899 16745 16911 16748
rect 16853 16739 16911 16745
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 20990 16776 20996 16788
rect 20036 16748 20996 16776
rect 20036 16736 20042 16748
rect 20990 16736 20996 16748
rect 21048 16776 21054 16788
rect 22281 16779 22339 16785
rect 22281 16776 22293 16779
rect 21048 16748 22293 16776
rect 21048 16736 21054 16748
rect 22281 16745 22293 16748
rect 22327 16776 22339 16779
rect 22922 16776 22928 16788
rect 22327 16748 22928 16776
rect 22327 16745 22339 16748
rect 22281 16739 22339 16745
rect 22922 16736 22928 16748
rect 22980 16776 22986 16788
rect 24210 16776 24216 16788
rect 22980 16748 24216 16776
rect 22980 16736 22986 16748
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 24578 16736 24584 16788
rect 24636 16736 24642 16788
rect 16132 16708 16160 16736
rect 17862 16708 17868 16720
rect 13596 16680 15148 16708
rect 15212 16680 16160 16708
rect 16684 16680 17868 16708
rect 13596 16668 13602 16680
rect 15120 16649 15148 16680
rect 12860 16612 13216 16640
rect 12860 16600 12866 16612
rect 13188 16546 13216 16612
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16609 15163 16643
rect 15105 16603 15163 16609
rect 16206 16600 16212 16652
rect 16264 16640 16270 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 16264 16612 16313 16640
rect 16264 16600 16270 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16684 16640 16712 16680
rect 17862 16668 17868 16680
rect 17920 16708 17926 16720
rect 17920 16680 18000 16708
rect 17920 16668 17926 16680
rect 17972 16649 18000 16680
rect 22554 16668 22560 16720
rect 22612 16708 22618 16720
rect 23566 16708 23572 16720
rect 22612 16680 23572 16708
rect 22612 16668 22618 16680
rect 23566 16668 23572 16680
rect 23624 16668 23630 16720
rect 16448 16612 16712 16640
rect 17957 16643 18015 16649
rect 16448 16600 16454 16612
rect 17957 16609 17969 16643
rect 18003 16609 18015 16643
rect 17957 16603 18015 16609
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 13630 16572 13636 16584
rect 13504 16544 13636 16572
rect 13504 16532 13510 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16572 14979 16575
rect 15654 16572 15660 16584
rect 14967 16544 15660 16572
rect 14967 16541 14979 16544
rect 14921 16535 14979 16541
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 16546 16544 18889 16572
rect 10410 16504 10416 16516
rect 9968 16476 10416 16504
rect 9968 16448 9996 16476
rect 10410 16464 10416 16476
rect 10468 16504 10474 16516
rect 10597 16507 10655 16513
rect 10597 16504 10609 16507
rect 10468 16476 10609 16504
rect 10468 16464 10474 16476
rect 10597 16473 10609 16476
rect 10643 16473 10655 16507
rect 10597 16467 10655 16473
rect 12069 16507 12127 16513
rect 12069 16473 12081 16507
rect 12115 16473 12127 16507
rect 14090 16504 14096 16516
rect 12069 16467 12127 16473
rect 13464 16476 14096 16504
rect 9950 16396 9956 16448
rect 10008 16396 10014 16448
rect 10226 16396 10232 16448
rect 10284 16396 10290 16448
rect 12084 16436 12112 16467
rect 13464 16436 13492 16476
rect 14090 16464 14096 16476
rect 14148 16464 14154 16516
rect 16546 16504 16574 16544
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 19076 16544 19564 16572
rect 14568 16476 16574 16504
rect 12084 16408 13492 16436
rect 13541 16439 13599 16445
rect 13541 16405 13553 16439
rect 13587 16436 13599 16439
rect 13630 16436 13636 16448
rect 13587 16408 13636 16436
rect 13587 16405 13599 16408
rect 13541 16399 13599 16405
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14274 16396 14280 16448
rect 14332 16396 14338 16448
rect 14568 16445 14596 16476
rect 17218 16464 17224 16516
rect 17276 16504 17282 16516
rect 17770 16504 17776 16516
rect 17276 16476 17776 16504
rect 17276 16464 17282 16476
rect 17770 16464 17776 16476
rect 17828 16464 17834 16516
rect 14553 16439 14611 16445
rect 14553 16405 14565 16439
rect 14599 16405 14611 16439
rect 14553 16399 14611 16405
rect 15010 16396 15016 16448
rect 15068 16396 15074 16448
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 16117 16439 16175 16445
rect 16117 16436 16129 16439
rect 15528 16408 16129 16436
rect 15528 16396 15534 16408
rect 16117 16405 16129 16408
rect 16163 16405 16175 16439
rect 16117 16399 16175 16405
rect 16206 16396 16212 16448
rect 16264 16396 16270 16448
rect 18693 16439 18751 16445
rect 18693 16405 18705 16439
rect 18739 16436 18751 16439
rect 19076 16436 19104 16544
rect 18739 16408 19104 16436
rect 19245 16439 19303 16445
rect 18739 16405 18751 16408
rect 18693 16399 18751 16405
rect 19245 16405 19257 16439
rect 19291 16436 19303 16439
rect 19426 16436 19432 16448
rect 19291 16408 19432 16436
rect 19291 16405 19303 16408
rect 19245 16399 19303 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 19536 16436 19564 16544
rect 20162 16532 20168 16584
rect 20220 16572 20226 16584
rect 20257 16575 20315 16581
rect 20257 16572 20269 16575
rect 20220 16544 20269 16572
rect 20220 16532 20226 16544
rect 20257 16541 20269 16544
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 22554 16532 22560 16584
rect 22612 16572 22618 16584
rect 22649 16575 22707 16581
rect 22649 16572 22661 16575
rect 22612 16544 22661 16572
rect 22612 16532 22618 16544
rect 22649 16541 22661 16544
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 23842 16532 23848 16584
rect 23900 16532 23906 16584
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 20533 16507 20591 16513
rect 20533 16473 20545 16507
rect 20579 16504 20591 16507
rect 20622 16504 20628 16516
rect 20579 16476 20628 16504
rect 20579 16473 20591 16476
rect 20533 16467 20591 16473
rect 20622 16464 20628 16476
rect 20680 16464 20686 16516
rect 20990 16464 20996 16516
rect 21048 16464 21054 16516
rect 24780 16504 24808 16535
rect 21836 16476 24808 16504
rect 21836 16436 21864 16476
rect 19536 16408 21864 16436
rect 21910 16396 21916 16448
rect 21968 16436 21974 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 21968 16408 22017 16436
rect 21968 16396 21974 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8478 16232 8484 16244
rect 8343 16204 8484 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 8665 16235 8723 16241
rect 8665 16201 8677 16235
rect 8711 16232 8723 16235
rect 9122 16232 9128 16244
rect 8711 16204 9128 16232
rect 8711 16201 8723 16204
rect 8665 16195 8723 16201
rect 8570 16164 8576 16176
rect 8050 16136 8576 16164
rect 8570 16124 8576 16136
rect 8628 16164 8634 16176
rect 8680 16164 8708 16195
rect 9122 16192 9128 16204
rect 9180 16232 9186 16244
rect 9306 16232 9312 16244
rect 9180 16204 9312 16232
rect 9180 16192 9186 16204
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 13357 16235 13415 16241
rect 13357 16232 13369 16235
rect 11664 16204 13369 16232
rect 11664 16192 11670 16204
rect 13357 16201 13369 16204
rect 13403 16201 13415 16235
rect 13357 16195 13415 16201
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 13596 16204 13829 16232
rect 13596 16192 13602 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 13817 16195 13875 16201
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 15010 16232 15016 16244
rect 14599 16204 15016 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 15712 16204 15761 16232
rect 15712 16192 15718 16204
rect 15749 16201 15761 16204
rect 15795 16201 15807 16235
rect 15749 16195 15807 16201
rect 16853 16235 16911 16241
rect 16853 16201 16865 16235
rect 16899 16232 16911 16235
rect 17218 16232 17224 16244
rect 16899 16204 17224 16232
rect 16899 16201 16911 16204
rect 16853 16195 16911 16201
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 21177 16235 21235 16241
rect 21177 16201 21189 16235
rect 21223 16232 21235 16235
rect 21358 16232 21364 16244
rect 21223 16204 21364 16232
rect 21223 16201 21235 16204
rect 21177 16195 21235 16201
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 23290 16232 23296 16244
rect 22664 16204 23296 16232
rect 8628 16136 8708 16164
rect 8628 16124 8634 16136
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 12529 16167 12587 16173
rect 11848 16136 12434 16164
rect 11848 16124 11854 16136
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 8386 16028 8392 16040
rect 6871 16000 8392 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 8386 15988 8392 16000
rect 8444 16028 8450 16040
rect 9582 16028 9588 16040
rect 8444 16000 9588 16028
rect 8444 15988 8450 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 12158 15920 12164 15972
rect 12216 15920 12222 15972
rect 12250 15920 12256 15972
rect 12308 15960 12314 15972
rect 12406 15960 12434 16136
rect 12529 16133 12541 16167
rect 12575 16164 12587 16167
rect 13998 16164 14004 16176
rect 12575 16136 14004 16164
rect 12575 16133 12587 16136
rect 12529 16127 12587 16133
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 14090 16124 14096 16176
rect 14148 16164 14154 16176
rect 19794 16164 19800 16176
rect 14148 16136 15148 16164
rect 14148 16124 14154 16136
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 13725 16099 13783 16105
rect 12667 16068 13676 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12713 16031 12771 16037
rect 12713 15997 12725 16031
rect 12759 15997 12771 16031
rect 13648 16028 13676 16068
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 14274 16096 14280 16108
rect 13771 16068 14280 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14792 16068 14933 16096
rect 14792 16056 14798 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 13814 16028 13820 16040
rect 13648 16000 13820 16028
rect 12713 15991 12771 15997
rect 12728 15960 12756 15991
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 14458 16028 14464 16040
rect 14047 16000 14464 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 14458 15988 14464 16000
rect 14516 15988 14522 16040
rect 15120 16037 15148 16136
rect 18708 16136 19800 16164
rect 17218 16056 17224 16108
rect 17276 16056 17282 16108
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18506 16096 18512 16108
rect 18095 16068 18512 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 18708 16105 18736 16136
rect 19794 16124 19800 16136
rect 19852 16124 19858 16176
rect 20073 16167 20131 16173
rect 20073 16133 20085 16167
rect 20119 16164 20131 16167
rect 20162 16164 20168 16176
rect 20119 16136 20168 16164
rect 20119 16133 20131 16136
rect 20073 16127 20131 16133
rect 20162 16124 20168 16136
rect 20220 16164 20226 16176
rect 22278 16164 22284 16176
rect 20220 16136 22284 16164
rect 20220 16124 20226 16136
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16096 19303 16099
rect 19426 16096 19432 16108
rect 19291 16068 19432 16096
rect 19291 16065 19303 16068
rect 19245 16059 19303 16065
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 15997 15071 16031
rect 15013 15991 15071 15997
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 15997 15163 16031
rect 15105 15991 15163 15997
rect 12308 15932 12756 15960
rect 15028 15960 15056 15991
rect 17770 15988 17776 16040
rect 17828 16028 17834 16040
rect 19260 16028 19288 16059
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20864 16068 21097 16096
rect 20864 16056 20870 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21910 16096 21916 16108
rect 21085 16059 21143 16065
rect 21284 16068 21916 16096
rect 17828 16000 19288 16028
rect 17828 15988 17834 16000
rect 20530 15988 20536 16040
rect 20588 16028 20594 16040
rect 21284 16028 21312 16068
rect 21910 16056 21916 16068
rect 21968 16056 21974 16108
rect 22020 16105 22048 16136
rect 22278 16124 22284 16136
rect 22336 16164 22342 16176
rect 22664 16164 22692 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 22336 16136 22692 16164
rect 22336 16124 22342 16136
rect 22922 16124 22928 16176
rect 22980 16124 22986 16176
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 20588 16000 21312 16028
rect 21361 16031 21419 16037
rect 20588 15988 20594 16000
rect 21361 15997 21373 16031
rect 21407 16028 21419 16031
rect 22281 16031 22339 16037
rect 22281 16028 22293 16031
rect 21407 16000 21864 16028
rect 21407 15997 21419 16000
rect 21361 15991 21419 15997
rect 15470 15960 15476 15972
rect 15028 15932 15476 15960
rect 12308 15920 12314 15932
rect 15470 15920 15476 15932
rect 15528 15960 15534 15972
rect 16666 15960 16672 15972
rect 15528 15932 16672 15960
rect 15528 15920 15534 15932
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 16206 15892 16212 15904
rect 15436 15864 16212 15892
rect 15436 15852 15442 15864
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 17184 15864 17325 15892
rect 17184 15852 17190 15864
rect 17313 15861 17325 15864
rect 17359 15861 17371 15895
rect 17313 15855 17371 15861
rect 17862 15852 17868 15904
rect 17920 15852 17926 15904
rect 18506 15852 18512 15904
rect 18564 15852 18570 15904
rect 20714 15852 20720 15904
rect 20772 15852 20778 15904
rect 21836 15892 21864 16000
rect 22066 16000 22293 16028
rect 21910 15920 21916 15972
rect 21968 15960 21974 15972
rect 22066 15960 22094 16000
rect 22281 15997 22293 16000
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 24489 16031 24547 16037
rect 24489 15997 24501 16031
rect 24535 16028 24547 16031
rect 24578 16028 24584 16040
rect 24535 16000 24584 16028
rect 24535 15997 24547 16000
rect 24489 15991 24547 15997
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 24765 16031 24823 16037
rect 24765 15997 24777 16031
rect 24811 15997 24823 16031
rect 24765 15991 24823 15997
rect 21968 15932 22094 15960
rect 21968 15920 21974 15932
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 24780 15960 24808 15991
rect 23532 15932 24808 15960
rect 23532 15920 23538 15932
rect 22646 15892 22652 15904
rect 21836 15864 22652 15892
rect 22646 15852 22652 15864
rect 22704 15892 22710 15904
rect 23753 15895 23811 15901
rect 23753 15892 23765 15895
rect 22704 15864 23765 15892
rect 22704 15852 22710 15864
rect 23753 15861 23765 15864
rect 23799 15861 23811 15895
rect 23753 15855 23811 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 9125 15691 9183 15697
rect 9125 15657 9137 15691
rect 9171 15688 9183 15691
rect 9214 15688 9220 15700
rect 9171 15660 9220 15688
rect 9171 15657 9183 15660
rect 9125 15651 9183 15657
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 9364 15660 10149 15688
rect 9364 15648 9370 15660
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 10137 15651 10195 15657
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11112 15660 11621 15688
rect 11112 15648 11118 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 15470 15648 15476 15700
rect 15528 15648 15534 15700
rect 18690 15688 18696 15700
rect 15580 15660 18696 15688
rect 5166 15580 5172 15632
rect 5224 15620 5230 15632
rect 12066 15620 12072 15632
rect 5224 15592 12072 15620
rect 5224 15580 5230 15592
rect 12066 15580 12072 15592
rect 12124 15580 12130 15632
rect 14274 15580 14280 15632
rect 14332 15620 14338 15632
rect 15580 15620 15608 15660
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 20714 15648 20720 15700
rect 20772 15688 20778 15700
rect 24394 15688 24400 15700
rect 20772 15660 24400 15688
rect 20772 15648 20778 15660
rect 24394 15648 24400 15660
rect 24452 15648 24458 15700
rect 14332 15592 15608 15620
rect 14332 15580 14338 15592
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9640 15524 9689 15552
rect 9640 15512 9646 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12308 15524 12633 15552
rect 12308 15512 12314 15524
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 16390 15512 16396 15564
rect 16448 15512 16454 15564
rect 16669 15555 16727 15561
rect 16669 15521 16681 15555
rect 16715 15552 16727 15555
rect 18598 15552 18604 15564
rect 16715 15524 18604 15552
rect 16715 15521 16727 15524
rect 16669 15515 16727 15521
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 20162 15552 20168 15564
rect 19475 15524 20168 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 20162 15512 20168 15524
rect 20220 15512 20226 15564
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15552 22615 15555
rect 22646 15552 22652 15564
rect 22603 15524 22652 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15552 24639 15555
rect 24670 15552 24676 15564
rect 24627 15524 24676 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 13173 15487 13231 15493
rect 13173 15484 13185 15487
rect 5500 15456 13185 15484
rect 5500 15444 5506 15456
rect 13173 15453 13185 15456
rect 13219 15484 13231 15487
rect 13538 15484 13544 15496
rect 13219 15456 13544 15484
rect 13219 15453 13231 15456
rect 13173 15447 13231 15453
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 21692 15456 21833 15484
rect 21692 15444 21698 15456
rect 21821 15453 21833 15456
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 9585 15419 9643 15425
rect 9585 15416 9597 15419
rect 9272 15388 9597 15416
rect 9272 15376 9278 15388
rect 9585 15385 9597 15388
rect 9631 15385 9643 15419
rect 9585 15379 9643 15385
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12526 15416 12532 15428
rect 12023 15388 12532 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 17894 15388 18460 15416
rect 18432 15360 18460 15388
rect 19610 15376 19616 15428
rect 19668 15416 19674 15428
rect 19705 15419 19763 15425
rect 19705 15416 19717 15419
rect 19668 15388 19717 15416
rect 19668 15376 19674 15388
rect 19705 15385 19717 15388
rect 19751 15385 19763 15419
rect 20990 15416 20996 15428
rect 20930 15388 20996 15416
rect 19705 15379 19763 15385
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 10042 15348 10048 15360
rect 9539 15320 10048 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 12710 15348 12716 15360
rect 12115 15320 12716 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14182 15348 14188 15360
rect 13872 15320 14188 15348
rect 13872 15308 13878 15320
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 15746 15308 15752 15360
rect 15804 15308 15810 15360
rect 17678 15308 17684 15360
rect 17736 15348 17742 15360
rect 18141 15351 18199 15357
rect 18141 15348 18153 15351
rect 17736 15320 18153 15348
rect 17736 15308 17742 15320
rect 18141 15317 18153 15320
rect 18187 15317 18199 15351
rect 18141 15311 18199 15317
rect 18414 15308 18420 15360
rect 18472 15348 18478 15360
rect 18969 15351 19027 15357
rect 18969 15348 18981 15351
rect 18472 15320 18981 15348
rect 18472 15308 18478 15320
rect 18969 15317 18981 15320
rect 19015 15317 19027 15351
rect 19720 15348 19748 15379
rect 20990 15376 20996 15388
rect 21048 15416 21054 15428
rect 21450 15416 21456 15428
rect 21048 15388 21456 15416
rect 21048 15376 21054 15388
rect 21450 15376 21456 15388
rect 21508 15416 21514 15428
rect 22646 15416 22652 15428
rect 21508 15388 22652 15416
rect 21508 15376 21514 15388
rect 22646 15376 22652 15388
rect 22704 15416 22710 15428
rect 22704 15388 23046 15416
rect 22704 15376 22710 15388
rect 20346 15348 20352 15360
rect 19720 15320 20352 15348
rect 18969 15311 19027 15317
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 20622 15308 20628 15360
rect 20680 15348 20686 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 20680 15320 21189 15348
rect 20680 15308 20686 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 21637 15351 21695 15357
rect 21637 15317 21649 15351
rect 21683 15348 21695 15351
rect 21910 15348 21916 15360
rect 21683 15320 21916 15348
rect 21683 15317 21695 15320
rect 21637 15311 21695 15317
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 23566 15308 23572 15360
rect 23624 15348 23630 15360
rect 24029 15351 24087 15357
rect 24029 15348 24041 15351
rect 23624 15320 24041 15348
rect 23624 15308 23630 15320
rect 24029 15317 24041 15320
rect 24075 15317 24087 15351
rect 24029 15311 24087 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 10134 15104 10140 15156
rect 10192 15104 10198 15156
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 11330 15144 11336 15156
rect 10284 15116 11336 15144
rect 10284 15104 10290 15116
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 12066 15104 12072 15156
rect 12124 15144 12130 15156
rect 12802 15144 12808 15156
rect 12124 15116 12808 15144
rect 12124 15104 12130 15116
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14274 15144 14280 15156
rect 14139 15116 14280 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15804 15116 15945 15144
rect 15804 15104 15810 15116
rect 15933 15113 15945 15116
rect 15979 15113 15991 15147
rect 15933 15107 15991 15113
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 17497 15147 17555 15153
rect 17497 15144 17509 15147
rect 17276 15116 17509 15144
rect 17276 15104 17282 15116
rect 17497 15113 17509 15116
rect 17543 15113 17555 15147
rect 17497 15107 17555 15113
rect 20070 15104 20076 15156
rect 20128 15104 20134 15156
rect 22830 15144 22836 15156
rect 20180 15116 22836 15144
rect 8570 15036 8576 15088
rect 8628 15036 8634 15088
rect 18693 15079 18751 15085
rect 18693 15045 18705 15079
rect 18739 15076 18751 15079
rect 18782 15076 18788 15088
rect 18739 15048 18788 15076
rect 18739 15045 18751 15048
rect 18693 15039 18751 15045
rect 18782 15036 18788 15048
rect 18840 15036 18846 15088
rect 20180 15076 20208 15116
rect 22830 15104 22836 15116
rect 22888 15104 22894 15156
rect 23198 15076 23204 15088
rect 18892 15048 20208 15076
rect 21008 15048 23204 15076
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 9640 14980 9812 15008
rect 9640 14968 9646 14980
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7929 14943 7987 14949
rect 7699 14912 7788 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7760 14804 7788 14912
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8478 14940 8484 14952
rect 7975 14912 8484 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 9784 14940 9812 14980
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 11606 15008 11612 15020
rect 10643 14980 11612 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 14458 15008 14464 15020
rect 11848 14980 14464 15008
rect 11848 14968 11854 14980
rect 14458 14968 14464 14980
rect 14516 14968 14522 15020
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 16025 15011 16083 15017
rect 16025 15008 16037 15011
rect 15252 14980 16037 15008
rect 15252 14968 15258 14980
rect 16025 14977 16037 14980
rect 16071 14977 16083 15011
rect 16025 14971 16083 14977
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 18892 15008 18920 15048
rect 18656 14980 18920 15008
rect 18656 14968 18662 14980
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 21008 15017 21036 15048
rect 23198 15036 23204 15048
rect 23256 15036 23262 15088
rect 23290 15036 23296 15088
rect 23348 15036 23354 15088
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21450 14968 21456 15020
rect 21508 15008 21514 15020
rect 21545 15011 21603 15017
rect 21545 15008 21557 15011
rect 21508 14980 21557 15008
rect 21508 14968 21514 14980
rect 21545 14977 21557 14980
rect 21591 14977 21603 15011
rect 21545 14971 21603 14977
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 22060 14980 22109 15008
rect 22060 14968 22066 14980
rect 22097 14977 22109 14980
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 9784 14912 10701 14940
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 10689 14903 10747 14909
rect 13372 14912 14197 14940
rect 11422 14832 11428 14884
rect 11480 14872 11486 14884
rect 13372 14881 13400 14912
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 15654 14940 15660 14952
rect 14415 14912 15660 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 16850 14940 16856 14952
rect 16255 14912 16856 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 20257 14943 20315 14949
rect 20257 14909 20269 14943
rect 20303 14940 20315 14943
rect 20622 14940 20628 14952
rect 20303 14912 20628 14940
rect 20303 14909 20315 14912
rect 20257 14903 20315 14909
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 24762 14900 24768 14952
rect 24820 14900 24826 14952
rect 13357 14875 13415 14881
rect 13357 14872 13369 14875
rect 11480 14844 13369 14872
rect 11480 14832 11486 14844
rect 13357 14841 13369 14844
rect 13403 14841 13415 14875
rect 13357 14835 13415 14841
rect 13725 14875 13783 14881
rect 13725 14841 13737 14875
rect 13771 14872 13783 14875
rect 14642 14872 14648 14884
rect 13771 14844 14648 14872
rect 13771 14841 13783 14844
rect 13725 14835 13783 14841
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 15565 14875 15623 14881
rect 15565 14841 15577 14875
rect 15611 14872 15623 14875
rect 18966 14872 18972 14884
rect 15611 14844 18972 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 19613 14875 19671 14881
rect 19613 14841 19625 14875
rect 19659 14872 19671 14875
rect 24670 14872 24676 14884
rect 19659 14844 24676 14872
rect 19659 14841 19671 14844
rect 19613 14835 19671 14841
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 8294 14804 8300 14816
rect 7760 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 12066 14804 12072 14816
rect 11204 14776 12072 14804
rect 11204 14764 11210 14776
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 12529 14807 12587 14813
rect 12529 14773 12541 14807
rect 12575 14804 12587 14807
rect 12802 14804 12808 14816
rect 12575 14776 12808 14804
rect 12575 14773 12587 14776
rect 12529 14767 12587 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 15194 14764 15200 14816
rect 15252 14764 15258 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 18785 14807 18843 14813
rect 18785 14804 18797 14807
rect 17000 14776 18797 14804
rect 17000 14764 17006 14776
rect 18785 14773 18797 14776
rect 18831 14773 18843 14807
rect 18785 14767 18843 14773
rect 20809 14807 20867 14813
rect 20809 14773 20821 14807
rect 20855 14804 20867 14807
rect 21450 14804 21456 14816
rect 20855 14776 21456 14804
rect 20855 14773 20867 14776
rect 20809 14767 20867 14773
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7892 14572 8217 14600
rect 7892 14560 7898 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 8570 14560 8576 14612
rect 8628 14600 8634 14612
rect 9585 14603 9643 14609
rect 9585 14600 9597 14603
rect 8628 14572 9597 14600
rect 8628 14560 8634 14572
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 8294 14464 8300 14476
rect 6512 14436 8300 14464
rect 6512 14424 6518 14436
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8570 14396 8576 14408
rect 7866 14368 8576 14396
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 6733 14331 6791 14337
rect 6733 14297 6745 14331
rect 6779 14297 6791 14331
rect 9030 14328 9036 14340
rect 6733 14291 6791 14297
rect 8404 14300 9036 14328
rect 6748 14260 6776 14291
rect 8404 14260 8432 14300
rect 9030 14288 9036 14300
rect 9088 14288 9094 14340
rect 9508 14328 9536 14572
rect 9585 14569 9597 14572
rect 9631 14569 9643 14603
rect 9585 14563 9643 14569
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10216 14603 10274 14609
rect 10216 14600 10228 14603
rect 9916 14572 10228 14600
rect 9916 14560 9922 14572
rect 10216 14569 10228 14572
rect 10262 14600 10274 14603
rect 11790 14600 11796 14612
rect 10262 14572 11796 14600
rect 10262 14569 10274 14572
rect 10216 14563 10274 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 12437 14603 12495 14609
rect 12437 14569 12449 14603
rect 12483 14600 12495 14603
rect 12618 14600 12624 14612
rect 12483 14572 12624 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 15746 14600 15752 14612
rect 14844 14572 15752 14600
rect 14844 14532 14872 14572
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 20162 14600 20168 14612
rect 16632 14572 20168 14600
rect 16632 14560 16638 14572
rect 20162 14560 20168 14572
rect 20220 14560 20226 14612
rect 11256 14504 14872 14532
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 11256 14464 11284 14504
rect 9732 14436 11284 14464
rect 9732 14424 9738 14436
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11756 14436 11989 14464
rect 11756 14424 11762 14436
rect 11977 14433 11989 14436
rect 12023 14464 12035 14467
rect 12158 14464 12164 14476
rect 12023 14436 12164 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 12158 14424 12164 14436
rect 12216 14464 12222 14476
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 12216 14436 13001 14464
rect 12216 14424 12222 14436
rect 12989 14433 13001 14436
rect 13035 14433 13047 14467
rect 14734 14464 14740 14476
rect 12989 14427 13047 14433
rect 13832 14436 14740 14464
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 13832 14405 13860 14436
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 14844 14473 14872 14504
rect 15562 14492 15568 14544
rect 15620 14532 15626 14544
rect 15620 14504 17080 14532
rect 15620 14492 15626 14504
rect 14829 14467 14887 14473
rect 14829 14433 14841 14467
rect 14875 14433 14887 14467
rect 14829 14427 14887 14433
rect 14918 14424 14924 14476
rect 14976 14464 14982 14476
rect 17052 14473 17080 14504
rect 17586 14492 17592 14544
rect 17644 14532 17650 14544
rect 19334 14532 19340 14544
rect 17644 14504 19340 14532
rect 17644 14492 17650 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 19702 14492 19708 14544
rect 19760 14532 19766 14544
rect 20438 14532 20444 14544
rect 19760 14504 20444 14532
rect 19760 14492 19766 14504
rect 20438 14492 20444 14504
rect 20496 14492 20502 14544
rect 21453 14535 21511 14541
rect 21453 14501 21465 14535
rect 21499 14532 21511 14535
rect 22462 14532 22468 14544
rect 21499 14504 22468 14532
rect 21499 14501 21511 14504
rect 21453 14495 21511 14501
rect 22462 14492 22468 14504
rect 22520 14492 22526 14544
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 14976 14436 16957 14464
rect 14976 14424 14982 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17037 14467 17095 14473
rect 17037 14433 17049 14467
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 21542 14424 21548 14476
rect 21600 14464 21606 14476
rect 21913 14467 21971 14473
rect 21913 14464 21925 14467
rect 21600 14436 21925 14464
rect 21600 14424 21606 14436
rect 21913 14433 21925 14436
rect 21959 14433 21971 14467
rect 21913 14427 21971 14433
rect 22094 14424 22100 14476
rect 22152 14424 22158 14476
rect 23845 14467 23903 14473
rect 23845 14433 23857 14467
rect 23891 14464 23903 14467
rect 24854 14464 24860 14476
rect 23891 14436 24860 14464
rect 23891 14433 23903 14436
rect 23845 14427 23903 14433
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9640 14368 9965 14396
rect 9640 14356 9646 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 9953 14359 10011 14365
rect 12406 14368 13829 14396
rect 9508 14300 10718 14328
rect 6748 14232 8432 14260
rect 10612 14260 10640 14300
rect 11146 14260 11152 14272
rect 10612 14232 11152 14260
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 12406 14260 12434 14368
rect 13817 14365 13829 14368
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14396 14703 14399
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 14691 14368 15393 14396
rect 14691 14365 14703 14368
rect 14645 14359 14703 14365
rect 15381 14365 15393 14368
rect 15427 14396 15439 14399
rect 16574 14396 16580 14408
rect 15427 14368 16580 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16666 14356 16672 14408
rect 16724 14396 16730 14408
rect 20254 14396 20260 14408
rect 16724 14368 20260 14396
rect 16724 14356 16730 14368
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 21818 14396 21824 14408
rect 20487 14368 21824 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 21818 14356 21824 14368
rect 21876 14356 21882 14408
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14396 22891 14399
rect 23934 14396 23940 14408
rect 22879 14368 23940 14396
rect 22879 14365 22891 14368
rect 22833 14359 22891 14365
rect 23934 14356 23940 14368
rect 23992 14356 23998 14408
rect 25038 14356 25044 14408
rect 25096 14356 25102 14408
rect 12897 14331 12955 14337
rect 12897 14297 12909 14331
rect 12943 14328 12955 14331
rect 13906 14328 13912 14340
rect 12943 14300 13912 14328
rect 12943 14297 12955 14300
rect 12897 14291 12955 14297
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 16853 14331 16911 14337
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 17681 14331 17739 14337
rect 17681 14328 17693 14331
rect 16899 14300 17693 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 17681 14297 17693 14300
rect 17727 14297 17739 14331
rect 17681 14291 17739 14297
rect 11296 14232 12434 14260
rect 11296 14220 11302 14232
rect 12802 14220 12808 14272
rect 12860 14220 12866 14272
rect 13538 14220 13544 14272
rect 13596 14220 13602 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 14366 14260 14372 14272
rect 14323 14232 14372 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 16485 14263 16543 14269
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 19610 14260 19616 14272
rect 16531 14232 19616 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 19610 14220 19616 14232
rect 19668 14220 19674 14272
rect 19794 14220 19800 14272
rect 19852 14260 19858 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 19852 14232 20269 14260
rect 19852 14220 19858 14232
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 21818 14220 21824 14272
rect 21876 14220 21882 14272
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 8294 14056 8300 14068
rect 7760 14028 8300 14056
rect 7760 13929 7788 14028
rect 8294 14016 8300 14028
rect 8352 14056 8358 14068
rect 9582 14056 9588 14068
rect 8352 14028 9588 14056
rect 8352 14016 8358 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 9824 14028 12633 14056
rect 9824 14016 9830 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 12989 14059 13047 14065
rect 12989 14025 13001 14059
rect 13035 14056 13047 14059
rect 13538 14056 13544 14068
rect 13035 14028 13544 14056
rect 13035 14025 13047 14028
rect 12989 14019 13047 14025
rect 13538 14016 13544 14028
rect 13596 14056 13602 14068
rect 16666 14056 16672 14068
rect 13596 14028 16672 14056
rect 13596 14016 13602 14028
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17310 14056 17316 14068
rect 16816 14028 17316 14056
rect 16816 14016 16822 14028
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 19613 14059 19671 14065
rect 19613 14056 19625 14059
rect 17512 14028 19625 14056
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 8021 13991 8079 13997
rect 8021 13988 8033 13991
rect 7984 13960 8033 13988
rect 7984 13948 7990 13960
rect 8021 13957 8033 13960
rect 8067 13957 8079 13991
rect 8021 13951 8079 13957
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 12434 13988 12440 14000
rect 10284 13960 12440 13988
rect 10284 13948 10290 13960
rect 12434 13948 12440 13960
rect 12492 13988 12498 14000
rect 13814 13988 13820 14000
rect 12492 13960 13820 13988
rect 12492 13948 12498 13960
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 15318 13960 15945 13988
rect 15933 13957 15945 13960
rect 15979 13988 15991 13991
rect 16114 13988 16120 14000
rect 15979 13960 16120 13988
rect 15979 13957 15991 13960
rect 15933 13951 15991 13957
rect 16114 13948 16120 13960
rect 16172 13948 16178 14000
rect 17512 13988 17540 14028
rect 19613 14025 19625 14028
rect 19659 14025 19671 14059
rect 19613 14019 19671 14025
rect 20165 14059 20223 14065
rect 20165 14025 20177 14059
rect 20211 14056 20223 14059
rect 23382 14056 23388 14068
rect 20211 14028 23388 14056
rect 20211 14025 20223 14028
rect 20165 14019 20223 14025
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 18414 13988 18420 14000
rect 16546 13960 17540 13988
rect 18354 13960 18420 13988
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 9640 13892 10977 13920
rect 9640 13880 9646 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16546 13920 16574 13960
rect 18414 13948 18420 13960
rect 18472 13988 18478 14000
rect 19061 13991 19119 13997
rect 19061 13988 19073 13991
rect 18472 13960 19073 13988
rect 18472 13948 18478 13960
rect 19061 13957 19073 13960
rect 19107 13957 19119 13991
rect 19061 13951 19119 13957
rect 19518 13948 19524 14000
rect 19576 13948 19582 14000
rect 19702 13948 19708 14000
rect 19760 13988 19766 14000
rect 22557 13991 22615 13997
rect 19760 13960 22140 13988
rect 19760 13948 19766 13960
rect 15712 13892 16574 13920
rect 15712 13880 15718 13892
rect 19610 13880 19616 13932
rect 19668 13920 19674 13932
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 19668 13892 20361 13920
rect 19668 13880 19674 13892
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13920 21143 13923
rect 21358 13920 21364 13932
rect 21131 13892 21364 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 22112 13924 22140 13960
rect 22557 13957 22569 13991
rect 22603 13988 22615 13991
rect 22646 13988 22652 14000
rect 22603 13960 22652 13988
rect 22603 13957 22615 13960
rect 22557 13951 22615 13957
rect 22646 13948 22652 13960
rect 22704 13988 22710 14000
rect 22830 13988 22836 14000
rect 22704 13960 22836 13988
rect 22704 13948 22710 13960
rect 22830 13948 22836 13960
rect 22888 13988 22894 14000
rect 22888 13960 23598 13988
rect 22888 13948 22894 13960
rect 22189 13924 22247 13929
rect 22112 13923 22247 13924
rect 22112 13896 22201 13923
rect 22189 13889 22201 13896
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 9858 13852 9864 13864
rect 9815 13824 9864 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11112 13824 11713 13852
rect 11112 13812 11118 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12308 13824 13093 13852
rect 12308 13812 12314 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 12894 13744 12900 13796
rect 12952 13784 12958 13796
rect 13280 13784 13308 13815
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13504 13824 13829 13852
rect 13504 13812 13510 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 13924 13824 15148 13852
rect 13924 13784 13952 13824
rect 12952 13756 13952 13784
rect 15120 13784 15148 13824
rect 15562 13812 15568 13864
rect 15620 13812 15626 13864
rect 16850 13812 16856 13864
rect 16908 13812 16914 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17494 13852 17500 13864
rect 17175 13824 17500 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17494 13812 17500 13824
rect 17552 13852 17558 13864
rect 18601 13855 18659 13861
rect 17552 13824 18184 13852
rect 17552 13812 17558 13824
rect 15838 13784 15844 13796
rect 15120 13756 15844 13784
rect 12952 13744 12958 13756
rect 15838 13744 15844 13756
rect 15896 13744 15902 13796
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 12158 13716 12164 13728
rect 11940 13688 12164 13716
rect 11940 13676 11946 13688
rect 12158 13676 12164 13688
rect 12216 13716 12222 13728
rect 14090 13725 14096 13728
rect 12253 13719 12311 13725
rect 12253 13716 12265 13719
rect 12216 13688 12265 13716
rect 12216 13676 12222 13688
rect 12253 13685 12265 13688
rect 12299 13685 12311 13719
rect 12253 13679 12311 13685
rect 14080 13719 14096 13725
rect 14080 13685 14092 13719
rect 14080 13679 14096 13685
rect 14090 13676 14096 13679
rect 14148 13676 14154 13728
rect 18156 13716 18184 13824
rect 18601 13821 18613 13855
rect 18647 13852 18659 13855
rect 18874 13852 18880 13864
rect 18647 13824 18880 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 21634 13852 21640 13864
rect 20916 13824 21640 13852
rect 20916 13793 20944 13824
rect 21634 13812 21640 13824
rect 21692 13812 21698 13864
rect 22554 13852 22560 13864
rect 22020 13824 22560 13852
rect 22020 13793 22048 13824
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 22646 13812 22652 13864
rect 22704 13852 22710 13864
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22704 13824 22845 13852
rect 22704 13812 22710 13824
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 23109 13855 23167 13861
rect 23109 13852 23121 13855
rect 22833 13815 22891 13821
rect 22940 13824 23121 13852
rect 20901 13787 20959 13793
rect 20901 13753 20913 13787
rect 20947 13753 20959 13787
rect 20901 13747 20959 13753
rect 22005 13787 22063 13793
rect 22005 13753 22017 13787
rect 22051 13753 22063 13787
rect 22005 13747 22063 13753
rect 22278 13744 22284 13796
rect 22336 13784 22342 13796
rect 22940 13784 22968 13824
rect 23109 13821 23121 13824
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 23198 13812 23204 13864
rect 23256 13852 23262 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 23256 13824 24593 13852
rect 23256 13812 23262 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 22336 13756 22968 13784
rect 22336 13744 22342 13756
rect 18966 13716 18972 13728
rect 18156 13688 18972 13716
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 22940 13716 22968 13756
rect 23566 13716 23572 13728
rect 22940 13688 23572 13716
rect 23566 13676 23572 13688
rect 23624 13676 23630 13728
rect 25038 13676 25044 13728
rect 25096 13676 25102 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8386 13512 8392 13524
rect 8343 13484 8392 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8570 13472 8576 13524
rect 8628 13472 8634 13524
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9217 13515 9275 13521
rect 9217 13512 9229 13515
rect 8812 13484 9229 13512
rect 8812 13472 8818 13484
rect 9217 13481 9229 13484
rect 9263 13481 9275 13515
rect 9217 13475 9275 13481
rect 10676 13515 10734 13521
rect 10676 13481 10688 13515
rect 10722 13512 10734 13515
rect 13630 13512 13636 13524
rect 10722 13484 13636 13512
rect 10722 13481 10734 13484
rect 10676 13475 10734 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 13814 13472 13820 13524
rect 13872 13472 13878 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17368 13484 17417 13512
rect 17368 13472 17374 13484
rect 17405 13481 17417 13484
rect 17451 13512 17463 13515
rect 17954 13512 17960 13524
rect 17451 13484 17960 13512
rect 17451 13481 17463 13484
rect 17405 13475 17463 13481
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 18414 13472 18420 13524
rect 18472 13512 18478 13524
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 18472 13484 21005 13512
rect 18472 13472 18478 13484
rect 20993 13481 21005 13484
rect 21039 13512 21051 13515
rect 21082 13512 21088 13524
rect 21039 13484 21088 13512
rect 21039 13481 21051 13484
rect 20993 13475 21051 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 23934 13472 23940 13524
rect 23992 13512 23998 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 23992 13484 24593 13512
rect 23992 13472 23998 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 9030 13404 9036 13456
rect 9088 13444 9094 13456
rect 9306 13444 9312 13456
rect 9088 13416 9312 13444
rect 9088 13404 9094 13416
rect 9306 13404 9312 13416
rect 9364 13444 9370 13456
rect 9364 13416 9628 13444
rect 9364 13404 9370 13416
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 6512 13348 6561 13376
rect 6512 13336 6518 13348
rect 6549 13345 6561 13348
rect 6595 13345 6607 13379
rect 9600 13376 9628 13416
rect 12894 13404 12900 13456
rect 12952 13444 12958 13456
rect 15286 13444 15292 13456
rect 12952 13416 15292 13444
rect 12952 13404 12958 13416
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 21450 13444 21456 13456
rect 17328 13416 21456 13444
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9600 13348 9781 13376
rect 6549 13339 6607 13345
rect 9769 13345 9781 13348
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 11698 13376 11704 13388
rect 10459 13348 11704 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 11698 13336 11704 13348
rect 11756 13376 11762 13388
rect 13446 13376 13452 13388
rect 11756 13348 13452 13376
rect 11756 13336 11762 13348
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 13538 13336 13544 13388
rect 13596 13376 13602 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 13596 13348 14657 13376
rect 13596 13336 13602 13348
rect 14645 13345 14657 13348
rect 14691 13376 14703 13379
rect 15194 13376 15200 13388
rect 14691 13348 15200 13376
rect 14691 13345 14703 13348
rect 14645 13339 14703 13345
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15470 13336 15476 13388
rect 15528 13376 15534 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15528 13348 15669 13376
rect 15528 13336 15534 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15746 13336 15752 13388
rect 15804 13336 15810 13388
rect 16114 13336 16120 13388
rect 16172 13376 16178 13388
rect 17328 13376 17356 13416
rect 21450 13404 21456 13416
rect 21508 13404 21514 13456
rect 18785 13379 18843 13385
rect 18785 13376 18797 13379
rect 16172 13348 17356 13376
rect 17604 13348 18797 13376
rect 16172 13336 16178 13348
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 12492 13280 12633 13308
rect 12492 13268 12498 13280
rect 12621 13277 12633 13280
rect 12667 13277 12679 13311
rect 17310 13308 17316 13320
rect 12621 13271 12679 13277
rect 16224 13280 17316 13308
rect 6825 13243 6883 13249
rect 6825 13209 6837 13243
rect 6871 13209 6883 13243
rect 8570 13240 8576 13252
rect 8050 13212 8576 13240
rect 6825 13203 6883 13209
rect 6840 13172 6868 13203
rect 8570 13200 8576 13212
rect 8628 13240 8634 13252
rect 9122 13240 9128 13252
rect 8628 13212 9128 13240
rect 8628 13200 8634 13212
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 9631 13212 11100 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 9030 13172 9036 13184
rect 6840 13144 9036 13172
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 11072 13172 11100 13212
rect 11146 13200 11152 13252
rect 11204 13200 11210 13252
rect 16224 13249 16252 13280
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17604 13308 17632 13348
rect 18785 13345 18797 13348
rect 18831 13345 18843 13379
rect 18785 13339 18843 13345
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 21637 13379 21695 13385
rect 21637 13376 21649 13379
rect 20772 13348 21649 13376
rect 20772 13336 20778 13348
rect 21637 13345 21649 13348
rect 21683 13345 21695 13379
rect 25038 13376 25044 13388
rect 21637 13339 21695 13345
rect 22848 13348 25044 13376
rect 17552 13280 17632 13308
rect 17865 13311 17923 13317
rect 17552 13268 17558 13280
rect 17865 13277 17877 13311
rect 17911 13308 17923 13311
rect 17954 13308 17960 13320
rect 17911 13280 17960 13308
rect 17911 13277 17923 13280
rect 17865 13271 17923 13277
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 19484 13280 20821 13308
rect 19484 13268 19490 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21358 13268 21364 13320
rect 21416 13268 21422 13320
rect 22848 13317 22876 13348
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 22833 13311 22891 13317
rect 22833 13277 22845 13311
rect 22879 13277 22891 13311
rect 22833 13271 22891 13277
rect 23842 13268 23848 13320
rect 23900 13268 23906 13320
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 15565 13243 15623 13249
rect 15565 13209 15577 13243
rect 15611 13240 15623 13243
rect 16209 13243 16267 13249
rect 16209 13240 16221 13243
rect 15611 13212 16221 13240
rect 15611 13209 15623 13212
rect 15565 13203 15623 13209
rect 16209 13209 16221 13212
rect 16255 13209 16267 13243
rect 16209 13203 16267 13209
rect 18601 13243 18659 13249
rect 18601 13209 18613 13243
rect 18647 13209 18659 13243
rect 18601 13203 18659 13209
rect 12066 13172 12072 13184
rect 11072 13144 12072 13172
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 12158 13132 12164 13184
rect 12216 13132 12222 13184
rect 14734 13132 14740 13184
rect 14792 13172 14798 13184
rect 14829 13175 14887 13181
rect 14829 13172 14841 13175
rect 14792 13144 14841 13172
rect 14792 13132 14798 13144
rect 14829 13141 14841 13144
rect 14875 13141 14887 13175
rect 14829 13135 14887 13141
rect 15197 13175 15255 13181
rect 15197 13141 15209 13175
rect 15243 13172 15255 13175
rect 15378 13172 15384 13184
rect 15243 13144 15384 13172
rect 15243 13141 15255 13144
rect 15197 13135 15255 13141
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17957 13175 18015 13181
rect 17957 13172 17969 13175
rect 17184 13144 17969 13172
rect 17184 13132 17190 13144
rect 17957 13141 17969 13144
rect 18003 13141 18015 13175
rect 18616 13172 18644 13203
rect 20254 13200 20260 13252
rect 20312 13200 20318 13252
rect 20717 13243 20775 13249
rect 20717 13209 20729 13243
rect 20763 13240 20775 13243
rect 21266 13240 21272 13252
rect 20763 13212 21272 13240
rect 20763 13209 20775 13212
rect 20717 13203 20775 13209
rect 18690 13172 18696 13184
rect 18616 13144 18696 13172
rect 17957 13135 18015 13141
rect 18690 13132 18696 13144
rect 18748 13172 18754 13184
rect 20732 13172 20760 13203
rect 21266 13200 21272 13212
rect 21324 13200 21330 13252
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 24780 13240 24808 13271
rect 23440 13212 24808 13240
rect 23440 13200 23446 13212
rect 18748 13144 20760 13172
rect 18748 13132 18754 13144
rect 20990 13132 20996 13184
rect 21048 13172 21054 13184
rect 22370 13172 22376 13184
rect 21048 13144 22376 13172
rect 21048 13132 21054 13144
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 7742 12968 7748 12980
rect 6687 12940 7748 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9214 12968 9220 12980
rect 9079 12940 9220 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 9493 12971 9551 12977
rect 9493 12937 9505 12971
rect 9539 12968 9551 12971
rect 9766 12968 9772 12980
rect 9539 12940 9772 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10100 12940 10425 12968
rect 10100 12928 10106 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 11054 12968 11060 12980
rect 10827 12940 11060 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 12584 12940 12633 12968
rect 12584 12928 12590 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 12621 12931 12679 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13446 12968 13452 12980
rect 13127 12940 13452 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 14918 12968 14924 12980
rect 13863 12940 14924 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 14918 12928 14924 12940
rect 14976 12928 14982 12980
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 16114 12968 16120 12980
rect 15427 12940 16120 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 16853 12971 16911 12977
rect 16853 12937 16865 12971
rect 16899 12937 16911 12971
rect 16853 12931 16911 12937
rect 17313 12971 17371 12977
rect 17313 12937 17325 12971
rect 17359 12968 17371 12971
rect 17402 12968 17408 12980
rect 17359 12940 17408 12968
rect 17359 12937 17371 12940
rect 17313 12931 17371 12937
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 6972 12872 7236 12900
rect 6972 12860 6978 12872
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7098 12724 7104 12776
rect 7156 12724 7162 12776
rect 7208 12773 7236 12872
rect 7650 12860 7656 12912
rect 7708 12900 7714 12912
rect 12342 12900 12348 12912
rect 7708 12872 12348 12900
rect 7708 12860 7714 12872
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 12989 12903 13047 12909
rect 12989 12869 13001 12903
rect 13035 12900 13047 12903
rect 15562 12900 15568 12912
rect 13035 12872 15568 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 16868 12900 16896 12931
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 17770 12928 17776 12980
rect 17828 12968 17834 12980
rect 19981 12971 20039 12977
rect 19981 12968 19993 12971
rect 17828 12940 19993 12968
rect 17828 12928 17834 12940
rect 19981 12937 19993 12940
rect 20027 12937 20039 12971
rect 19981 12931 20039 12937
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 21174 12928 21180 12980
rect 21232 12928 21238 12980
rect 21266 12928 21272 12980
rect 21324 12968 21330 12980
rect 21450 12968 21456 12980
rect 21324 12940 21456 12968
rect 21324 12928 21330 12940
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 22002 12928 22008 12980
rect 22060 12928 22066 12980
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 22888 12940 23520 12968
rect 22888 12928 22894 12940
rect 16868 12872 18460 12900
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 10919 12804 11529 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7892 12736 8309 12764
rect 7892 12724 7898 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 8662 12764 8668 12776
rect 8527 12736 8668 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 9585 12767 9643 12773
rect 9585 12764 9597 12767
rect 9088 12736 9597 12764
rect 9088 12724 9094 12736
rect 9585 12733 9597 12736
rect 9631 12764 9643 12767
rect 11054 12764 11060 12776
rect 9631 12736 11060 12764
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 11532 12764 11560 12795
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 11940 12804 13216 12832
rect 11940 12792 11946 12804
rect 12526 12764 12532 12776
rect 11532 12736 12532 12764
rect 12526 12724 12532 12736
rect 12584 12764 12590 12776
rect 12894 12764 12900 12776
rect 12584 12736 12900 12764
rect 12584 12724 12590 12736
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13188 12773 13216 12804
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13688 12804 14197 12832
rect 13688 12792 13694 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 14550 12832 14556 12844
rect 14323 12804 14556 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 18322 12832 18328 12844
rect 18279 12804 18328 12832
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 18432 12832 18460 12872
rect 18506 12860 18512 12912
rect 18564 12900 18570 12912
rect 19245 12903 19303 12909
rect 19245 12900 19257 12903
rect 18564 12872 19257 12900
rect 18564 12860 18570 12872
rect 19245 12869 19257 12872
rect 19291 12869 19303 12903
rect 20898 12900 20904 12912
rect 19245 12863 19303 12869
rect 19352 12872 20904 12900
rect 18432 12804 19104 12832
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14148 12736 14381 12764
rect 14148 12724 14154 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 15252 12736 15485 12764
rect 15252 12724 15258 12736
rect 15473 12733 15485 12736
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 15657 12767 15715 12773
rect 15657 12733 15669 12767
rect 15703 12764 15715 12767
rect 15838 12764 15844 12776
rect 15703 12736 15844 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 17497 12767 17555 12773
rect 17497 12733 17509 12767
rect 17543 12764 17555 12767
rect 18874 12764 18880 12776
rect 17543 12736 18880 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 19076 12764 19104 12804
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 19352 12764 19380 12872
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12832 20223 12835
rect 20990 12832 20996 12844
rect 20211 12804 20996 12832
rect 20211 12801 20223 12804
rect 20165 12795 20223 12801
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 21192 12832 21220 12928
rect 22094 12860 22100 12912
rect 22152 12900 22158 12912
rect 23290 12900 23296 12912
rect 22152 12872 23296 12900
rect 22152 12860 22158 12872
rect 23290 12860 23296 12872
rect 23348 12900 23354 12912
rect 23385 12903 23443 12909
rect 23385 12900 23397 12903
rect 23348 12872 23397 12900
rect 23348 12860 23354 12872
rect 23385 12869 23397 12872
rect 23431 12869 23443 12903
rect 23492 12900 23520 12940
rect 23492 12872 23874 12900
rect 23385 12863 23443 12869
rect 21192 12804 21680 12832
rect 19076 12736 19380 12764
rect 19429 12767 19487 12773
rect 19429 12733 19441 12767
rect 19475 12764 19487 12767
rect 20530 12764 20536 12776
rect 19475 12736 20536 12764
rect 19475 12733 19487 12736
rect 19429 12727 19487 12733
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12733 21419 12767
rect 21652 12764 21680 12804
rect 22002 12792 22008 12844
rect 22060 12832 22066 12844
rect 22189 12835 22247 12841
rect 22189 12832 22201 12835
rect 22060 12804 22201 12832
rect 22060 12792 22066 12804
rect 22189 12801 22201 12804
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 22465 12767 22523 12773
rect 22465 12764 22477 12767
rect 21652 12736 22477 12764
rect 21361 12727 21419 12733
rect 22465 12733 22477 12736
rect 22511 12733 22523 12767
rect 22465 12727 22523 12733
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 11204 12668 11468 12696
rect 11204 12656 11210 12668
rect 7837 12631 7895 12637
rect 7837 12597 7849 12631
rect 7883 12628 7895 12631
rect 11330 12628 11336 12640
rect 7883 12600 11336 12628
rect 7883 12597 7895 12600
rect 7837 12591 7895 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 11440 12628 11468 12668
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 15013 12699 15071 12705
rect 15013 12696 15025 12699
rect 11848 12668 15025 12696
rect 11848 12656 11854 12668
rect 15013 12665 15025 12668
rect 15059 12665 15071 12699
rect 15013 12659 15071 12665
rect 18049 12699 18107 12705
rect 18049 12665 18061 12699
rect 18095 12696 18107 12699
rect 19702 12696 19708 12708
rect 18095 12668 19708 12696
rect 18095 12665 18107 12668
rect 18049 12659 18107 12665
rect 19702 12656 19708 12668
rect 19760 12656 19766 12708
rect 20806 12696 20812 12708
rect 19904 12668 20812 12696
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 11440 12600 12081 12628
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 12069 12591 12127 12597
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 14734 12628 14740 12640
rect 12400 12600 14740 12628
rect 12400 12588 12406 12600
rect 14734 12588 14740 12600
rect 14792 12628 14798 12640
rect 15470 12628 15476 12640
rect 14792 12600 15476 12628
rect 14792 12588 14798 12600
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 18690 12628 18696 12640
rect 17368 12600 18696 12628
rect 17368 12588 17374 12600
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 18785 12631 18843 12637
rect 18785 12597 18797 12631
rect 18831 12628 18843 12631
rect 19904 12628 19932 12668
rect 20806 12656 20812 12668
rect 20864 12656 20870 12708
rect 21376 12696 21404 12727
rect 22646 12724 22652 12776
rect 22704 12764 22710 12776
rect 23109 12767 23167 12773
rect 23109 12764 23121 12767
rect 22704 12736 23121 12764
rect 22704 12724 22710 12736
rect 23109 12733 23121 12736
rect 23155 12733 23167 12767
rect 23109 12727 23167 12733
rect 22554 12696 22560 12708
rect 21376 12668 22560 12696
rect 22554 12656 22560 12668
rect 22612 12696 22618 12708
rect 22612 12668 23152 12696
rect 22612 12656 22618 12668
rect 18831 12600 19932 12628
rect 20717 12631 20775 12637
rect 18831 12597 18843 12600
rect 18785 12591 18843 12597
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 22370 12628 22376 12640
rect 20763 12600 22376 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 22370 12588 22376 12600
rect 22428 12588 22434 12640
rect 23124 12628 23152 12668
rect 24857 12631 24915 12637
rect 24857 12628 24869 12631
rect 23124 12600 24869 12628
rect 24857 12597 24869 12600
rect 24903 12597 24915 12631
rect 24857 12591 24915 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 9548 12396 10241 12424
rect 9548 12384 9554 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 11425 12427 11483 12433
rect 11425 12424 11437 12427
rect 10560 12396 11437 12424
rect 10560 12384 10566 12396
rect 11425 12393 11437 12396
rect 11471 12393 11483 12427
rect 11425 12387 11483 12393
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 12158 12424 12164 12436
rect 11940 12396 12164 12424
rect 11940 12384 11946 12396
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12618 12384 12624 12436
rect 12676 12384 12682 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 13872 12396 16313 12424
rect 13872 12384 13878 12396
rect 16301 12393 16313 12396
rect 16347 12424 16359 12427
rect 17310 12424 17316 12436
rect 16347 12396 17316 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18782 12384 18788 12436
rect 18840 12424 18846 12436
rect 20070 12424 20076 12436
rect 18840 12396 20076 12424
rect 18840 12384 18846 12396
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 21726 12424 21732 12436
rect 20220 12396 21732 12424
rect 20220 12384 20226 12396
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 24176 12396 24593 12424
rect 24176 12384 24182 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 11054 12316 11060 12368
rect 11112 12356 11118 12368
rect 11112 12328 12204 12356
rect 11112 12316 11118 12328
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7064 12260 7389 12288
rect 7064 12248 7070 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 9306 12288 9312 12300
rect 9088 12260 9312 12288
rect 9088 12248 9094 12260
rect 9306 12248 9312 12260
rect 9364 12288 9370 12300
rect 11992 12297 12020 12328
rect 12176 12300 12204 12328
rect 13998 12316 14004 12368
rect 14056 12356 14062 12368
rect 14277 12359 14335 12365
rect 14277 12356 14289 12359
rect 14056 12328 14289 12356
rect 14056 12316 14062 12328
rect 14277 12325 14289 12328
rect 14323 12325 14335 12359
rect 14277 12319 14335 12325
rect 14550 12316 14556 12368
rect 14608 12356 14614 12368
rect 15381 12359 15439 12365
rect 15381 12356 15393 12359
rect 14608 12328 15393 12356
rect 14608 12316 14614 12328
rect 15381 12325 15393 12328
rect 15427 12356 15439 12359
rect 19242 12356 19248 12368
rect 15427 12328 19248 12356
rect 15427 12325 15439 12328
rect 15381 12319 15439 12325
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 22830 12316 22836 12368
rect 22888 12316 22894 12368
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 9364 12260 10793 12288
rect 9364 12248 9370 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 11977 12291 12035 12297
rect 10781 12251 10839 12257
rect 11716 12260 11928 12288
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 11716 12220 11744 12260
rect 7524 12192 11744 12220
rect 7524 12180 7530 12192
rect 11790 12180 11796 12232
rect 11848 12180 11854 12232
rect 11900 12220 11928 12260
rect 11977 12257 11989 12291
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12158 12248 12164 12300
rect 12216 12248 12222 12300
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13722 12288 13728 12300
rect 13311 12260 13728 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14660 12260 14841 12288
rect 13740 12220 13768 12248
rect 14660 12220 14688 12260
rect 14829 12257 14841 12260
rect 14875 12288 14887 12291
rect 14918 12288 14924 12300
rect 14875 12260 14924 12288
rect 14875 12257 14887 12260
rect 14829 12251 14887 12257
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12288 15623 12291
rect 15838 12288 15844 12300
rect 15611 12260 15844 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 19150 12288 19156 12300
rect 18739 12260 19156 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19260 12260 19993 12288
rect 11900 12192 12020 12220
rect 13740 12192 14688 12220
rect 11514 12112 11520 12164
rect 11572 12152 11578 12164
rect 11885 12155 11943 12161
rect 11885 12152 11897 12155
rect 11572 12124 11897 12152
rect 11572 12112 11578 12124
rect 11885 12121 11897 12124
rect 11931 12121 11943 12155
rect 11992 12152 12020 12192
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 19260 12220 19288 12260
rect 19981 12257 19993 12260
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20254 12248 20260 12300
rect 20312 12288 20318 12300
rect 20441 12291 20499 12297
rect 20441 12288 20453 12291
rect 20312 12260 20453 12288
rect 20312 12248 20318 12260
rect 20441 12257 20453 12260
rect 20487 12257 20499 12291
rect 22002 12288 22008 12300
rect 20441 12251 20499 12257
rect 21928 12260 22008 12288
rect 18840 12192 19288 12220
rect 19521 12223 19579 12229
rect 18840 12180 18846 12192
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 20162 12220 20168 12232
rect 19567 12192 20168 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 21928 12220 21956 12260
rect 22002 12248 22008 12260
rect 22060 12288 22066 12300
rect 22848 12288 22876 12316
rect 23290 12288 23296 12300
rect 22060 12260 23296 12288
rect 22060 12248 22066 12260
rect 23290 12248 23296 12260
rect 23348 12248 23354 12300
rect 21850 12192 21956 12220
rect 22830 12180 22836 12232
rect 22888 12180 22894 12232
rect 24762 12180 24768 12232
rect 24820 12180 24826 12232
rect 13081 12155 13139 12161
rect 13081 12152 13093 12155
rect 11992 12124 13093 12152
rect 11885 12115 11943 12121
rect 13081 12121 13093 12124
rect 13127 12152 13139 12155
rect 13630 12152 13636 12164
rect 13127 12124 13636 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 13630 12112 13636 12124
rect 13688 12112 13694 12164
rect 13725 12155 13783 12161
rect 13725 12121 13737 12155
rect 13771 12152 13783 12155
rect 16482 12152 16488 12164
rect 13771 12124 16488 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8536 12056 8953 12084
rect 8536 12044 8542 12056
rect 8941 12053 8953 12056
rect 8987 12084 8999 12087
rect 9398 12084 9404 12096
rect 8987 12056 9404 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 10686 12044 10692 12096
rect 10744 12044 10750 12096
rect 11422 12044 11428 12096
rect 11480 12084 11486 12096
rect 12342 12084 12348 12096
rect 11480 12056 12348 12084
rect 11480 12044 11486 12056
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 13740 12084 13768 12115
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 18141 12155 18199 12161
rect 18141 12152 18153 12155
rect 16908 12124 18153 12152
rect 16908 12112 16914 12124
rect 18141 12121 18153 12124
rect 18187 12152 18199 12155
rect 18187 12124 18552 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 13035 12056 13768 12084
rect 13909 12087 13967 12093
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 13998 12084 14004 12096
rect 13955 12056 14004 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 13998 12044 14004 12056
rect 14056 12084 14062 12096
rect 14550 12084 14556 12096
rect 14056 12056 14556 12084
rect 14056 12044 14062 12056
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 15286 12084 15292 12096
rect 14691 12056 15292 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15286 12044 15292 12056
rect 15344 12084 15350 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 15344 12056 15761 12084
rect 15344 12044 15350 12056
rect 15749 12053 15761 12056
rect 15795 12084 15807 12087
rect 16298 12084 16304 12096
rect 15795 12056 16304 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 16669 12087 16727 12093
rect 16669 12053 16681 12087
rect 16715 12084 16727 12087
rect 18414 12084 18420 12096
rect 16715 12056 18420 12084
rect 16715 12053 16727 12056
rect 16669 12047 16727 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18524 12084 18552 12124
rect 18690 12112 18696 12164
rect 18748 12152 18754 12164
rect 19426 12152 19432 12164
rect 18748 12124 19432 12152
rect 18748 12112 18754 12124
rect 19426 12112 19432 12124
rect 19484 12112 19490 12164
rect 20714 12112 20720 12164
rect 20772 12112 20778 12164
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24946 12152 24952 12164
rect 23891 12124 24952 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24946 12112 24952 12124
rect 25004 12112 25010 12164
rect 18874 12084 18880 12096
rect 18524 12056 18880 12084
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19300 12056 19625 12084
rect 19300 12044 19306 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 20346 12084 20352 12096
rect 19852 12056 20352 12084
rect 19852 12044 19858 12056
rect 20346 12044 20352 12056
rect 20404 12084 20410 12096
rect 22189 12087 22247 12093
rect 22189 12084 22201 12087
rect 20404 12056 22201 12084
rect 20404 12044 20410 12056
rect 22189 12053 22201 12056
rect 22235 12053 22247 12087
rect 22189 12047 22247 12053
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 5408 11852 8892 11880
rect 5408 11840 5414 11852
rect 8864 11812 8892 11852
rect 9030 11840 9036 11892
rect 9088 11840 9094 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9732 11852 9873 11880
rect 9732 11840 9738 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 11931 11852 12664 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 9493 11815 9551 11821
rect 9493 11812 9505 11815
rect 8864 11784 9505 11812
rect 9493 11781 9505 11784
rect 9539 11812 9551 11815
rect 10226 11812 10232 11824
rect 9539 11784 10232 11812
rect 9539 11781 9551 11784
rect 9493 11775 9551 11781
rect 10226 11772 10232 11784
rect 10284 11772 10290 11824
rect 10321 11815 10379 11821
rect 10321 11781 10333 11815
rect 10367 11812 10379 11815
rect 12636 11812 12664 11852
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 12768 11852 13093 11880
rect 12768 11840 12774 11852
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 13081 11843 13139 11849
rect 13449 11883 13507 11889
rect 13449 11849 13461 11883
rect 13495 11880 13507 11883
rect 13538 11880 13544 11892
rect 13495 11852 13544 11880
rect 13495 11849 13507 11852
rect 13449 11843 13507 11849
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 14240 11852 14289 11880
rect 14240 11840 14246 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 16942 11880 16948 11892
rect 14277 11843 14335 11849
rect 15028 11852 16948 11880
rect 15028 11824 15056 11852
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 17092 11852 17325 11880
rect 17092 11840 17098 11852
rect 17313 11849 17325 11852
rect 17359 11849 17371 11883
rect 17313 11843 17371 11849
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11849 18107 11883
rect 18049 11843 18107 11849
rect 12802 11812 12808 11824
rect 10367 11784 12572 11812
rect 12636 11784 12808 11812
rect 10367 11781 10379 11784
rect 10321 11775 10379 11781
rect 9122 11744 9128 11756
rect 8694 11716 9128 11744
rect 9122 11704 9128 11716
rect 9180 11744 9186 11756
rect 9398 11744 9404 11756
rect 9180 11716 9404 11744
rect 9180 11704 9186 11716
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 11609 11747 11667 11753
rect 11609 11713 11621 11747
rect 11655 11744 11667 11747
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 11655 11716 12265 11744
rect 11655 11713 11667 11716
rect 11609 11707 11667 11713
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 7561 11679 7619 11685
rect 7331 11648 7420 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 7392 11540 7420 11648
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 7607 11648 10425 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 10413 11645 10425 11648
rect 10459 11676 10471 11679
rect 11054 11676 11060 11688
rect 10459 11648 11060 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 12268 11676 12296 11707
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12544 11744 12572 11784
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 14366 11812 14372 11824
rect 12912 11784 14372 11812
rect 12912 11744 12940 11784
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 15010 11812 15016 11824
rect 14660 11784 15016 11812
rect 14660 11753 14688 11784
rect 15010 11772 15016 11784
rect 15068 11772 15074 11824
rect 15194 11772 15200 11824
rect 15252 11812 15258 11824
rect 17678 11812 17684 11824
rect 15252 11784 17684 11812
rect 15252 11772 15258 11784
rect 17678 11772 17684 11784
rect 17736 11772 17742 11824
rect 18064 11812 18092 11843
rect 18414 11840 18420 11892
rect 18472 11840 18478 11892
rect 21358 11880 21364 11892
rect 19352 11852 21364 11880
rect 19352 11821 19380 11852
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 21637 11883 21695 11889
rect 21637 11849 21649 11883
rect 21683 11880 21695 11883
rect 22002 11880 22008 11892
rect 21683 11852 22008 11880
rect 21683 11849 21695 11852
rect 21637 11843 21695 11849
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 19337 11815 19395 11821
rect 18064 11784 19012 11812
rect 12544 11716 12940 11744
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11713 14703 11747
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 14645 11707 14703 11713
rect 15028 11716 17233 11744
rect 12268 11648 12388 11676
rect 12360 11620 12388 11648
rect 12434 11636 12440 11688
rect 12492 11636 12498 11688
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 12676 11648 13553 11676
rect 12676 11636 12682 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 13722 11636 13728 11688
rect 13780 11636 13786 11688
rect 14734 11636 14740 11688
rect 14792 11636 14798 11688
rect 14918 11636 14924 11688
rect 14976 11636 14982 11688
rect 12342 11568 12348 11620
rect 12400 11568 12406 11620
rect 12710 11568 12716 11620
rect 12768 11608 12774 11620
rect 15028 11608 15056 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 18984 11744 19012 11784
rect 19337 11781 19349 11815
rect 19383 11781 19395 11815
rect 19337 11775 19395 11781
rect 19978 11772 19984 11824
rect 20036 11772 20042 11824
rect 20070 11772 20076 11824
rect 20128 11812 20134 11824
rect 20622 11812 20628 11824
rect 20128 11784 20628 11812
rect 20128 11772 20134 11784
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 21269 11815 21327 11821
rect 21269 11781 21281 11815
rect 21315 11812 21327 11815
rect 21726 11812 21732 11824
rect 21315 11784 21732 11812
rect 21315 11781 21327 11784
rect 21269 11775 21327 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 19996 11744 20024 11772
rect 18984 11716 20024 11744
rect 20257 11747 20315 11753
rect 17221 11707 17279 11713
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20530 11744 20536 11756
rect 20303 11716 20536 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 23934 11744 23940 11756
rect 22327 11716 23940 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 23934 11704 23940 11716
rect 23992 11704 23998 11756
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24946 11744 24952 11756
rect 24167 11716 24952 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11676 15623 11679
rect 16022 11676 16028 11688
rect 15611 11648 16028 11676
rect 15611 11645 15623 11648
rect 15565 11639 15623 11645
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16724 11648 17417 11676
rect 16724 11636 16730 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 17770 11636 17776 11688
rect 17828 11676 17834 11688
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17828 11648 18521 11676
rect 17828 11636 17834 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11676 18751 11679
rect 19794 11676 19800 11688
rect 18739 11648 19800 11676
rect 18739 11645 18751 11648
rect 18693 11639 18751 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20036 11648 20729 11676
rect 20036 11636 20042 11648
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 24210 11676 24216 11688
rect 20956 11648 24216 11676
rect 20956 11636 20962 11648
rect 24210 11636 24216 11648
rect 24268 11636 24274 11688
rect 12768 11580 15056 11608
rect 16853 11611 16911 11617
rect 12768 11568 12774 11580
rect 16853 11577 16865 11611
rect 16899 11608 16911 11611
rect 20162 11608 20168 11620
rect 16899 11580 20168 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 20162 11568 20168 11580
rect 20220 11568 20226 11620
rect 20346 11568 20352 11620
rect 20404 11608 20410 11620
rect 22278 11608 22284 11620
rect 20404 11580 22284 11608
rect 20404 11568 20410 11580
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 8294 11540 8300 11552
rect 7392 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10134 11540 10140 11552
rect 9456 11512 10140 11540
rect 9456 11500 9462 11512
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 11238 11500 11244 11552
rect 11296 11500 11302 11552
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15289 11543 15347 11549
rect 15289 11540 15301 11543
rect 15068 11512 15301 11540
rect 15068 11500 15074 11512
rect 15289 11509 15301 11512
rect 15335 11509 15347 11543
rect 15289 11503 15347 11509
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 15654 11540 15660 11552
rect 15528 11512 15660 11540
rect 15528 11500 15534 11512
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 19334 11540 19340 11552
rect 16080 11512 19340 11540
rect 16080 11500 16086 11512
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 19794 11540 19800 11552
rect 19475 11512 19800 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 22002 11540 22008 11552
rect 20680 11512 22008 11540
rect 20680 11500 20686 11512
rect 22002 11500 22008 11512
rect 22060 11540 22066 11552
rect 25774 11540 25780 11552
rect 22060 11512 25780 11540
rect 22060 11500 22066 11512
rect 25774 11500 25780 11512
rect 25832 11500 25838 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7248 11308 10548 11336
rect 7248 11296 7254 11308
rect 10520 11268 10548 11308
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 12621 11339 12679 11345
rect 12621 11336 12633 11339
rect 10652 11308 12633 11336
rect 10652 11296 10658 11308
rect 12621 11305 12633 11308
rect 12667 11305 12679 11339
rect 15378 11336 15384 11348
rect 12621 11299 12679 11305
rect 14200 11308 15384 11336
rect 11238 11268 11244 11280
rect 10520 11240 11244 11268
rect 11238 11228 11244 11240
rect 11296 11228 11302 11280
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 12802 11268 12808 11280
rect 11471 11240 12808 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 13538 11268 13544 11280
rect 12952 11240 13544 11268
rect 12952 11228 12958 11240
rect 13538 11228 13544 11240
rect 13596 11268 13602 11280
rect 13725 11271 13783 11277
rect 13725 11268 13737 11271
rect 13596 11240 13737 11268
rect 13596 11228 13602 11240
rect 13725 11237 13737 11240
rect 13771 11237 13783 11271
rect 13725 11231 13783 11237
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 11882 11200 11888 11212
rect 9447 11172 11888 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 11882 11160 11888 11172
rect 11940 11200 11946 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11940 11172 11989 11200
rect 11940 11160 11946 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 11977 11163 12035 11169
rect 12406 11172 13277 11200
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 12406 11132 12434 11172
rect 13265 11169 13277 11172
rect 13311 11200 13323 11203
rect 13630 11200 13636 11212
rect 13311 11172 13636 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 11112 11104 12434 11132
rect 12989 11135 13047 11141
rect 11112 11092 11118 11104
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 14200 11132 14228 11308
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 17589 11339 17647 11345
rect 17589 11336 17601 11339
rect 15712 11308 17601 11336
rect 15712 11296 15718 11308
rect 17589 11305 17601 11308
rect 17635 11336 17647 11339
rect 17635 11308 18092 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 16666 11228 16672 11280
rect 16724 11228 16730 11280
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 16942 11200 16948 11212
rect 14967 11172 16948 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17770 11160 17776 11212
rect 17828 11160 17834 11212
rect 13035 11104 14228 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16816 11104 17141 11132
rect 16816 11092 16822 11104
rect 17129 11101 17141 11104
rect 17175 11132 17187 11135
rect 17175 11104 18000 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 7098 11064 7104 11076
rect 4212 11036 7104 11064
rect 4212 11024 4218 11036
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 10134 11024 10140 11076
rect 10192 11024 10198 11076
rect 11885 11067 11943 11073
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 12894 11064 12900 11076
rect 11931 11036 12900 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 13081 11067 13139 11073
rect 13081 11033 13093 11067
rect 13127 11064 13139 11067
rect 15102 11064 15108 11076
rect 13127 11036 15108 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 15194 11024 15200 11076
rect 15252 11024 15258 11076
rect 16482 11064 16488 11076
rect 16422 11036 16488 11064
rect 16482 11024 16488 11036
rect 16540 11064 16546 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 16540 11036 16957 11064
rect 16540 11024 16546 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 16945 11027 17003 11033
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10870 10996 10876 11008
rect 9732 10968 10876 10996
rect 9732 10956 9738 10968
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 11238 10956 11244 11008
rect 11296 10996 11302 11008
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 11296 10968 11805 10996
rect 11296 10956 11302 10968
rect 11793 10965 11805 10968
rect 11839 10996 11851 10999
rect 12250 10996 12256 11008
rect 11839 10968 12256 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 14274 10956 14280 11008
rect 14332 10956 14338 11008
rect 14366 10956 14372 11008
rect 14424 10996 14430 11008
rect 17862 10996 17868 11008
rect 14424 10968 17868 10996
rect 14424 10956 14430 10968
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 17972 10996 18000 11104
rect 18064 11064 18092 11308
rect 20162 11296 20168 11348
rect 20220 11336 20226 11348
rect 20622 11336 20628 11348
rect 20220 11308 20628 11336
rect 20220 11296 20226 11308
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 21545 11339 21603 11345
rect 21545 11305 21557 11339
rect 21591 11336 21603 11339
rect 22462 11336 22468 11348
rect 21591 11308 22468 11336
rect 21591 11305 21603 11308
rect 21545 11299 21603 11305
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 22830 11296 22836 11348
rect 22888 11336 22894 11348
rect 25041 11339 25099 11345
rect 25041 11336 25053 11339
rect 22888 11308 25053 11336
rect 22888 11296 22894 11308
rect 25041 11305 25053 11308
rect 25087 11305 25099 11339
rect 25041 11299 25099 11305
rect 18141 11271 18199 11277
rect 18141 11237 18153 11271
rect 18187 11268 18199 11271
rect 19518 11268 19524 11280
rect 18187 11240 19524 11268
rect 18187 11237 18199 11240
rect 18141 11231 18199 11237
rect 19518 11228 19524 11240
rect 19576 11228 19582 11280
rect 19613 11271 19671 11277
rect 19613 11237 19625 11271
rect 19659 11268 19671 11271
rect 21818 11268 21824 11280
rect 19659 11240 21824 11268
rect 19659 11237 19671 11240
rect 19613 11231 19671 11237
rect 21818 11228 21824 11240
rect 21876 11228 21882 11280
rect 22002 11228 22008 11280
rect 22060 11268 22066 11280
rect 22097 11271 22155 11277
rect 22097 11268 22109 11271
rect 22060 11240 22109 11268
rect 22060 11228 22066 11240
rect 22097 11237 22109 11240
rect 22143 11237 22155 11271
rect 22097 11231 22155 11237
rect 22278 11228 22284 11280
rect 22336 11268 22342 11280
rect 25590 11268 25596 11280
rect 22336 11240 25596 11268
rect 22336 11228 22342 11240
rect 25590 11228 25596 11240
rect 25648 11228 25654 11280
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 19426 11200 19432 11212
rect 18831 11172 19432 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 20257 11203 20315 11209
rect 20257 11169 20269 11203
rect 20303 11169 20315 11203
rect 20257 11163 20315 11169
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 19150 11132 19156 11144
rect 18647 11104 19156 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 19150 11092 19156 11104
rect 19208 11132 19214 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 19208 11104 19257 11132
rect 19208 11092 19214 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19978 11092 19984 11144
rect 20036 11092 20042 11144
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 18064 11036 18521 11064
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 20272 11064 20300 11163
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 21085 11203 21143 11209
rect 21085 11200 21097 11203
rect 21048 11172 21097 11200
rect 21048 11160 21054 11172
rect 21085 11169 21097 11172
rect 21131 11169 21143 11203
rect 21085 11163 21143 11169
rect 21910 11160 21916 11212
rect 21968 11200 21974 11212
rect 21968 11172 25268 11200
rect 21968 11160 21974 11172
rect 20622 11092 20628 11144
rect 20680 11132 20686 11144
rect 21729 11135 21787 11141
rect 21729 11132 21741 11135
rect 20680 11104 21741 11132
rect 20680 11092 20686 11104
rect 21729 11101 21741 11104
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11132 22891 11135
rect 23290 11132 23296 11144
rect 22879 11104 23296 11132
rect 22879 11101 22891 11104
rect 22833 11095 22891 11101
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 25240 11141 25268 11172
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11101 25283 11135
rect 25225 11095 25283 11101
rect 20346 11064 20352 11076
rect 18509 11027 18567 11033
rect 18616 11036 20208 11064
rect 20272 11036 20352 11064
rect 18616 10996 18644 11036
rect 17972 10968 18644 10996
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 20073 10999 20131 11005
rect 20073 10996 20085 10999
rect 20036 10968 20085 10996
rect 20036 10956 20042 10968
rect 20073 10965 20085 10968
rect 20119 10965 20131 10999
rect 20180 10996 20208 11036
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 20901 11067 20959 11073
rect 20901 11033 20913 11067
rect 20947 11064 20959 11067
rect 21266 11064 21272 11076
rect 20947 11036 21272 11064
rect 20947 11033 20959 11036
rect 20901 11027 20959 11033
rect 21266 11024 21272 11036
rect 21324 11064 21330 11076
rect 22278 11064 22284 11076
rect 21324 11036 22284 11064
rect 21324 11024 21330 11036
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 23382 11024 23388 11076
rect 23440 11064 23446 11076
rect 23569 11067 23627 11073
rect 23569 11064 23581 11067
rect 23440 11036 23581 11064
rect 23440 11024 23446 11036
rect 23569 11033 23581 11036
rect 23615 11033 23627 11067
rect 23569 11027 23627 11033
rect 21450 10996 21456 11008
rect 20180 10968 21456 10996
rect 20073 10959 20131 10965
rect 21450 10956 21456 10968
rect 21508 10996 21514 11008
rect 24026 10996 24032 11008
rect 21508 10968 24032 10996
rect 21508 10956 21514 10968
rect 24026 10956 24032 10968
rect 24084 10956 24090 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 12158 10792 12164 10804
rect 9999 10764 12164 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12345 10795 12403 10801
rect 12345 10761 12357 10795
rect 12391 10761 12403 10795
rect 12345 10755 12403 10761
rect 8202 10724 8208 10736
rect 7852 10696 8208 10724
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7852 10461 7880 10696
rect 8202 10684 8208 10696
rect 8260 10724 8266 10736
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 8260 10696 8493 10724
rect 8260 10684 8266 10696
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 8481 10687 8539 10693
rect 10134 10656 10140 10668
rect 9614 10628 10140 10656
rect 10134 10616 10140 10628
rect 10192 10656 10198 10668
rect 12360 10656 12388 10755
rect 12802 10752 12808 10804
rect 12860 10752 12866 10804
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 13906 10792 13912 10804
rect 13863 10764 13912 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 14185 10795 14243 10801
rect 14185 10761 14197 10795
rect 14231 10792 14243 10795
rect 14366 10792 14372 10804
rect 14231 10764 14372 10792
rect 14231 10761 14243 10764
rect 14185 10755 14243 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15562 10752 15568 10804
rect 15620 10752 15626 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16758 10792 16764 10804
rect 15979 10764 16764 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 18233 10795 18291 10801
rect 16899 10764 18184 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 12713 10727 12771 10733
rect 12713 10693 12725 10727
rect 12759 10724 12771 10727
rect 14274 10724 14280 10736
rect 12759 10696 14280 10724
rect 12759 10693 12771 10696
rect 12713 10687 12771 10693
rect 14274 10684 14280 10696
rect 14332 10684 14338 10736
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 14884 10696 17172 10724
rect 14884 10684 14890 10696
rect 10192 10628 10456 10656
rect 12360 10628 16620 10656
rect 10192 10616 10198 10628
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7156 10424 7849 10452
rect 7156 10412 7162 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8220 10452 8248 10551
rect 8294 10452 8300 10464
rect 8220 10424 8300 10452
rect 7837 10415 7895 10421
rect 8294 10412 8300 10424
rect 8352 10452 8358 10464
rect 9122 10452 9128 10464
rect 8352 10424 9128 10452
rect 8352 10412 8358 10424
rect 9122 10412 9128 10424
rect 9180 10452 9186 10464
rect 9582 10452 9588 10464
rect 9180 10424 9588 10452
rect 9180 10412 9186 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 10428 10461 10456 10628
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10588 11759 10591
rect 12802 10588 12808 10600
rect 11747 10560 12808 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 12912 10520 12940 10551
rect 14274 10548 14280 10600
rect 14332 10548 14338 10600
rect 14458 10548 14464 10600
rect 14516 10548 14522 10600
rect 15378 10548 15384 10600
rect 15436 10588 15442 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15436 10560 16037 10588
rect 15436 10548 15442 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10588 16267 10591
rect 16482 10588 16488 10600
rect 16255 10560 16488 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 14476 10520 14504 10548
rect 16224 10520 16252 10551
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 16592 10588 16620 10628
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 17144 10656 17172 10696
rect 17586 10684 17592 10736
rect 17644 10684 17650 10736
rect 18156 10724 18184 10764
rect 18233 10761 18245 10795
rect 18279 10792 18291 10795
rect 22002 10792 22008 10804
rect 18279 10764 22008 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 22833 10795 22891 10801
rect 22833 10761 22845 10795
rect 22879 10792 22891 10795
rect 23198 10792 23204 10804
rect 22879 10764 23204 10792
rect 22879 10761 22891 10764
rect 22833 10755 22891 10761
rect 23198 10752 23204 10764
rect 23256 10792 23262 10804
rect 23256 10764 23520 10792
rect 23256 10752 23262 10764
rect 19518 10724 19524 10736
rect 18156 10696 19524 10724
rect 19518 10684 19524 10696
rect 19576 10684 19582 10736
rect 20070 10724 20076 10736
rect 19996 10696 20076 10724
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 17144 10628 18429 10656
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 19996 10656 20024 10696
rect 20070 10684 20076 10696
rect 20128 10684 20134 10736
rect 21082 10684 21088 10736
rect 21140 10684 21146 10736
rect 21174 10684 21180 10736
rect 21232 10684 21238 10736
rect 22465 10727 22523 10733
rect 22465 10724 22477 10727
rect 21284 10696 22477 10724
rect 21284 10656 21312 10696
rect 22465 10693 22477 10696
rect 22511 10693 22523 10727
rect 22465 10687 22523 10693
rect 22554 10684 22560 10736
rect 22612 10724 22618 10736
rect 23385 10727 23443 10733
rect 23385 10724 23397 10727
rect 22612 10696 23397 10724
rect 22612 10684 22618 10696
rect 23385 10693 23397 10696
rect 23431 10693 23443 10727
rect 23492 10724 23520 10764
rect 23842 10724 23848 10736
rect 23492 10696 23848 10724
rect 23385 10687 23443 10693
rect 23842 10684 23848 10696
rect 23900 10684 23906 10736
rect 19935 10628 20024 10656
rect 20088 10628 21312 10656
rect 22189 10659 22247 10665
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 18322 10588 18328 10600
rect 16592 10560 18328 10588
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 18782 10520 18788 10532
rect 10928 10492 12940 10520
rect 13096 10492 16252 10520
rect 17236 10492 18788 10520
rect 10928 10480 10934 10492
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10452 10471 10455
rect 10962 10452 10968 10464
rect 10459 10424 10968 10452
rect 10459 10421 10471 10424
rect 10413 10415 10471 10421
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11238 10412 11244 10464
rect 11296 10412 11302 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 13096 10452 13124 10492
rect 12492 10424 13124 10452
rect 12492 10412 12498 10424
rect 13446 10412 13452 10464
rect 13504 10412 13510 10464
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15378 10452 15384 10464
rect 15335 10424 15384 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15378 10412 15384 10424
rect 15436 10452 15442 10464
rect 17236 10452 17264 10492
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 19076 10520 19104 10619
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19981 10591 20039 10597
rect 19392 10560 19748 10588
rect 19392 10548 19398 10560
rect 19720 10520 19748 10560
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 20088 10588 20116 10628
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22235 10628 22600 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 20027 10560 20116 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 19996 10520 20024 10551
rect 20162 10548 20168 10600
rect 20220 10548 20226 10600
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 21266 10588 21272 10600
rect 20772 10560 21272 10588
rect 20772 10548 20778 10560
rect 21266 10548 21272 10560
rect 21324 10548 21330 10600
rect 22572 10588 22600 10628
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 23109 10659 23167 10665
rect 23109 10656 23121 10659
rect 22704 10628 23121 10656
rect 22704 10616 22710 10628
rect 23109 10625 23121 10628
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 22738 10588 22744 10600
rect 22572 10560 22744 10588
rect 22738 10548 22744 10560
rect 22796 10548 22802 10600
rect 19076 10492 19656 10520
rect 19720 10492 20024 10520
rect 15436 10424 17264 10452
rect 15436 10412 15442 10424
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 17368 10424 17693 10452
rect 17368 10412 17374 10424
rect 17681 10421 17693 10424
rect 17727 10421 17739 10455
rect 17681 10415 17739 10421
rect 18414 10412 18420 10464
rect 18472 10452 18478 10464
rect 18877 10455 18935 10461
rect 18877 10452 18889 10455
rect 18472 10424 18889 10452
rect 18472 10412 18478 10424
rect 18877 10421 18889 10424
rect 18923 10421 18935 10455
rect 18877 10415 18935 10421
rect 19518 10412 19524 10464
rect 19576 10412 19582 10464
rect 19628 10452 19656 10492
rect 21358 10480 21364 10532
rect 21416 10520 21422 10532
rect 22005 10523 22063 10529
rect 22005 10520 22017 10523
rect 21416 10492 22017 10520
rect 21416 10480 21422 10492
rect 22005 10489 22017 10492
rect 22051 10489 22063 10523
rect 22005 10483 22063 10489
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 19628 10424 20729 10452
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 20717 10415 20775 10421
rect 23382 10412 23388 10464
rect 23440 10452 23446 10464
rect 24857 10455 24915 10461
rect 24857 10452 24869 10455
rect 23440 10424 24869 10452
rect 23440 10412 23446 10424
rect 24857 10421 24869 10424
rect 24903 10421 24915 10455
rect 24857 10415 24915 10421
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8260 10220 11008 10248
rect 8260 10208 8266 10220
rect 10980 10180 11008 10220
rect 11054 10208 11060 10260
rect 11112 10208 11118 10260
rect 11606 10208 11612 10260
rect 11664 10208 11670 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12124 10220 12817 10248
rect 12124 10208 12130 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 14550 10208 14556 10260
rect 14608 10208 14614 10260
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 15657 10251 15715 10257
rect 15657 10248 15669 10251
rect 14976 10220 15669 10248
rect 14976 10208 14982 10220
rect 15657 10217 15669 10220
rect 15703 10248 15715 10251
rect 20438 10248 20444 10260
rect 15703 10220 20444 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 21266 10208 21272 10260
rect 21324 10248 21330 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 21324 10220 22293 10248
rect 21324 10208 21330 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 24302 10248 24308 10260
rect 22281 10211 22339 10217
rect 22388 10220 24308 10248
rect 10980 10152 12296 10180
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9582 10112 9588 10124
rect 9355 10084 9588 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 12158 10072 12164 10124
rect 12216 10072 12222 10124
rect 12268 10112 12296 10152
rect 12434 10140 12440 10192
rect 12492 10180 12498 10192
rect 17034 10180 17040 10192
rect 12492 10152 17040 10180
rect 12492 10140 12498 10152
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 20346 10180 20352 10192
rect 17920 10152 20352 10180
rect 17920 10140 17926 10152
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 21818 10140 21824 10192
rect 21876 10180 21882 10192
rect 22388 10180 22416 10220
rect 24302 10208 24308 10220
rect 24360 10208 24366 10260
rect 24578 10208 24584 10260
rect 24636 10208 24642 10260
rect 21876 10152 22416 10180
rect 21876 10140 21882 10152
rect 22554 10140 22560 10192
rect 22612 10180 22618 10192
rect 23842 10180 23848 10192
rect 22612 10152 23848 10180
rect 22612 10140 22618 10152
rect 23842 10140 23848 10152
rect 23900 10180 23906 10192
rect 24118 10180 24124 10192
rect 23900 10152 24124 10180
rect 23900 10140 23906 10152
rect 24118 10140 24124 10152
rect 24176 10140 24182 10192
rect 13449 10115 13507 10121
rect 12268 10084 13400 10112
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12860 10016 13185 10044
rect 12860 10004 12866 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13372 10044 13400 10084
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13630 10112 13636 10124
rect 13495 10084 13636 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10112 14335 10115
rect 14458 10112 14464 10124
rect 14323 10084 14464 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 14292 10044 14320 10075
rect 14458 10072 14464 10084
rect 14516 10112 14522 10124
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 14516 10084 15117 10112
rect 14516 10072 14522 10084
rect 15105 10081 15117 10084
rect 15151 10112 15163 10115
rect 15838 10112 15844 10124
rect 15151 10084 15844 10112
rect 15151 10081 15163 10084
rect 15105 10075 15163 10081
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 17770 10112 17776 10124
rect 16868 10084 17776 10112
rect 13372 10016 14320 10044
rect 13173 10007 13231 10013
rect 14918 10004 14924 10056
rect 14976 10004 14982 10056
rect 16868 10044 16896 10084
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18012 10084 18276 10112
rect 18012 10072 18018 10084
rect 15028 10016 16896 10044
rect 18248 10044 18276 10084
rect 18322 10072 18328 10124
rect 18380 10112 18386 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 18380 10084 18429 10112
rect 18380 10072 18386 10084
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 18417 10075 18475 10081
rect 18601 10115 18659 10121
rect 18601 10081 18613 10115
rect 18647 10112 18659 10115
rect 18782 10112 18788 10124
rect 18647 10084 18788 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19576 10084 22094 10112
rect 19576 10072 19582 10084
rect 18248 10016 18368 10044
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9548 9948 9597 9976
rect 9548 9936 9554 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 10962 9976 10968 9988
rect 10810 9948 10968 9976
rect 9585 9939 9643 9945
rect 10962 9936 10968 9948
rect 11020 9976 11026 9988
rect 11514 9976 11520 9988
rect 11020 9948 11520 9976
rect 11020 9936 11026 9948
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 11977 9979 12035 9985
rect 11977 9945 11989 9979
rect 12023 9976 12035 9979
rect 13906 9976 13912 9988
rect 12023 9948 13912 9976
rect 12023 9945 12035 9948
rect 11977 9939 12035 9945
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 12066 9868 12072 9920
rect 12124 9868 12130 9920
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9908 13323 9911
rect 13354 9908 13360 9920
rect 13311 9880 13360 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 13354 9868 13360 9880
rect 13412 9908 13418 9920
rect 13538 9908 13544 9920
rect 13412 9880 13544 9908
rect 13412 9868 13418 9880
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 13817 9911 13875 9917
rect 13817 9877 13829 9911
rect 13863 9908 13875 9911
rect 14734 9908 14740 9920
rect 13863 9880 14740 9908
rect 13863 9877 13875 9880
rect 13817 9871 13875 9877
rect 14734 9868 14740 9880
rect 14792 9908 14798 9920
rect 15028 9917 15056 10016
rect 16114 9936 16120 9988
rect 16172 9936 16178 9988
rect 16850 9936 16856 9988
rect 16908 9936 16914 9988
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14792 9880 15025 9908
rect 14792 9868 14798 9880
rect 15013 9877 15025 9880
rect 15059 9877 15071 9911
rect 15013 9871 15071 9877
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16816 9880 16957 9908
rect 16816 9868 16822 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 17957 9911 18015 9917
rect 17957 9877 17969 9911
rect 18003 9908 18015 9911
rect 18230 9908 18236 9920
rect 18003 9880 18236 9908
rect 18003 9877 18015 9880
rect 17957 9871 18015 9877
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18340 9917 18368 10016
rect 18874 10004 18880 10056
rect 18932 10044 18938 10056
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 18932 10016 20545 10044
rect 18932 10004 18938 10016
rect 20533 10013 20545 10016
rect 20579 10013 20591 10047
rect 22066 10044 22094 10084
rect 22370 10072 22376 10124
rect 22428 10112 22434 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 22428 10084 23305 10112
rect 22428 10072 22434 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23382 10072 23388 10124
rect 23440 10072 23446 10124
rect 22066 10016 22692 10044
rect 20533 10007 20591 10013
rect 19521 9979 19579 9985
rect 19521 9945 19533 9979
rect 19567 9976 19579 9979
rect 19886 9976 19892 9988
rect 19567 9948 19892 9976
rect 19567 9945 19579 9948
rect 19521 9939 19579 9945
rect 19886 9936 19892 9948
rect 19944 9936 19950 9988
rect 20714 9936 20720 9988
rect 20772 9976 20778 9988
rect 20809 9979 20867 9985
rect 20809 9976 20821 9979
rect 20772 9948 20821 9976
rect 20772 9936 20778 9948
rect 20809 9945 20821 9948
rect 20855 9945 20867 9979
rect 22554 9976 22560 9988
rect 22034 9948 22560 9976
rect 20809 9939 20867 9945
rect 22554 9936 22560 9948
rect 22612 9936 22618 9988
rect 22664 9976 22692 10016
rect 22738 10004 22744 10056
rect 22796 10044 22802 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 22796 10016 23213 10044
rect 22796 10004 22802 10016
rect 23201 10013 23213 10016
rect 23247 10013 23259 10047
rect 23201 10007 23259 10013
rect 24670 10004 24676 10056
rect 24728 10044 24734 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 24728 10016 24777 10044
rect 24728 10004 24734 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 22664 9948 24716 9976
rect 24688 9920 24716 9948
rect 18325 9911 18383 9917
rect 18325 9877 18337 9911
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 18690 9868 18696 9920
rect 18748 9908 18754 9920
rect 18969 9911 19027 9917
rect 18969 9908 18981 9911
rect 18748 9880 18981 9908
rect 18748 9868 18754 9880
rect 18969 9877 18981 9880
rect 19015 9908 19027 9911
rect 19150 9908 19156 9920
rect 19015 9880 19156 9908
rect 19015 9877 19027 9880
rect 18969 9871 19027 9877
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19392 9880 19625 9908
rect 19392 9868 19398 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 19978 9868 19984 9920
rect 20036 9868 20042 9920
rect 20162 9868 20168 9920
rect 20220 9868 20226 9920
rect 20438 9868 20444 9920
rect 20496 9908 20502 9920
rect 21818 9908 21824 9920
rect 20496 9880 21824 9908
rect 20496 9868 20502 9880
rect 21818 9868 21824 9880
rect 21876 9868 21882 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22833 9911 22891 9917
rect 22833 9908 22845 9911
rect 22152 9880 22845 9908
rect 22152 9868 22158 9880
rect 22833 9877 22845 9880
rect 22879 9877 22891 9911
rect 22833 9871 22891 9877
rect 24670 9868 24676 9920
rect 24728 9868 24734 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 13446 9704 13452 9716
rect 12406 9676 13452 9704
rect 11514 9596 11520 9648
rect 11572 9636 11578 9648
rect 12406 9636 12434 9676
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 13906 9664 13912 9716
rect 13964 9664 13970 9716
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 17862 9704 17868 9716
rect 14608 9676 17868 9704
rect 14608 9664 14614 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 18506 9664 18512 9716
rect 18564 9704 18570 9716
rect 18564 9676 18920 9704
rect 18564 9664 18570 9676
rect 14277 9639 14335 9645
rect 11572 9608 12466 9636
rect 11572 9596 11578 9608
rect 14277 9605 14289 9639
rect 14323 9636 14335 9639
rect 15286 9636 15292 9648
rect 14323 9608 15292 9636
rect 14323 9605 14335 9608
rect 14277 9599 14335 9605
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 16117 9639 16175 9645
rect 16117 9636 16129 9639
rect 15396 9608 16129 9636
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 15396 9568 15424 9608
rect 16117 9605 16129 9608
rect 16163 9605 16175 9639
rect 16117 9599 16175 9605
rect 14056 9540 15424 9568
rect 15473 9571 15531 9577
rect 14056 9528 14062 9540
rect 14384 9512 14412 9540
rect 15473 9537 15485 9571
rect 15519 9537 15531 9571
rect 18892 9568 18920 9676
rect 18966 9664 18972 9716
rect 19024 9704 19030 9716
rect 19024 9676 19472 9704
rect 19024 9664 19030 9676
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 19300 9608 19380 9636
rect 19300 9596 19306 9608
rect 15473 9531 15531 9537
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 12710 9500 12716 9512
rect 12023 9472 12716 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9500 13507 9503
rect 14090 9500 14096 9512
rect 13495 9472 14096 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14366 9460 14372 9512
rect 14424 9460 14430 9512
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 15102 9392 15108 9444
rect 15160 9392 15166 9444
rect 11330 9324 11336 9376
rect 11388 9324 11394 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 15378 9364 15384 9376
rect 13872 9336 15384 9364
rect 13872 9324 13878 9336
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15488 9364 15516 9531
rect 15562 9460 15568 9512
rect 15620 9460 15626 9512
rect 15746 9460 15752 9512
rect 15804 9460 15810 9512
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 17000 9472 17325 9500
rect 17000 9460 17006 9472
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9500 17647 9503
rect 18230 9500 18236 9512
rect 17635 9472 18236 9500
rect 17635 9469 17647 9472
rect 17589 9463 17647 9469
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18708 9500 18736 9554
rect 18892 9540 19288 9568
rect 18874 9500 18880 9512
rect 18708 9472 18880 9500
rect 18874 9460 18880 9472
rect 18932 9460 18938 9512
rect 19260 9432 19288 9540
rect 19352 9500 19380 9608
rect 19444 9592 19472 9676
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 20162 9704 20168 9716
rect 19576 9676 20168 9704
rect 19576 9664 19582 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 21082 9664 21088 9716
rect 21140 9704 21146 9716
rect 21818 9704 21824 9716
rect 21140 9676 21824 9704
rect 21140 9664 21146 9676
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 22002 9704 22008 9716
rect 21928 9676 22008 9704
rect 21928 9636 21956 9676
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 22278 9664 22284 9716
rect 22336 9704 22342 9716
rect 24397 9707 24455 9713
rect 24397 9704 24409 9707
rect 22336 9676 24409 9704
rect 22336 9664 22342 9676
rect 24397 9673 24409 9676
rect 24443 9673 24455 9707
rect 24397 9667 24455 9673
rect 19812 9608 21956 9636
rect 19444 9568 19564 9592
rect 19812 9568 19840 9608
rect 19444 9564 19840 9568
rect 19536 9540 19840 9564
rect 20070 9528 20076 9580
rect 20128 9528 20134 9580
rect 19352 9472 20668 9500
rect 20162 9432 20168 9444
rect 19260 9404 20168 9432
rect 20162 9392 20168 9404
rect 20220 9392 20226 9444
rect 20640 9432 20668 9472
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 21174 9500 21180 9512
rect 20772 9472 21180 9500
rect 20772 9460 20778 9472
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 21818 9500 21824 9512
rect 21315 9472 21824 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 21910 9460 21916 9512
rect 21968 9500 21974 9512
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 21968 9472 22017 9500
rect 21968 9460 21974 9472
rect 22005 9469 22017 9472
rect 22051 9469 22063 9503
rect 22005 9463 22063 9469
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22646 9500 22652 9512
rect 22152 9472 22652 9500
rect 22152 9460 22158 9472
rect 22646 9460 22652 9472
rect 22704 9460 22710 9512
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23382 9500 23388 9512
rect 22971 9472 23388 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 24044 9500 24072 9554
rect 24394 9528 24400 9580
rect 24452 9568 24458 9580
rect 25041 9571 25099 9577
rect 25041 9568 25053 9571
rect 24452 9540 25053 9568
rect 24452 9528 24458 9540
rect 25041 9537 25053 9540
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 24118 9500 24124 9512
rect 24044 9472 24124 9500
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 20640 9404 22129 9432
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 15488 9336 16405 9364
rect 16393 9333 16405 9336
rect 16439 9364 16451 9367
rect 18690 9364 18696 9376
rect 16439 9336 18696 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 18690 9324 18696 9336
rect 18748 9324 18754 9376
rect 19058 9324 19064 9376
rect 19116 9324 19122 9376
rect 19242 9324 19248 9376
rect 19300 9364 19306 9376
rect 19426 9364 19432 9376
rect 19300 9336 19432 9364
rect 19300 9324 19306 9336
rect 19426 9324 19432 9336
rect 19484 9364 19490 9376
rect 19797 9367 19855 9373
rect 19797 9364 19809 9367
rect 19484 9336 19809 9364
rect 19484 9324 19490 9336
rect 19797 9333 19809 9336
rect 19843 9364 19855 9367
rect 19886 9364 19892 9376
rect 19843 9336 19892 9364
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 19886 9324 19892 9336
rect 19944 9364 19950 9376
rect 21634 9364 21640 9376
rect 19944 9336 21640 9364
rect 19944 9324 19950 9336
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 22101 9364 22129 9404
rect 24857 9367 24915 9373
rect 24857 9364 24869 9367
rect 22101 9336 24869 9364
rect 24857 9333 24869 9336
rect 24903 9333 24915 9367
rect 24857 9327 24915 9333
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 12066 9120 12072 9172
rect 12124 9160 12130 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 12124 9132 14289 9160
rect 12124 9120 12130 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 19058 9160 19064 9172
rect 15068 9132 19064 9160
rect 15068 9120 15074 9132
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 19260 9132 20944 9160
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 10744 9064 13001 9092
rect 10744 9052 10750 9064
rect 12989 9061 13001 9064
rect 13035 9061 13047 9095
rect 12989 9055 13047 9061
rect 13722 9052 13728 9104
rect 13780 9092 13786 9104
rect 15933 9095 15991 9101
rect 15933 9092 15945 9095
rect 13780 9064 15945 9092
rect 13780 9052 13786 9064
rect 15933 9061 15945 9064
rect 15979 9061 15991 9095
rect 15933 9055 15991 9061
rect 17221 9095 17279 9101
rect 17221 9061 17233 9095
rect 17267 9092 17279 9095
rect 19260 9092 19288 9132
rect 17267 9064 19288 9092
rect 19337 9095 19395 9101
rect 17267 9061 17279 9064
rect 17221 9055 17279 9061
rect 19337 9061 19349 9095
rect 19383 9092 19395 9095
rect 19426 9092 19432 9104
rect 19383 9064 19432 9092
rect 19383 9061 19395 9064
rect 19337 9055 19395 9061
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 11054 9024 11060 9036
rect 9171 8996 11060 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 11054 8984 11060 8996
rect 11112 9024 11118 9036
rect 11698 9024 11704 9036
rect 11112 8996 11704 9024
rect 11112 8984 11118 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 14829 9027 14887 9033
rect 14829 9024 14841 9027
rect 14516 8996 14841 9024
rect 14516 8984 14522 8996
rect 14829 8993 14841 8996
rect 14875 8993 14887 9027
rect 14829 8987 14887 8993
rect 15286 8984 15292 9036
rect 15344 8984 15350 9036
rect 16482 8984 16488 9036
rect 16540 8984 16546 9036
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 15838 8956 15844 8968
rect 13495 8928 15844 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 17236 8956 17264 9055
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 20916 9092 20944 9132
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 21361 9163 21419 9169
rect 21361 9160 21373 9163
rect 21232 9132 21373 9160
rect 21232 9120 21238 9132
rect 21361 9129 21373 9132
rect 21407 9129 21419 9163
rect 21361 9123 21419 9129
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 23290 9160 23296 9172
rect 22888 9132 23296 9160
rect 22888 9120 22894 9132
rect 23290 9120 23296 9132
rect 23348 9120 23354 9172
rect 23934 9120 23940 9172
rect 23992 9160 23998 9172
rect 24581 9163 24639 9169
rect 24581 9160 24593 9163
rect 23992 9132 24593 9160
rect 23992 9120 23998 9132
rect 24581 9129 24593 9132
rect 24627 9129 24639 9163
rect 24581 9123 24639 9129
rect 21542 9092 21548 9104
rect 20916 9064 21548 9092
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 25041 9095 25099 9101
rect 25041 9092 25053 9095
rect 22756 9064 25053 9092
rect 18230 8984 18236 9036
rect 18288 9024 18294 9036
rect 19242 9024 19248 9036
rect 18288 8996 19248 9024
rect 18288 8984 18294 8996
rect 19242 8984 19248 8996
rect 19300 8984 19306 9036
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 9024 19671 9027
rect 20254 9024 20260 9036
rect 19659 8996 20260 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 20254 8984 20260 8996
rect 20312 8984 20318 9036
rect 20346 8984 20352 9036
rect 20404 9024 20410 9036
rect 22756 9024 22784 9064
rect 25041 9061 25053 9064
rect 25087 9061 25099 9095
rect 25041 9055 25099 9061
rect 20404 8996 21956 9024
rect 20404 8984 20410 8996
rect 16347 8928 17264 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 19518 8956 19524 8968
rect 18616 8928 19524 8956
rect 9401 8891 9459 8897
rect 9401 8857 9413 8891
rect 9447 8888 9459 8891
rect 9674 8888 9680 8900
rect 9447 8860 9680 8888
rect 9447 8857 9459 8860
rect 9401 8851 9459 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 11149 8891 11207 8897
rect 11149 8888 11161 8891
rect 10626 8860 11161 8888
rect 11149 8857 11161 8860
rect 11195 8888 11207 8891
rect 11330 8888 11336 8900
rect 11195 8860 11336 8888
rect 11195 8857 11207 8860
rect 11149 8851 11207 8857
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 12894 8888 12900 8900
rect 12584 8860 12900 8888
rect 12584 8848 12590 8860
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 13357 8891 13415 8897
rect 13357 8857 13369 8891
rect 13403 8888 13415 8891
rect 13998 8888 14004 8900
rect 13403 8860 14004 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13998 8848 14004 8860
rect 14056 8848 14062 8900
rect 14645 8891 14703 8897
rect 14645 8857 14657 8891
rect 14691 8888 14703 8891
rect 14918 8888 14924 8900
rect 14691 8860 14924 8888
rect 14691 8857 14703 8860
rect 14645 8851 14703 8857
rect 14918 8848 14924 8860
rect 14976 8888 14982 8900
rect 15378 8888 15384 8900
rect 14976 8860 15384 8888
rect 14976 8848 14982 8860
rect 15378 8848 15384 8860
rect 15436 8848 15442 8900
rect 15473 8891 15531 8897
rect 15473 8857 15485 8891
rect 15519 8888 15531 8891
rect 15562 8888 15568 8900
rect 15519 8860 15568 8888
rect 15519 8857 15531 8860
rect 15473 8851 15531 8857
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 10962 8820 10968 8832
rect 10919 8792 10968 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 12713 8823 12771 8829
rect 12713 8789 12725 8823
rect 12759 8820 12771 8823
rect 14458 8820 14464 8832
rect 12759 8792 14464 8820
rect 12759 8789 12771 8792
rect 12713 8783 12771 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 14608 8792 14749 8820
rect 14608 8780 14614 8792
rect 14737 8789 14749 8792
rect 14783 8789 14795 8823
rect 14737 8783 14795 8789
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 15160 8792 16405 8820
rect 15160 8780 15166 8792
rect 16393 8789 16405 8792
rect 16439 8820 16451 8823
rect 16945 8823 17003 8829
rect 16945 8820 16957 8823
rect 16439 8792 16957 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 16945 8789 16957 8792
rect 16991 8820 17003 8823
rect 18616 8820 18644 8928
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 21928 8965 21956 8996
rect 22664 8996 22784 9024
rect 21913 8959 21971 8965
rect 21913 8925 21925 8959
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 22554 8916 22560 8968
rect 22612 8956 22618 8968
rect 22664 8965 22692 8996
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 22612 8928 22661 8956
rect 22612 8916 22618 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 22649 8919 22707 8925
rect 22940 8928 24777 8956
rect 18693 8891 18751 8897
rect 18693 8857 18705 8891
rect 18739 8888 18751 8891
rect 18739 8860 19380 8888
rect 18739 8857 18751 8860
rect 18693 8851 18751 8857
rect 16991 8792 18644 8820
rect 19352 8820 19380 8860
rect 19426 8848 19432 8900
rect 19484 8888 19490 8900
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 19484 8860 19901 8888
rect 19484 8848 19490 8860
rect 19889 8857 19901 8860
rect 19935 8857 19947 8891
rect 21634 8888 21640 8900
rect 21114 8860 21640 8888
rect 19889 8851 19947 8857
rect 21634 8848 21640 8860
rect 21692 8848 21698 8900
rect 22462 8848 22468 8900
rect 22520 8888 22526 8900
rect 22940 8888 22968 8928
rect 24765 8925 24777 8928
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 22520 8860 22968 8888
rect 23845 8891 23903 8897
rect 22520 8848 22526 8860
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24946 8888 24952 8900
rect 23891 8860 24952 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 21174 8820 21180 8832
rect 19352 8792 21180 8820
rect 16991 8789 17003 8792
rect 16945 8783 17003 8789
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 21726 8780 21732 8832
rect 21784 8820 21790 8832
rect 22005 8823 22063 8829
rect 22005 8820 22017 8823
rect 21784 8792 22017 8820
rect 21784 8780 21790 8792
rect 22005 8789 22017 8792
rect 22051 8789 22063 8823
rect 22005 8783 22063 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 9916 8588 12848 8616
rect 9916 8576 9922 8588
rect 12820 8548 12848 8588
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 12952 8588 13952 8616
rect 12952 8576 12958 8588
rect 13814 8548 13820 8560
rect 12820 8520 13820 8548
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 13924 8557 13952 8588
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 15672 8588 23980 8616
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8517 13967 8551
rect 13909 8511 13967 8517
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 15010 8480 15016 8492
rect 11664 8452 15016 8480
rect 11664 8440 11670 8452
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8480 15163 8483
rect 15672 8480 15700 8588
rect 15746 8508 15752 8560
rect 15804 8548 15810 8560
rect 17586 8548 17592 8560
rect 15804 8520 17592 8548
rect 15804 8508 15810 8520
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 18690 8508 18696 8560
rect 18748 8548 18754 8560
rect 21269 8551 21327 8557
rect 18748 8520 20392 8548
rect 18748 8508 18754 8520
rect 15151 8452 15700 8480
rect 17405 8483 17463 8489
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17451 8452 18184 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8412 13231 8415
rect 13354 8412 13360 8424
rect 13219 8384 13360 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 13464 8384 14841 8412
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 4798 8344 4804 8356
rect 3844 8316 4804 8344
rect 3844 8304 3850 8316
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 11146 8344 11152 8356
rect 5316 8316 11152 8344
rect 5316 8304 5322 8316
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 13464 8344 13492 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 16114 8372 16120 8424
rect 16172 8372 16178 8424
rect 16761 8415 16819 8421
rect 16761 8381 16773 8415
rect 16807 8412 16819 8415
rect 17497 8415 17555 8421
rect 17497 8412 17509 8415
rect 16807 8384 17509 8412
rect 16807 8381 16819 8384
rect 16761 8375 16819 8381
rect 17497 8381 17509 8384
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 12584 8316 13492 8344
rect 12584 8304 12590 8316
rect 13998 8304 14004 8356
rect 14056 8304 14062 8356
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8344 14151 8347
rect 14642 8344 14648 8356
rect 14139 8316 14648 8344
rect 14139 8313 14151 8316
rect 14093 8307 14151 8313
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 17037 8347 17095 8353
rect 17037 8344 17049 8347
rect 15580 8316 17049 8344
rect 14016 8276 14044 8304
rect 15580 8276 15608 8316
rect 17037 8313 17049 8316
rect 17083 8313 17095 8347
rect 17512 8344 17540 8375
rect 17586 8372 17592 8424
rect 17644 8372 17650 8424
rect 18156 8412 18184 8452
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 19702 8480 19708 8492
rect 18524 8452 19708 8480
rect 18524 8424 18552 8452
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 18506 8412 18512 8424
rect 18156 8384 18512 8412
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 18690 8372 18696 8424
rect 18748 8372 18754 8424
rect 19978 8344 19984 8356
rect 17512 8316 19984 8344
rect 17037 8307 17095 8313
rect 17604 8288 17632 8316
rect 19978 8304 19984 8316
rect 20036 8304 20042 8356
rect 20272 8344 20300 8443
rect 20364 8412 20392 8520
rect 21269 8517 21281 8551
rect 21315 8548 21327 8551
rect 22830 8548 22836 8560
rect 21315 8520 22836 8548
rect 21315 8517 21327 8520
rect 21269 8511 21327 8517
rect 22830 8508 22836 8520
rect 22888 8508 22894 8560
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 23952 8489 23980 8588
rect 23937 8483 23995 8489
rect 22388 8452 23888 8480
rect 22388 8412 22416 8452
rect 20364 8384 22416 8412
rect 22462 8372 22468 8424
rect 22520 8412 22526 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 22520 8384 22569 8412
rect 22520 8372 22526 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 23860 8412 23888 8452
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24578 8412 24584 8424
rect 22557 8375 22615 8381
rect 22664 8384 22876 8412
rect 23860 8384 24584 8412
rect 22664 8344 22692 8384
rect 20272 8316 22692 8344
rect 22848 8344 22876 8384
rect 24578 8372 24584 8384
rect 24636 8372 24642 8424
rect 24762 8372 24768 8424
rect 24820 8372 24826 8424
rect 23842 8344 23848 8356
rect 22848 8316 23848 8344
rect 23842 8304 23848 8316
rect 23900 8304 23906 8356
rect 14016 8248 15608 8276
rect 17586 8236 17592 8288
rect 17644 8236 17650 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 11974 8072 11980 8084
rect 11103 8044 11980 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 13722 8072 13728 8084
rect 12768 8044 13728 8072
rect 12768 8032 12774 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14277 8075 14335 8081
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 14826 8072 14832 8084
rect 14323 8044 14832 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 19150 8072 19156 8084
rect 17920 8044 19156 8072
rect 17920 8032 17926 8044
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 20772 8044 22232 8072
rect 20772 8032 20778 8044
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 15194 8004 15200 8016
rect 8444 7976 13492 8004
rect 8444 7964 8450 7976
rect 11606 7896 11612 7948
rect 11664 7936 11670 7948
rect 11882 7936 11888 7948
rect 11664 7908 11888 7936
rect 11664 7896 11670 7908
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 13464 7945 13492 7976
rect 13556 7976 15200 8004
rect 13556 7945 13584 7976
rect 15194 7964 15200 7976
rect 15252 7964 15258 8016
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7905 13599 7939
rect 13541 7899 13599 7905
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 13780 7908 14841 7936
rect 13780 7896 13786 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15470 7936 15476 7948
rect 14976 7908 15476 7936
rect 14976 7896 14982 7908
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 15804 7908 16405 7936
rect 15804 7896 15810 7908
rect 16393 7905 16405 7908
rect 16439 7905 16451 7939
rect 21266 7936 21272 7948
rect 16393 7899 16451 7905
rect 17604 7908 21272 7936
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11698 7868 11704 7880
rect 11471 7840 11704 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12618 7868 12624 7880
rect 12492 7840 12624 7868
rect 12492 7828 12498 7840
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 16114 7868 16120 7880
rect 14691 7840 16120 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7868 16267 7871
rect 17604 7868 17632 7908
rect 21266 7896 21272 7908
rect 21324 7896 21330 7948
rect 21910 7896 21916 7948
rect 21968 7936 21974 7948
rect 22094 7936 22100 7948
rect 21968 7908 22100 7936
rect 21968 7896 21974 7908
rect 22094 7896 22100 7908
rect 22152 7896 22158 7948
rect 22204 7936 22232 8044
rect 23382 8032 23388 8084
rect 23440 8072 23446 8084
rect 24765 8075 24823 8081
rect 24765 8072 24777 8075
rect 23440 8044 24777 8072
rect 23440 8032 23446 8044
rect 24765 8041 24777 8044
rect 24811 8041 24823 8075
rect 24765 8035 24823 8041
rect 23934 7964 23940 8016
rect 23992 8004 23998 8016
rect 25317 8007 25375 8013
rect 25317 8004 25329 8007
rect 23992 7976 25329 8004
rect 23992 7964 23998 7976
rect 25317 7973 25329 7976
rect 25363 7973 25375 8007
rect 25317 7967 25375 7973
rect 25133 7939 25191 7945
rect 25133 7936 25145 7939
rect 22204 7908 25145 7936
rect 25133 7905 25145 7908
rect 25179 7905 25191 7939
rect 25133 7899 25191 7905
rect 16255 7840 17632 7868
rect 17681 7871 17739 7877
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 17681 7837 17693 7871
rect 17727 7868 17739 7871
rect 18598 7868 18604 7880
rect 17727 7840 18604 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 19518 7828 19524 7880
rect 19576 7828 19582 7880
rect 20438 7828 20444 7880
rect 20496 7828 20502 7880
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 24118 7868 24124 7880
rect 20680 7840 22094 7868
rect 23506 7840 24124 7868
rect 20680 7828 20686 7840
rect 12802 7760 12808 7812
rect 12860 7800 12866 7812
rect 14737 7803 14795 7809
rect 14737 7800 14749 7803
rect 12860 7772 14749 7800
rect 12860 7760 12866 7772
rect 14737 7769 14749 7772
rect 14783 7769 14795 7803
rect 17218 7800 17224 7812
rect 14737 7763 14795 7769
rect 14844 7772 17224 7800
rect 11517 7735 11575 7741
rect 11517 7701 11529 7735
rect 11563 7732 11575 7735
rect 11606 7732 11612 7744
rect 11563 7704 11612 7732
rect 11563 7701 11575 7704
rect 11517 7695 11575 7701
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12618 7732 12624 7744
rect 12391 7704 12624 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12952 7704 13001 7732
rect 12952 7692 12958 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 12989 7695 13047 7701
rect 14274 7692 14280 7744
rect 14332 7732 14338 7744
rect 14844 7732 14872 7772
rect 17218 7760 17224 7772
rect 17276 7760 17282 7812
rect 18693 7803 18751 7809
rect 18693 7769 18705 7803
rect 18739 7769 18751 7803
rect 18693 7763 18751 7769
rect 14332 7704 14872 7732
rect 15381 7735 15439 7741
rect 14332 7692 14338 7704
rect 15381 7701 15393 7735
rect 15427 7732 15439 7735
rect 15470 7732 15476 7744
rect 15427 7704 15476 7732
rect 15427 7701 15439 7704
rect 15381 7695 15439 7701
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15565 7735 15623 7741
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 15654 7732 15660 7744
rect 15611 7704 15660 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 16080 7704 16313 7732
rect 16080 7692 16086 7704
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 16850 7692 16856 7744
rect 16908 7692 16914 7744
rect 18708 7732 18736 7763
rect 19702 7760 19708 7812
rect 19760 7760 19766 7812
rect 21450 7760 21456 7812
rect 21508 7760 21514 7812
rect 22066 7800 22094 7840
rect 24118 7828 24124 7840
rect 24176 7828 24182 7880
rect 22066 7772 22324 7800
rect 21358 7732 21364 7744
rect 18708 7704 21364 7732
rect 21358 7692 21364 7704
rect 21416 7692 21422 7744
rect 22296 7732 22324 7772
rect 22370 7760 22376 7812
rect 22428 7760 22434 7812
rect 24673 7803 24731 7809
rect 24673 7800 24685 7803
rect 23676 7772 24685 7800
rect 23676 7732 23704 7772
rect 24673 7769 24685 7772
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 22296 7704 23704 7732
rect 23750 7692 23756 7744
rect 23808 7732 23814 7744
rect 23845 7735 23903 7741
rect 23845 7732 23857 7735
rect 23808 7704 23857 7732
rect 23808 7692 23814 7704
rect 23845 7701 23857 7704
rect 23891 7701 23903 7735
rect 23845 7695 23903 7701
rect 24118 7692 24124 7744
rect 24176 7692 24182 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 11149 7531 11207 7537
rect 9180 7500 10640 7528
rect 9180 7488 9186 7500
rect 9582 7460 9588 7472
rect 9048 7432 9588 7460
rect 9048 7401 9076 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 10612 7460 10640 7500
rect 11149 7497 11161 7531
rect 11195 7528 11207 7531
rect 11330 7528 11336 7540
rect 11195 7500 11336 7528
rect 11195 7497 11207 7500
rect 11149 7491 11207 7497
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11882 7488 11888 7540
rect 11940 7488 11946 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12342 7528 12348 7540
rect 12299 7500 12348 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12618 7488 12624 7540
rect 12676 7488 12682 7540
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 13688 7500 15485 7528
rect 13688 7488 13694 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 17218 7488 17224 7540
rect 17276 7488 17282 7540
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 17402 7528 17408 7540
rect 17359 7500 17408 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 17402 7488 17408 7500
rect 17460 7528 17466 7540
rect 17862 7528 17868 7540
rect 17460 7500 17868 7528
rect 17460 7488 17466 7500
rect 17862 7488 17868 7500
rect 17920 7528 17926 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 17920 7500 18061 7528
rect 17920 7488 17926 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 19610 7528 19616 7540
rect 18049 7491 18107 7497
rect 18524 7500 19616 7528
rect 14274 7460 14280 7472
rect 10612 7432 14280 7460
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 14734 7420 14740 7472
rect 14792 7420 14798 7472
rect 16117 7463 16175 7469
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 16574 7460 16580 7472
rect 16163 7432 16580 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 16574 7420 16580 7432
rect 16632 7460 16638 7472
rect 16850 7460 16856 7472
rect 16632 7432 16856 7460
rect 16632 7420 16638 7432
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 11330 7392 11336 7404
rect 10442 7364 11336 7392
rect 9033 7355 9091 7361
rect 11330 7352 11336 7364
rect 11388 7392 11394 7404
rect 11514 7392 11520 7404
rect 11388 7364 11520 7392
rect 11388 7352 11394 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 18524 7401 18552 7500
rect 19610 7488 19616 7500
rect 19668 7528 19674 7540
rect 20254 7528 20260 7540
rect 19668 7500 20260 7528
rect 19668 7488 19674 7500
rect 20254 7488 20260 7500
rect 20312 7528 20318 7540
rect 21910 7528 21916 7540
rect 20312 7500 21916 7528
rect 20312 7488 20318 7500
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 22922 7488 22928 7540
rect 22980 7528 22986 7540
rect 23382 7528 23388 7540
rect 22980 7500 23388 7528
rect 22980 7488 22986 7500
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 23293 7463 23351 7469
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24854 7460 24860 7472
rect 23339 7432 24860 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 20346 7392 20352 7404
rect 19944 7364 20352 7392
rect 19944 7352 19950 7364
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 20438 7352 20444 7404
rect 20496 7392 20502 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 20496 7364 21097 7392
rect 20496 7352 20502 7364
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 23474 7392 23480 7404
rect 22327 7364 23480 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 23474 7352 23480 7364
rect 23532 7352 23538 7404
rect 23934 7352 23940 7404
rect 23992 7352 23998 7404
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 10962 7324 10968 7336
rect 9355 7296 10968 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 11204 7296 12725 7324
rect 11204 7284 11210 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 16666 7324 16672 7336
rect 14047 7296 16672 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 12820 7256 12848 7287
rect 10796 7228 12848 7256
rect 10796 7200 10824 7228
rect 10778 7148 10784 7200
rect 10836 7148 10842 7200
rect 13740 7188 13768 7287
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7324 17555 7327
rect 17678 7324 17684 7336
rect 17543 7296 17684 7324
rect 17543 7293 17555 7296
rect 17497 7287 17555 7293
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 19242 7324 19248 7336
rect 18932 7296 19248 7324
rect 18932 7284 18938 7296
rect 19242 7284 19248 7296
rect 19300 7324 19306 7336
rect 20257 7327 20315 7333
rect 20257 7324 20269 7327
rect 19300 7296 20269 7324
rect 19300 7284 19306 7296
rect 20257 7293 20269 7296
rect 20303 7293 20315 7327
rect 20257 7287 20315 7293
rect 20714 7284 20720 7336
rect 20772 7324 20778 7336
rect 21177 7327 21235 7333
rect 21177 7324 21189 7327
rect 20772 7296 21189 7324
rect 20772 7284 20778 7296
rect 21177 7293 21189 7296
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7293 21327 7327
rect 21269 7287 21327 7293
rect 16301 7259 16359 7265
rect 16301 7225 16313 7259
rect 16347 7256 16359 7259
rect 16390 7256 16396 7268
rect 16347 7228 16396 7256
rect 16347 7225 16359 7228
rect 16301 7219 16359 7225
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 16482 7216 16488 7268
rect 16540 7256 16546 7268
rect 18414 7256 18420 7268
rect 16540 7228 18420 7256
rect 16540 7216 16546 7228
rect 18414 7216 18420 7228
rect 18472 7216 18478 7268
rect 19812 7228 20852 7256
rect 15102 7188 15108 7200
rect 13740 7160 15108 7188
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7188 16911 7191
rect 17770 7188 17776 7200
rect 16899 7160 17776 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 17957 7191 18015 7197
rect 17957 7157 17969 7191
rect 18003 7188 18015 7191
rect 18506 7188 18512 7200
rect 18003 7160 18512 7188
rect 18003 7157 18015 7160
rect 17957 7151 18015 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 18782 7197 18788 7200
rect 18772 7191 18788 7197
rect 18772 7157 18784 7191
rect 18840 7188 18846 7200
rect 19812 7188 19840 7228
rect 18840 7160 19840 7188
rect 18772 7151 18788 7157
rect 18782 7148 18788 7151
rect 18840 7148 18846 7160
rect 20714 7148 20720 7200
rect 20772 7148 20778 7200
rect 20824 7188 20852 7228
rect 21082 7216 21088 7268
rect 21140 7256 21146 7268
rect 21284 7256 21312 7287
rect 21358 7284 21364 7336
rect 21416 7324 21422 7336
rect 21416 7296 22094 7324
rect 21416 7284 21422 7296
rect 21140 7228 21312 7256
rect 22066 7256 22094 7296
rect 24762 7256 24768 7268
rect 22066 7228 24768 7256
rect 21140 7216 21146 7228
rect 24762 7216 24768 7228
rect 24820 7216 24826 7268
rect 21358 7188 21364 7200
rect 20824 7160 21364 7188
rect 21358 7148 21364 7160
rect 21416 7148 21422 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 11572 6956 12817 6984
rect 11572 6944 11578 6956
rect 12805 6953 12817 6956
rect 12851 6984 12863 6987
rect 13906 6984 13912 6996
rect 12851 6956 13912 6984
rect 12851 6953 12863 6956
rect 12805 6947 12863 6953
rect 13906 6944 13912 6956
rect 13964 6984 13970 6996
rect 14734 6984 14740 6996
rect 13964 6956 14740 6984
rect 13964 6944 13970 6956
rect 14734 6944 14740 6956
rect 14792 6984 14798 6996
rect 15654 6984 15660 6996
rect 14792 6956 15660 6984
rect 14792 6944 14798 6956
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16022 6944 16028 6996
rect 16080 6984 16086 6996
rect 20438 6984 20444 6996
rect 16080 6956 20444 6984
rect 16080 6944 16086 6956
rect 20438 6944 20444 6956
rect 20496 6944 20502 6996
rect 21450 6944 21456 6996
rect 21508 6984 21514 6996
rect 22554 6984 22560 6996
rect 21508 6956 22560 6984
rect 21508 6944 21514 6956
rect 22554 6944 22560 6956
rect 22612 6944 22618 6996
rect 12894 6876 12900 6928
rect 12952 6916 12958 6928
rect 16482 6916 16488 6928
rect 12952 6888 16488 6916
rect 12952 6876 12958 6888
rect 16482 6876 16488 6888
rect 16540 6876 16546 6928
rect 19518 6876 19524 6928
rect 19576 6916 19582 6928
rect 19886 6916 19892 6928
rect 19576 6888 19892 6916
rect 19576 6876 19582 6888
rect 19886 6876 19892 6888
rect 19944 6876 19950 6928
rect 21266 6876 21272 6928
rect 21324 6916 21330 6928
rect 22646 6916 22652 6928
rect 21324 6888 22652 6916
rect 21324 6876 21330 6888
rect 22646 6876 22652 6888
rect 22704 6876 22710 6928
rect 23658 6876 23664 6928
rect 23716 6916 23722 6928
rect 23716 6888 25176 6916
rect 23716 6876 23722 6888
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 11054 6848 11060 6860
rect 10827 6820 11060 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6848 12587 6851
rect 12710 6848 12716 6860
rect 12575 6820 12716 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 14366 6808 14372 6860
rect 14424 6848 14430 6860
rect 14424 6820 14872 6848
rect 14424 6808 14430 6820
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 14844 6789 14872 6820
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 19981 6851 20039 6857
rect 19981 6848 19993 6851
rect 16632 6820 19993 6848
rect 16632 6808 16638 6820
rect 19981 6817 19993 6820
rect 20027 6817 20039 6851
rect 19981 6811 20039 6817
rect 20346 6808 20352 6860
rect 20404 6848 20410 6860
rect 20441 6851 20499 6857
rect 20441 6848 20453 6851
rect 20404 6820 20453 6848
rect 20404 6808 20410 6820
rect 20441 6817 20453 6820
rect 20487 6817 20499 6851
rect 20441 6811 20499 6817
rect 22370 6808 22376 6860
rect 22428 6848 22434 6860
rect 25148 6857 25176 6888
rect 24397 6851 24455 6857
rect 24397 6848 24409 6851
rect 22428 6820 24409 6848
rect 22428 6808 22434 6820
rect 24397 6817 24409 6820
rect 24443 6848 24455 6851
rect 25133 6851 25191 6857
rect 24443 6820 24992 6848
rect 24443 6817 24455 6820
rect 24397 6811 24455 6817
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6780 15531 6783
rect 16298 6780 16304 6792
rect 15519 6752 16304 6780
rect 15519 6749 15531 6752
rect 15473 6743 15531 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 17000 6752 17141 6780
rect 17000 6740 17006 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 20364 6780 20392 6808
rect 18840 6752 20392 6780
rect 18840 6740 18846 6752
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 20898 6740 20904 6792
rect 20956 6780 20962 6792
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 20956 6752 22661 6780
rect 20956 6740 20962 6752
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 23934 6780 23940 6792
rect 22649 6743 22707 6749
rect 23768 6752 23940 6780
rect 11057 6715 11115 6721
rect 11057 6681 11069 6715
rect 11103 6712 11115 6715
rect 11330 6712 11336 6724
rect 11103 6684 11336 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 11514 6672 11520 6724
rect 11572 6672 11578 6724
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 12676 6684 14688 6712
rect 12676 6672 12682 6684
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 7558 6644 7564 6656
rect 4120 6616 7564 6644
rect 4120 6604 4126 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 13446 6604 13452 6656
rect 13504 6644 13510 6656
rect 14660 6653 14688 6684
rect 16482 6672 16488 6724
rect 16540 6672 16546 6724
rect 17405 6715 17463 6721
rect 17405 6681 17417 6715
rect 17451 6712 17463 6715
rect 17678 6712 17684 6724
rect 17451 6684 17684 6712
rect 17451 6681 17463 6684
rect 17405 6675 17463 6681
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 17862 6672 17868 6724
rect 17920 6672 17926 6724
rect 19889 6715 19947 6721
rect 19889 6712 19901 6715
rect 18708 6684 19901 6712
rect 13541 6647 13599 6653
rect 13541 6644 13553 6647
rect 13504 6616 13553 6644
rect 13504 6604 13510 6616
rect 13541 6613 13553 6616
rect 13587 6613 13599 6647
rect 13541 6607 13599 6613
rect 14645 6647 14703 6653
rect 14645 6613 14657 6647
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 18708 6644 18736 6684
rect 19889 6681 19901 6684
rect 19935 6681 19947 6715
rect 19889 6675 19947 6681
rect 22005 6715 22063 6721
rect 22005 6681 22017 6715
rect 22051 6712 22063 6715
rect 23768 6712 23796 6752
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 24964 6789 24992 6820
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 24949 6783 25007 6789
rect 24949 6749 24961 6783
rect 24995 6749 25007 6783
rect 24949 6743 25007 6749
rect 22051 6684 23796 6712
rect 23845 6715 23903 6721
rect 22051 6681 22063 6684
rect 22005 6675 22063 6681
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 24854 6712 24860 6724
rect 23891 6684 24860 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 24854 6672 24860 6684
rect 24912 6672 24918 6724
rect 14792 6616 18736 6644
rect 18877 6647 18935 6653
rect 14792 6604 14798 6616
rect 18877 6613 18889 6647
rect 18923 6644 18935 6647
rect 19334 6644 19340 6656
rect 18923 6616 19340 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19426 6604 19432 6656
rect 19484 6604 19490 6656
rect 19794 6604 19800 6656
rect 19852 6604 19858 6656
rect 21082 6604 21088 6656
rect 21140 6644 21146 6656
rect 23750 6644 23756 6656
rect 21140 6616 23756 6644
rect 21140 6604 21146 6616
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 24486 6604 24492 6656
rect 24544 6644 24550 6656
rect 24581 6647 24639 6653
rect 24581 6644 24593 6647
rect 24544 6616 24593 6644
rect 24544 6604 24550 6616
rect 24581 6613 24593 6616
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 24670 6604 24676 6656
rect 24728 6644 24734 6656
rect 25041 6647 25099 6653
rect 25041 6644 25053 6647
rect 24728 6616 25053 6644
rect 24728 6604 24734 6616
rect 25041 6613 25053 6616
rect 25087 6613 25099 6647
rect 25041 6607 25099 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 11146 6440 11152 6452
rect 10459 6412 11152 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6440 11759 6443
rect 12802 6440 12808 6452
rect 11747 6412 12808 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 17313 6443 17371 6449
rect 17313 6440 17325 6443
rect 13403 6412 17325 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 17313 6409 17325 6412
rect 17359 6409 17371 6443
rect 17313 6403 17371 6409
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 20254 6440 20260 6452
rect 19392 6412 20260 6440
rect 19392 6400 19398 6412
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 23658 6440 23664 6452
rect 22296 6412 23664 6440
rect 12161 6375 12219 6381
rect 12161 6341 12173 6375
rect 12207 6372 12219 6375
rect 12710 6372 12716 6384
rect 12207 6344 12716 6372
rect 12207 6341 12219 6344
rect 12161 6335 12219 6341
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 13630 6332 13636 6384
rect 13688 6372 13694 6384
rect 13688 6344 13952 6372
rect 13688 6332 13694 6344
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 6604 6276 10793 6304
rect 6604 6264 6610 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 11204 6276 12081 6304
rect 11204 6264 11210 6276
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 12069 6267 12127 6273
rect 13096 6276 13737 6304
rect 10870 6196 10876 6248
rect 10928 6196 10934 6248
rect 10962 6196 10968 6248
rect 11020 6196 11026 6248
rect 11330 6196 11336 6248
rect 11388 6236 11394 6248
rect 12253 6239 12311 6245
rect 12253 6236 12265 6239
rect 11388 6208 12265 6236
rect 11388 6196 11394 6208
rect 12253 6205 12265 6208
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 12986 6196 12992 6248
rect 13044 6196 13050 6248
rect 4246 6060 4252 6112
rect 4304 6100 4310 6112
rect 7834 6100 7840 6112
rect 4304 6072 7840 6100
rect 4304 6060 4310 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 13096 6100 13124 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 13924 6245 13952 6344
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 20898 6372 20904 6384
rect 14056 6344 18276 6372
rect 14056 6332 14062 6344
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15378 6304 15384 6316
rect 15151 6276 15384 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 16666 6264 16672 6316
rect 16724 6304 16730 6316
rect 16724 6276 17080 6304
rect 16724 6264 16730 6276
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 13504 6208 13829 6236
rect 13504 6196 13510 6208
rect 9732 6072 13124 6100
rect 13648 6100 13676 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 16114 6196 16120 6248
rect 16172 6196 16178 6248
rect 16298 6196 16304 6248
rect 16356 6236 16362 6248
rect 17052 6236 17080 6276
rect 17218 6264 17224 6316
rect 17276 6264 17282 6316
rect 17954 6304 17960 6316
rect 17328 6276 17960 6304
rect 17328 6236 17356 6276
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 18248 6313 18276 6344
rect 18340 6344 20904 6372
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 16356 6208 16988 6236
rect 17052 6208 17356 6236
rect 16356 6196 16362 6208
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 16853 6171 16911 6177
rect 16853 6168 16865 6171
rect 13780 6140 16865 6168
rect 13780 6128 13786 6140
rect 16853 6137 16865 6140
rect 16899 6137 16911 6171
rect 16960 6168 16988 6208
rect 17402 6196 17408 6248
rect 17460 6196 17466 6248
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18340 6236 18368 6344
rect 20898 6332 20904 6344
rect 20956 6332 20962 6384
rect 21266 6332 21272 6384
rect 21324 6372 21330 6384
rect 21726 6372 21732 6384
rect 21324 6344 21732 6372
rect 21324 6332 21330 6344
rect 21726 6332 21732 6344
rect 21784 6332 21790 6384
rect 22296 6381 22324 6412
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 23750 6400 23756 6452
rect 23808 6400 23814 6452
rect 22281 6375 22339 6381
rect 22281 6341 22293 6375
rect 22327 6341 22339 6375
rect 24118 6372 24124 6384
rect 23506 6344 24124 6372
rect 22281 6335 22339 6341
rect 24118 6332 24124 6344
rect 24176 6332 24182 6384
rect 24302 6332 24308 6384
rect 24360 6332 24366 6384
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 20346 6304 20352 6316
rect 20303 6276 20352 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 20346 6264 20352 6276
rect 20404 6264 20410 6316
rect 21910 6264 21916 6316
rect 21968 6304 21974 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21968 6276 22017 6304
rect 21968 6264 21974 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 24670 6264 24676 6316
rect 24728 6304 24734 6316
rect 25041 6307 25099 6313
rect 25041 6304 25053 6307
rect 24728 6276 25053 6304
rect 24728 6264 24734 6276
rect 25041 6273 25053 6276
rect 25087 6273 25099 6307
rect 25041 6267 25099 6273
rect 17920 6208 18368 6236
rect 19429 6239 19487 6245
rect 17920 6196 17926 6208
rect 19429 6205 19441 6239
rect 19475 6236 19487 6239
rect 20622 6236 20628 6248
rect 19475 6208 20628 6236
rect 19475 6205 19487 6208
rect 19429 6199 19487 6205
rect 20622 6196 20628 6208
rect 20680 6196 20686 6248
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21726 6236 21732 6248
rect 21315 6208 21732 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21726 6196 21732 6208
rect 21784 6196 21790 6248
rect 23014 6196 23020 6248
rect 23072 6236 23078 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 23072 6208 25237 6236
rect 23072 6196 23078 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 24489 6171 24547 6177
rect 24489 6168 24501 6171
rect 16960 6140 22094 6168
rect 16853 6131 16911 6137
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 13648 6072 14381 6100
rect 9732 6060 9738 6072
rect 14369 6069 14381 6072
rect 14415 6069 14427 6103
rect 14369 6063 14427 6069
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 21450 6100 21456 6112
rect 16540 6072 21456 6100
rect 16540 6060 16546 6072
rect 21450 6060 21456 6072
rect 21508 6060 21514 6112
rect 22066 6100 22094 6140
rect 23308 6140 24501 6168
rect 23308 6100 23336 6140
rect 24489 6137 24501 6140
rect 24535 6137 24547 6171
rect 24489 6131 24547 6137
rect 22066 6072 23336 6100
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 11793 5899 11851 5905
rect 11793 5896 11805 5899
rect 11388 5868 11805 5896
rect 11388 5856 11394 5868
rect 11793 5865 11805 5868
rect 11839 5865 11851 5899
rect 11793 5859 11851 5865
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13998 5896 14004 5908
rect 13587 5868 14004 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14182 5856 14188 5908
rect 14240 5856 14246 5908
rect 14734 5856 14740 5908
rect 14792 5856 14798 5908
rect 15304 5868 17264 5896
rect 12897 5831 12955 5837
rect 12897 5797 12909 5831
rect 12943 5828 12955 5831
rect 13722 5828 13728 5840
rect 12943 5800 13728 5828
rect 12943 5797 12955 5800
rect 12897 5791 12955 5797
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10778 5760 10784 5772
rect 10367 5732 10784 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11514 5760 11520 5772
rect 11440 5732 11520 5760
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9640 5664 10057 5692
rect 9640 5652 9646 5664
rect 10045 5661 10057 5664
rect 10091 5661 10103 5695
rect 11440 5678 11468 5732
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 12253 5763 12311 5769
rect 12253 5729 12265 5763
rect 12299 5760 12311 5763
rect 15304 5760 15332 5868
rect 17236 5828 17264 5868
rect 17678 5856 17684 5908
rect 17736 5856 17742 5908
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 17828 5868 20208 5896
rect 17828 5856 17834 5868
rect 19794 5828 19800 5840
rect 17236 5800 19800 5828
rect 19794 5788 19800 5800
rect 19852 5788 19858 5840
rect 12299 5732 15332 5760
rect 12299 5729 12311 5732
rect 12253 5723 12311 5729
rect 15378 5720 15384 5772
rect 15436 5720 15442 5772
rect 16942 5760 16948 5772
rect 15948 5732 16948 5760
rect 13081 5695 13139 5701
rect 10045 5655 10103 5661
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13538 5692 13544 5704
rect 13127 5664 13544 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 13740 5624 13768 5655
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15948 5701 15976 5732
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 18380 5732 18613 5760
rect 18380 5720 18386 5732
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18785 5763 18843 5769
rect 18785 5729 18797 5763
rect 18831 5760 18843 5763
rect 18874 5760 18880 5772
rect 18831 5732 18880 5760
rect 18831 5729 18843 5732
rect 18785 5723 18843 5729
rect 18874 5720 18880 5732
rect 18932 5720 18938 5772
rect 19150 5720 19156 5772
rect 19208 5760 19214 5772
rect 19889 5763 19947 5769
rect 19889 5760 19901 5763
rect 19208 5732 19901 5760
rect 19208 5720 19214 5732
rect 19889 5729 19901 5732
rect 19935 5729 19947 5763
rect 20180 5760 20208 5868
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20312 5868 23704 5896
rect 20312 5856 20318 5868
rect 20438 5788 20444 5840
rect 20496 5828 20502 5840
rect 20496 5800 22232 5828
rect 20496 5788 20502 5800
rect 22204 5769 22232 5800
rect 23676 5769 23704 5868
rect 24118 5856 24124 5908
rect 24176 5856 24182 5908
rect 24302 5856 24308 5908
rect 24360 5896 24366 5908
rect 25133 5899 25191 5905
rect 25133 5896 25145 5899
rect 24360 5868 25145 5896
rect 24360 5856 24366 5868
rect 25133 5865 25145 5868
rect 25179 5865 25191 5899
rect 25133 5859 25191 5865
rect 24857 5831 24915 5837
rect 24857 5797 24869 5831
rect 24903 5828 24915 5831
rect 24946 5828 24952 5840
rect 24903 5800 24952 5828
rect 24903 5797 24915 5800
rect 24857 5791 24915 5797
rect 24946 5788 24952 5800
rect 25004 5788 25010 5840
rect 22189 5763 22247 5769
rect 20180 5732 21404 5760
rect 19889 5723 19947 5729
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15160 5664 15945 5692
rect 15160 5652 15166 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 20990 5692 20996 5704
rect 19659 5664 20996 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 20990 5652 20996 5664
rect 21048 5652 21054 5704
rect 21266 5652 21272 5704
rect 21324 5652 21330 5704
rect 21376 5692 21404 5732
rect 22189 5729 22201 5763
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 23661 5763 23719 5769
rect 23661 5729 23673 5763
rect 23707 5729 23719 5763
rect 23661 5723 23719 5729
rect 23569 5695 23627 5701
rect 23569 5692 23581 5695
rect 21376 5664 23581 5692
rect 23569 5661 23581 5664
rect 23615 5661 23627 5695
rect 23569 5655 23627 5661
rect 24578 5652 24584 5704
rect 24636 5692 24642 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 24636 5664 24685 5692
rect 24636 5652 24642 5664
rect 24673 5661 24685 5664
rect 24719 5692 24731 5695
rect 25317 5695 25375 5701
rect 25317 5692 25329 5695
rect 24719 5664 25329 5692
rect 24719 5661 24731 5664
rect 24673 5655 24731 5661
rect 25317 5661 25329 5664
rect 25363 5661 25375 5695
rect 25317 5655 25375 5661
rect 11624 5596 13768 5624
rect 14461 5627 14519 5633
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 11624 5556 11652 5596
rect 14461 5593 14473 5627
rect 14507 5624 14519 5627
rect 15194 5624 15200 5636
rect 14507 5596 15200 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 15194 5584 15200 5596
rect 15252 5584 15258 5636
rect 16209 5627 16267 5633
rect 16209 5593 16221 5627
rect 16255 5624 16267 5627
rect 16482 5624 16488 5636
rect 16255 5596 16488 5624
rect 16255 5593 16267 5596
rect 16209 5587 16267 5593
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 16666 5584 16672 5636
rect 16724 5584 16730 5636
rect 18509 5627 18567 5633
rect 18509 5593 18521 5627
rect 18555 5624 18567 5627
rect 19242 5624 19248 5636
rect 18555 5596 19248 5624
rect 18555 5593 18567 5596
rect 18509 5587 18567 5593
rect 19242 5584 19248 5596
rect 19300 5584 19306 5636
rect 20622 5584 20628 5636
rect 20680 5624 20686 5636
rect 23382 5624 23388 5636
rect 20680 5596 23388 5624
rect 20680 5584 20686 5596
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 23474 5584 23480 5636
rect 23532 5584 23538 5636
rect 10468 5528 11652 5556
rect 10468 5516 10474 5528
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 15105 5559 15163 5565
rect 15105 5556 15117 5559
rect 12492 5528 15117 5556
rect 12492 5516 12498 5528
rect 15105 5525 15117 5528
rect 15151 5525 15163 5559
rect 15105 5519 15163 5525
rect 18141 5559 18199 5565
rect 18141 5525 18153 5559
rect 18187 5556 18199 5559
rect 18322 5556 18328 5568
rect 18187 5528 18328 5556
rect 18187 5525 18199 5528
rect 18141 5519 18199 5525
rect 18322 5516 18328 5528
rect 18380 5516 18386 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 21910 5556 21916 5568
rect 19392 5528 21916 5556
rect 19392 5516 19398 5528
rect 21910 5516 21916 5528
rect 21968 5516 21974 5568
rect 23106 5516 23112 5568
rect 23164 5516 23170 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 11514 5312 11520 5364
rect 11572 5312 11578 5364
rect 12526 5312 12532 5364
rect 12584 5312 12590 5364
rect 13630 5312 13636 5364
rect 13688 5312 13694 5364
rect 14274 5312 14280 5364
rect 14332 5352 14338 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14332 5324 14933 5352
rect 14332 5312 14338 5324
rect 14921 5321 14933 5324
rect 14967 5352 14979 5355
rect 17402 5352 17408 5364
rect 14967 5324 17408 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 18932 5324 20208 5352
rect 18932 5312 18938 5324
rect 13354 5284 13360 5296
rect 10612 5256 13360 5284
rect 10612 5225 10640 5256
rect 13354 5244 13360 5256
rect 13412 5244 13418 5296
rect 13449 5287 13507 5293
rect 13449 5253 13461 5287
rect 13495 5284 13507 5287
rect 13648 5284 13676 5312
rect 13495 5256 13676 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 13906 5244 13912 5296
rect 13964 5244 13970 5296
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 19426 5284 19432 5296
rect 14792 5256 19432 5284
rect 14792 5244 14798 5256
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 20180 5284 20208 5324
rect 21358 5312 21364 5364
rect 21416 5312 21422 5364
rect 21542 5312 21548 5364
rect 21600 5352 21606 5364
rect 21910 5352 21916 5364
rect 21600 5324 21916 5352
rect 21600 5312 21606 5324
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 20180 5256 20378 5284
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 12713 5219 12771 5225
rect 11112 5188 12434 5216
rect 11112 5176 11118 5188
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 11422 5148 11428 5160
rect 10367 5120 11428 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5148 11851 5151
rect 12066 5148 12072 5160
rect 11839 5120 12072 5148
rect 11839 5117 11851 5120
rect 11793 5111 11851 5117
rect 12066 5108 12072 5120
rect 12124 5108 12130 5160
rect 12406 5148 12434 5188
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 13078 5216 13084 5228
rect 12759 5188 13084 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 15838 5176 15844 5228
rect 15896 5216 15902 5228
rect 16666 5216 16672 5228
rect 15896 5188 16672 5216
rect 15896 5176 15902 5188
rect 16666 5176 16672 5188
rect 16724 5216 16730 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 16724 5188 16865 5216
rect 16724 5176 16730 5188
rect 16853 5185 16865 5188
rect 16899 5216 16911 5219
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16899 5188 17049 5216
rect 16899 5185 16911 5188
rect 16853 5179 16911 5185
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 13173 5151 13231 5157
rect 13173 5148 13185 5151
rect 12406 5120 13185 5148
rect 13173 5117 13185 5120
rect 13219 5117 13231 5151
rect 13173 5111 13231 5117
rect 6086 4972 6092 5024
rect 6144 4972 6150 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6512 4984 7205 5012
rect 6512 4972 6518 4984
rect 7193 4981 7205 4984
rect 7239 5012 7251 5015
rect 11514 5012 11520 5024
rect 7239 4984 11520 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 13188 5012 13216 5111
rect 13998 5108 14004 5160
rect 14056 5148 14062 5160
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 14056 5120 15485 5148
rect 14056 5108 14062 5120
rect 15473 5117 15485 5120
rect 15519 5117 15531 5151
rect 15473 5111 15531 5117
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15712 5120 15761 5148
rect 15712 5108 15718 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 17422 5148 17450 5179
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 17828 5188 19564 5216
rect 17828 5176 17834 5188
rect 17422 5120 19472 5148
rect 15749 5111 15807 5117
rect 19334 5080 19340 5092
rect 14476 5052 19340 5080
rect 13906 5012 13912 5024
rect 13188 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14476 5012 14504 5052
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 14240 4984 14504 5012
rect 14240 4972 14246 4984
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 18693 5015 18751 5021
rect 18693 5012 18705 5015
rect 16724 4984 18705 5012
rect 16724 4972 16730 4984
rect 18693 4981 18705 4984
rect 18739 5012 18751 5015
rect 18874 5012 18880 5024
rect 18739 4984 18880 5012
rect 18739 4981 18751 4984
rect 18693 4975 18751 4981
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 19444 5012 19472 5120
rect 19536 5080 19564 5188
rect 19610 5176 19616 5228
rect 19668 5176 19674 5228
rect 22186 5176 22192 5228
rect 22244 5176 22250 5228
rect 24029 5219 24087 5225
rect 22848 5188 23060 5216
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5148 19947 5151
rect 21266 5148 21272 5160
rect 19935 5120 21272 5148
rect 19935 5117 19947 5120
rect 19889 5111 19947 5117
rect 21266 5108 21272 5120
rect 21324 5108 21330 5160
rect 21358 5108 21364 5160
rect 21416 5148 21422 5160
rect 22848 5148 22876 5188
rect 21416 5120 22876 5148
rect 22925 5151 22983 5157
rect 21416 5108 21422 5120
rect 22925 5117 22937 5151
rect 22971 5117 22983 5151
rect 23032 5148 23060 5188
rect 24029 5185 24041 5219
rect 24075 5216 24087 5219
rect 25038 5216 25044 5228
rect 24075 5188 25044 5216
rect 24075 5185 24087 5188
rect 24029 5179 24087 5185
rect 25038 5176 25044 5188
rect 25096 5176 25102 5228
rect 24305 5151 24363 5157
rect 24305 5148 24317 5151
rect 23032 5120 24317 5148
rect 22925 5111 22983 5117
rect 24305 5117 24317 5120
rect 24351 5117 24363 5151
rect 24305 5111 24363 5117
rect 19610 5080 19616 5092
rect 19536 5052 19616 5080
rect 19610 5040 19616 5052
rect 19668 5040 19674 5092
rect 20898 5040 20904 5092
rect 20956 5080 20962 5092
rect 22940 5080 22968 5111
rect 20956 5052 22968 5080
rect 20956 5040 20962 5052
rect 22094 5012 22100 5024
rect 19444 4984 22100 5012
rect 22094 4972 22100 4984
rect 22152 4972 22158 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 12066 4768 12072 4820
rect 12124 4808 12130 4820
rect 14182 4808 14188 4820
rect 12124 4780 14188 4808
rect 12124 4768 12130 4780
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 17218 4808 17224 4820
rect 15028 4780 17224 4808
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4709 1639 4743
rect 12802 4740 12808 4752
rect 1581 4703 1639 4709
rect 9692 4712 12808 4740
rect 1596 4672 1624 4703
rect 5077 4675 5135 4681
rect 1596 4644 2820 4672
rect 1762 4564 1768 4616
rect 1820 4564 1826 4616
rect 2792 4613 2820 4644
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 9582 4672 9588 4684
rect 5123 4644 9588 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 9692 4681 9720 4712
rect 12802 4700 12808 4712
rect 12860 4700 12866 4752
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9950 4632 9956 4684
rect 10008 4632 10014 4684
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 13998 4672 14004 4684
rect 11296 4644 14004 4672
rect 11296 4632 11302 4644
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 15028 4672 15056 4780
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 18969 4811 19027 4817
rect 18969 4808 18981 4811
rect 18932 4780 18981 4808
rect 18932 4768 18938 4780
rect 18969 4777 18981 4780
rect 19015 4808 19027 4811
rect 19015 4780 19334 4808
rect 19015 4777 19027 4780
rect 18969 4771 19027 4777
rect 16574 4700 16580 4752
rect 16632 4740 16638 4752
rect 16853 4743 16911 4749
rect 16853 4740 16865 4743
rect 16632 4712 16865 4740
rect 16632 4700 16638 4712
rect 16853 4709 16865 4712
rect 16899 4709 16911 4743
rect 19306 4740 19334 4780
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 19852 4780 20852 4808
rect 19852 4768 19858 4780
rect 20824 4740 20852 4780
rect 21266 4768 21272 4820
rect 21324 4768 21330 4820
rect 24394 4768 24400 4820
rect 24452 4808 24458 4820
rect 24765 4811 24823 4817
rect 24765 4808 24777 4811
rect 24452 4780 24777 4808
rect 24452 4768 24458 4780
rect 24765 4777 24777 4780
rect 24811 4777 24823 4811
rect 24765 4771 24823 4777
rect 19306 4712 19656 4740
rect 20824 4712 22094 4740
rect 16853 4703 16911 4709
rect 14507 4644 15056 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 15102 4632 15108 4684
rect 15160 4632 15166 4684
rect 15378 4632 15384 4684
rect 15436 4632 15442 4684
rect 19518 4632 19524 4684
rect 19576 4632 19582 4684
rect 19628 4672 19656 4712
rect 22066 4672 22094 4712
rect 22189 4675 22247 4681
rect 22189 4672 22201 4675
rect 19628 4644 21036 4672
rect 22066 4644 22201 4672
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3467 4576 3985 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 6454 4564 6460 4616
rect 6512 4564 6518 4616
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 6696 4576 7849 4604
rect 6696 4564 6702 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 11054 4564 11060 4616
rect 11112 4564 11118 4616
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4604 11391 4607
rect 12529 4607 12587 4613
rect 11379 4576 12434 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 4617 4539 4675 4545
rect 4617 4505 4629 4539
rect 4663 4536 4675 4539
rect 5353 4539 5411 4545
rect 5353 4536 5365 4539
rect 4663 4508 5365 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 5353 4505 5365 4508
rect 5399 4505 5411 4539
rect 5353 4499 5411 4505
rect 7098 4496 7104 4548
rect 7156 4496 7162 4548
rect 12406 4536 12434 4576
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12618 4604 12624 4616
rect 12575 4576 12624 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 14182 4564 14188 4616
rect 14240 4604 14246 4616
rect 14918 4604 14924 4616
rect 14240 4576 14924 4604
rect 14240 4564 14246 4576
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 17494 4564 17500 4616
rect 17552 4564 17558 4616
rect 13170 4536 13176 4548
rect 12406 4508 13176 4536
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 13262 4496 13268 4548
rect 13320 4496 13326 4548
rect 15654 4536 15660 4548
rect 13372 4508 15660 4536
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 7432 4440 7481 4468
rect 7432 4428 7438 4440
rect 7469 4437 7481 4440
rect 7515 4437 7527 4471
rect 7469 4431 7527 4437
rect 7742 4428 7748 4480
rect 7800 4428 7806 4480
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7892 4440 8033 4468
rect 7892 4428 7898 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 8294 4428 8300 4480
rect 8352 4428 8358 4480
rect 8570 4428 8576 4480
rect 8628 4428 8634 4480
rect 8754 4428 8760 4480
rect 8812 4428 8818 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 13372 4468 13400 4508
rect 15654 4496 15660 4508
rect 15712 4496 15718 4548
rect 15838 4496 15844 4548
rect 15896 4496 15902 4548
rect 18509 4539 18567 4545
rect 18509 4505 18521 4539
rect 18555 4536 18567 4539
rect 19518 4536 19524 4548
rect 18555 4508 19524 4536
rect 18555 4505 18567 4508
rect 18509 4499 18567 4505
rect 19518 4496 19524 4508
rect 19576 4496 19582 4548
rect 19797 4539 19855 4545
rect 19797 4505 19809 4539
rect 19843 4505 19855 4539
rect 21008 4536 21036 4644
rect 22189 4641 22201 4644
rect 22235 4641 22247 4675
rect 22189 4635 22247 4641
rect 21913 4607 21971 4613
rect 21913 4573 21925 4607
rect 21959 4604 21971 4607
rect 22002 4604 22008 4616
rect 21959 4576 22008 4604
rect 21959 4573 21971 4576
rect 21913 4567 21971 4573
rect 22002 4564 22008 4576
rect 22060 4564 22066 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 23584 4576 24685 4604
rect 21542 4536 21548 4548
rect 21008 4522 21548 4536
rect 21022 4508 21548 4522
rect 19797 4499 19855 4505
rect 12492 4440 13400 4468
rect 12492 4428 12498 4440
rect 13446 4428 13452 4480
rect 13504 4468 13510 4480
rect 17862 4468 17868 4480
rect 13504 4440 17868 4468
rect 13504 4428 13510 4440
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 19812 4468 19840 4499
rect 21542 4496 21548 4508
rect 21600 4496 21606 4548
rect 23584 4536 23612 4576
rect 24673 4573 24685 4576
rect 24719 4604 24731 4607
rect 25133 4607 25191 4613
rect 25133 4604 25145 4607
rect 24719 4576 25145 4604
rect 24719 4573 24731 4576
rect 24673 4567 24731 4573
rect 25133 4573 25145 4576
rect 25179 4573 25191 4607
rect 25133 4567 25191 4573
rect 22066 4508 23612 4536
rect 21082 4468 21088 4480
rect 19812 4440 21088 4468
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 21910 4428 21916 4480
rect 21968 4468 21974 4480
rect 22066 4468 22094 4508
rect 23658 4496 23664 4548
rect 23716 4536 23722 4548
rect 24121 4539 24179 4545
rect 24121 4536 24133 4539
rect 23716 4508 24133 4536
rect 23716 4496 23722 4508
rect 24121 4505 24133 4508
rect 24167 4505 24179 4539
rect 24121 4499 24179 4505
rect 24302 4496 24308 4548
rect 24360 4536 24366 4548
rect 25317 4539 25375 4545
rect 25317 4536 25329 4539
rect 24360 4508 25329 4536
rect 24360 4496 24366 4508
rect 25317 4505 25329 4508
rect 25363 4505 25375 4539
rect 25317 4499 25375 4505
rect 21968 4440 22094 4468
rect 21968 4428 21974 4440
rect 23750 4428 23756 4480
rect 23808 4428 23814 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 7190 4224 7196 4276
rect 7248 4224 7254 4276
rect 10042 4273 10048 4276
rect 9999 4267 10048 4273
rect 9999 4233 10011 4267
rect 10045 4233 10048 4267
rect 9999 4227 10048 4233
rect 10042 4224 10048 4227
rect 10100 4224 10106 4276
rect 11330 4264 11336 4276
rect 11256 4236 11336 4264
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1544 4100 1593 4128
rect 1544 4088 1550 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 2915 4100 3280 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 2774 4060 2780 4072
rect 2746 4020 2780 4060
rect 2832 4020 2838 4072
rect 3252 4069 3280 4100
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4120 4100 4353 4128
rect 4120 4088 4126 4100
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 5031 4100 5365 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5353 4097 5365 4100
rect 5399 4128 5411 4131
rect 5902 4128 5908 4140
rect 5399 4100 5908 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 5994 4088 6000 4140
rect 6052 4088 6058 4140
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 7006 4128 7012 4140
rect 6779 4100 7012 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7374 4088 7380 4140
rect 7432 4088 7438 4140
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 7616 4100 8033 4128
rect 7616 4088 7622 4100
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8352 4100 8677 4128
rect 8352 4088 8358 4100
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9272 4100 9321 4128
rect 9272 4088 9278 4100
rect 9309 4097 9321 4100
rect 9355 4128 9367 4131
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 9355 4100 11069 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 3694 4060 3700 4072
rect 3283 4032 3700 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 9674 4060 9680 4072
rect 7852 4032 9680 4060
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 2746 3992 2774 4020
rect 3329 3995 3387 4001
rect 3329 3992 3341 3995
rect 2271 3964 2774 3992
rect 2884 3964 3341 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2556 3896 2697 3924
rect 2556 3884 2562 3896
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 2685 3887 2743 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2884 3924 2912 3964
rect 3329 3961 3341 3964
rect 3375 3961 3387 3995
rect 3329 3955 3387 3961
rect 4154 3952 4160 4004
rect 4212 3952 4218 4004
rect 4816 3964 6500 3992
rect 2832 3896 2912 3924
rect 2832 3884 2838 3896
rect 3510 3884 3516 3936
rect 3568 3884 3574 3936
rect 3881 3927 3939 3933
rect 3881 3893 3893 3927
rect 3927 3924 3939 3927
rect 4062 3924 4068 3936
rect 3927 3896 4068 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4816 3933 4844 3964
rect 4801 3927 4859 3933
rect 4801 3893 4813 3927
rect 4847 3893 4859 3927
rect 4801 3887 4859 3893
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 5810 3884 5816 3936
rect 5868 3884 5874 3936
rect 6472 3924 6500 3964
rect 6546 3952 6552 4004
rect 6604 3952 6610 4004
rect 7852 4001 7880 4032
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4060 9827 4063
rect 9950 4060 9956 4072
rect 9815 4032 9956 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 11256 4060 11284 4236
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 13320 4236 15516 4264
rect 13320 4224 13326 4236
rect 13170 4156 13176 4208
rect 13228 4196 13234 4208
rect 13814 4196 13820 4208
rect 13228 4168 13820 4196
rect 13228 4156 13234 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 14185 4199 14243 4205
rect 14185 4165 14197 4199
rect 14231 4196 14243 4199
rect 14274 4196 14280 4208
rect 14231 4168 14280 4196
rect 14231 4165 14243 4168
rect 14185 4159 14243 4165
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 15488 4196 15516 4236
rect 21542 4224 21548 4276
rect 21600 4224 21606 4276
rect 21634 4224 21640 4276
rect 21692 4264 21698 4276
rect 22002 4264 22008 4276
rect 21692 4236 22008 4264
rect 21692 4224 21698 4236
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 22094 4224 22100 4276
rect 22152 4224 22158 4276
rect 22738 4224 22744 4276
rect 22796 4224 22802 4276
rect 15488 4168 17908 4196
rect 11333 4131 11391 4137
rect 11333 4097 11345 4131
rect 11379 4128 11391 4131
rect 11422 4128 11428 4140
rect 11379 4100 11428 4128
rect 11379 4097 11391 4100
rect 11333 4091 11391 4097
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 15838 4128 15844 4140
rect 15318 4100 15844 4128
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16390 4128 16396 4140
rect 16347 4100 16396 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17586 4128 17592 4140
rect 17083 4100 17592 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 17880 4128 17908 4168
rect 20162 4156 20168 4208
rect 20220 4196 20226 4208
rect 21910 4196 21916 4208
rect 20220 4168 21916 4196
rect 20220 4156 20226 4168
rect 21910 4156 21916 4168
rect 21968 4156 21974 4208
rect 23290 4156 23296 4208
rect 23348 4196 23354 4208
rect 23348 4168 24256 4196
rect 23348 4156 23354 4168
rect 18506 4128 18512 4140
rect 17880 4100 18512 4128
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4128 18935 4131
rect 19058 4128 19064 4140
rect 18923 4100 19064 4128
rect 18923 4097 18935 4100
rect 18877 4091 18935 4097
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 20898 4088 20904 4140
rect 20956 4088 20962 4140
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 23474 4128 23480 4140
rect 22327 4100 23480 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 23569 4131 23627 4137
rect 23569 4097 23581 4131
rect 23615 4128 23627 4131
rect 24026 4128 24032 4140
rect 23615 4100 24032 4128
rect 23615 4097 23627 4100
rect 23569 4091 23627 4097
rect 24026 4088 24032 4100
rect 24084 4088 24090 4140
rect 24228 4137 24256 4168
rect 24213 4131 24271 4137
rect 24213 4097 24225 4131
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 24302 4088 24308 4140
rect 24360 4128 24366 4140
rect 24673 4131 24731 4137
rect 24673 4128 24685 4131
rect 24360 4100 24685 4128
rect 24360 4088 24366 4100
rect 24673 4097 24685 4100
rect 24719 4097 24731 4131
rect 24673 4091 24731 4097
rect 12526 4060 12532 4072
rect 10100 4032 11284 4060
rect 12406 4032 12532 4060
rect 10100 4020 10106 4032
rect 7837 3995 7895 4001
rect 7837 3961 7849 3995
rect 7883 3961 7895 3995
rect 7837 3955 7895 3961
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 8846 3992 8852 4004
rect 8527 3964 8852 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 9125 3995 9183 4001
rect 9125 3961 9137 3995
rect 9171 3992 9183 3995
rect 12406 3992 12434 4032
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13311 4032 16160 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 9171 3964 12434 3992
rect 9171 3961 9183 3964
rect 9125 3955 9183 3961
rect 15378 3952 15384 4004
rect 15436 3992 15442 4004
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 15436 3964 15669 3992
rect 15436 3952 15442 3964
rect 15657 3961 15669 3964
rect 15703 3961 15715 3995
rect 16132 3992 16160 4032
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16264 4032 17325 4060
rect 16264 4020 16270 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17402 4020 17408 4072
rect 17460 4060 17466 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 17460 4032 19165 4060
rect 17460 4020 17466 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 20993 4063 21051 4069
rect 20993 4060 21005 4063
rect 20772 4032 21005 4060
rect 20772 4020 20778 4032
rect 20993 4029 21005 4032
rect 21039 4029 21051 4063
rect 20993 4023 21051 4029
rect 21177 4063 21235 4069
rect 21177 4029 21189 4063
rect 21223 4060 21235 4063
rect 21266 4060 21272 4072
rect 21223 4032 21272 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 17770 3992 17776 4004
rect 16132 3964 17776 3992
rect 15657 3955 15715 3961
rect 17770 3952 17776 3964
rect 17828 3952 17834 4004
rect 18690 3952 18696 4004
rect 18748 3992 18754 4004
rect 20254 3992 20260 4004
rect 18748 3964 20260 3992
rect 18748 3952 18754 3964
rect 20254 3952 20260 3964
rect 20312 3952 20318 4004
rect 20346 3952 20352 4004
rect 20404 3992 20410 4004
rect 23385 3995 23443 4001
rect 23385 3992 23397 3995
rect 20404 3964 23397 3992
rect 20404 3952 20410 3964
rect 23385 3961 23397 3964
rect 23431 3961 23443 3995
rect 23385 3955 23443 3961
rect 10042 3924 10048 3936
rect 6472 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10686 3924 10692 3936
rect 10192 3896 10692 3924
rect 10192 3884 10198 3896
rect 10686 3884 10692 3896
rect 10744 3924 10750 3936
rect 10873 3927 10931 3933
rect 10873 3924 10885 3927
rect 10744 3896 10885 3924
rect 10744 3884 10750 3896
rect 10873 3893 10885 3896
rect 10919 3893 10931 3927
rect 10873 3887 10931 3893
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 11698 3924 11704 3936
rect 11655 3896 11704 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 12526 3924 12532 3936
rect 11839 3896 12532 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 19058 3924 19064 3936
rect 16163 3896 19064 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 20530 3884 20536 3936
rect 20588 3884 20594 3936
rect 24026 3884 24032 3936
rect 24084 3884 24090 3936
rect 24578 3884 24584 3936
rect 24636 3924 24642 3936
rect 25317 3927 25375 3933
rect 25317 3924 25329 3927
rect 24636 3896 25329 3924
rect 24636 3884 24642 3896
rect 25317 3893 25329 3896
rect 25363 3893 25375 3927
rect 25317 3887 25375 3893
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 2593 3723 2651 3729
rect 2593 3720 2605 3723
rect 1820 3692 2605 3720
rect 1820 3680 1826 3692
rect 2593 3689 2605 3692
rect 2639 3689 2651 3723
rect 2593 3683 2651 3689
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3326 3720 3332 3732
rect 3099 3692 3332 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4246 3680 4252 3732
rect 4304 3680 4310 3732
rect 7006 3680 7012 3732
rect 7064 3680 7070 3732
rect 7466 3680 7472 3732
rect 7524 3680 7530 3732
rect 8386 3680 8392 3732
rect 8444 3680 8450 3732
rect 9122 3680 9128 3732
rect 9180 3680 9186 3732
rect 9769 3723 9827 3729
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 9858 3720 9864 3732
rect 9815 3692 9864 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10410 3680 10416 3732
rect 10468 3680 10474 3732
rect 11146 3720 11152 3732
rect 10520 3692 11152 3720
rect 2498 3612 2504 3664
rect 2556 3652 2562 3664
rect 3418 3652 3424 3664
rect 2556 3624 3424 3652
rect 2556 3612 2562 3624
rect 3418 3612 3424 3624
rect 3476 3612 3482 3664
rect 4614 3652 4620 3664
rect 3712 3624 4620 3652
rect 3712 3584 3740 3624
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 5810 3612 5816 3664
rect 5868 3652 5874 3664
rect 10520 3652 10548 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 18279 3723 18337 3729
rect 18279 3689 18291 3723
rect 18325 3720 18337 3723
rect 20070 3720 20076 3732
rect 18325 3692 20076 3720
rect 18325 3689 18337 3692
rect 18279 3683 18337 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 20312 3692 21864 3720
rect 20312 3680 20318 3692
rect 18598 3652 18604 3664
rect 5868 3624 10548 3652
rect 10612 3624 18604 3652
rect 5868 3612 5874 3624
rect 1964 3556 3740 3584
rect 3973 3587 4031 3593
rect 1964 3525 1992 3556
rect 3973 3553 3985 3587
rect 4019 3584 4031 3587
rect 4798 3584 4804 3596
rect 4019 3556 4804 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 4798 3544 4804 3556
rect 4856 3584 4862 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 4856 3556 4905 3584
rect 4856 3544 4862 3556
rect 4893 3553 4905 3556
rect 4939 3553 4951 3587
rect 4893 3547 4951 3553
rect 5166 3544 5172 3596
rect 5224 3544 5230 3596
rect 6089 3587 6147 3593
rect 6089 3553 6101 3587
rect 6135 3584 6147 3587
rect 7006 3584 7012 3596
rect 6135 3556 7012 3584
rect 6135 3553 6147 3556
rect 6089 3547 6147 3553
rect 7006 3544 7012 3556
rect 7064 3584 7070 3596
rect 7064 3556 7696 3584
rect 7064 3544 7070 3556
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 2682 3516 2688 3528
rect 2280 3488 2688 3516
rect 2280 3476 2286 3488
rect 2682 3476 2688 3488
rect 2740 3516 2746 3528
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2740 3488 3249 3516
rect 2740 3476 2746 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4430 3516 4436 3528
rect 3651 3488 4436 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 6270 3516 6276 3528
rect 5592 3488 6276 3516
rect 5592 3476 5598 3488
rect 6270 3476 6276 3488
rect 6328 3516 6334 3528
rect 7668 3525 7696 3556
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 6328 3488 6377 3516
rect 6328 3476 6334 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3485 7711 3519
rect 8478 3516 8484 3528
rect 7653 3479 7711 3485
rect 8036 3488 8484 3516
rect 3418 3408 3424 3460
rect 3476 3448 3482 3460
rect 8036 3448 8064 3488
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9582 3516 9588 3528
rect 9355 3488 9588 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10134 3516 10140 3528
rect 9999 3488 10140 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10612 3525 10640 3624
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 18874 3612 18880 3664
rect 18932 3652 18938 3664
rect 21836 3652 21864 3692
rect 21910 3680 21916 3732
rect 21968 3720 21974 3732
rect 22925 3723 22983 3729
rect 22925 3720 22937 3723
rect 21968 3692 22937 3720
rect 21968 3680 21974 3692
rect 22925 3689 22937 3692
rect 22971 3689 22983 3723
rect 22925 3683 22983 3689
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 24029 3723 24087 3729
rect 24029 3720 24041 3723
rect 23532 3692 24041 3720
rect 23532 3680 23538 3692
rect 24029 3689 24041 3692
rect 24075 3689 24087 3723
rect 24029 3683 24087 3689
rect 23198 3652 23204 3664
rect 18932 3624 21772 3652
rect 21836 3624 23204 3652
rect 18932 3612 18938 3624
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 12526 3584 12532 3596
rect 11103 3556 12532 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12802 3544 12808 3596
rect 12860 3544 12866 3596
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18690 3584 18696 3596
rect 18095 3556 18696 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 19058 3544 19064 3596
rect 19116 3584 19122 3596
rect 21744 3593 21772 3624
rect 23198 3612 23204 3624
rect 23256 3612 23262 3664
rect 21729 3587 21787 3593
rect 19116 3556 21404 3584
rect 19116 3544 19122 3556
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 14182 3516 14188 3528
rect 12483 3488 14188 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 3476 3420 8064 3448
rect 8113 3451 8171 3457
rect 3476 3408 3482 3420
rect 8113 3417 8125 3451
rect 8159 3448 8171 3451
rect 8159 3420 9352 3448
rect 8159 3417 8171 3420
rect 8113 3411 8171 3417
rect 9324 3392 9352 3420
rect 9398 3408 9404 3460
rect 9456 3448 9462 3460
rect 10612 3448 10640 3479
rect 9456 3420 10640 3448
rect 11348 3448 11376 3479
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 15930 3516 15936 3528
rect 14507 3488 15936 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 17310 3516 17316 3528
rect 16347 3488 17316 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 19576 3488 20484 3516
rect 19576 3476 19582 3488
rect 14550 3448 14556 3460
rect 11348 3420 14556 3448
rect 9456 3408 9462 3420
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 20349 3451 20407 3457
rect 20349 3448 20361 3451
rect 18340 3420 20361 3448
rect 18340 3392 18368 3420
rect 20349 3417 20361 3420
rect 20395 3417 20407 3451
rect 20456 3448 20484 3488
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20772 3488 21281 3516
rect 20772 3476 20778 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21376 3516 21404 3556
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 21376 3488 23397 3516
rect 21269 3479 21327 3485
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 24578 3476 24584 3528
rect 24636 3476 24642 3528
rect 22370 3448 22376 3460
rect 20456 3420 22376 3448
rect 20349 3411 20407 3417
rect 22370 3408 22376 3420
rect 22428 3408 22434 3460
rect 1486 3340 1492 3392
rect 1544 3340 1550 3392
rect 9306 3340 9312 3392
rect 9364 3340 9370 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 18230 3380 18236 3392
rect 11204 3352 18236 3380
rect 11204 3340 11210 3352
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 18322 3340 18328 3392
rect 18380 3340 18386 3392
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 21358 3380 21364 3392
rect 19576 3352 21364 3380
rect 19576 3340 19582 3352
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 22830 3380 22836 3392
rect 22152 3352 22836 3380
rect 22152 3340 22158 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 24578 3340 24584 3392
rect 24636 3380 24642 3392
rect 25225 3383 25283 3389
rect 25225 3380 25237 3383
rect 24636 3352 25237 3380
rect 24636 3340 24642 3352
rect 25225 3349 25237 3352
rect 25271 3349 25283 3383
rect 25225 3343 25283 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 7285 3179 7343 3185
rect 7285 3176 7297 3179
rect 6052 3148 7297 3176
rect 6052 3136 6058 3148
rect 7285 3145 7297 3148
rect 7331 3145 7343 3179
rect 7285 3139 7343 3145
rect 9398 3136 9404 3188
rect 9456 3136 9462 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 10008 3148 10333 3176
rect 10008 3136 10014 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 10321 3139 10379 3145
rect 10520 3148 17264 3176
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3384 3012 3433 3040
rect 3384 3000 3390 3012
rect 3421 3009 3433 3012
rect 3467 3040 3479 3043
rect 3510 3040 3516 3052
rect 3467 3012 3516 3040
rect 3467 3009 3479 3012
rect 3421 3003 3479 3009
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 5350 3040 5356 3052
rect 3743 3012 5356 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 10520 3049 10548 3148
rect 10962 3068 10968 3120
rect 11020 3108 11026 3120
rect 11238 3108 11244 3120
rect 11020 3080 11244 3108
rect 11020 3068 11026 3080
rect 11238 3068 11244 3080
rect 11296 3068 11302 3120
rect 14182 3108 14188 3120
rect 13188 3080 14188 3108
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7800 3012 7849 3040
rect 7800 3000 7806 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2972 1823 2975
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 1811 2944 2145 2972
rect 1811 2941 1823 2944
rect 1765 2935 1823 2941
rect 2133 2941 2145 2944
rect 2179 2972 2191 2975
rect 2590 2972 2596 2984
rect 2179 2944 2596 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 5166 2972 5172 2984
rect 4755 2944 5172 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8113 2975 8171 2981
rect 8113 2972 8125 2975
rect 7708 2944 8125 2972
rect 7708 2932 7714 2944
rect 8113 2941 8125 2944
rect 8159 2941 8171 2975
rect 8113 2935 8171 2941
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9876 2972 9904 3003
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11422 3000 11428 3052
rect 11480 3040 11486 3052
rect 11698 3040 11704 3052
rect 11480 3012 11704 3040
rect 11480 3000 11486 3012
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 13188 3049 13216 3080
rect 14182 3068 14188 3080
rect 14240 3108 14246 3120
rect 16298 3108 16304 3120
rect 14240 3080 16304 3108
rect 14240 3068 14246 3080
rect 16298 3068 16304 3080
rect 16356 3068 16362 3120
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14700 3012 14841 3040
rect 14700 3000 14706 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17126 3040 17132 3052
rect 17083 3012 17132 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17236 3040 17264 3148
rect 17494 3136 17500 3188
rect 17552 3176 17558 3188
rect 17552 3148 19380 3176
rect 17552 3136 17558 3148
rect 17310 3068 17316 3120
rect 17368 3108 17374 3120
rect 19352 3108 19380 3148
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21269 3179 21327 3185
rect 21269 3176 21281 3179
rect 20956 3148 21281 3176
rect 20956 3136 20962 3148
rect 21269 3145 21281 3148
rect 21315 3145 21327 3179
rect 22925 3179 22983 3185
rect 22925 3176 22937 3179
rect 21269 3139 21327 3145
rect 21376 3148 22937 3176
rect 21376 3108 21404 3148
rect 22925 3145 22937 3148
rect 22971 3145 22983 3179
rect 22925 3139 22983 3145
rect 23661 3179 23719 3185
rect 23661 3145 23673 3179
rect 23707 3176 23719 3179
rect 23842 3176 23848 3188
rect 23707 3148 23848 3176
rect 23707 3145 23719 3148
rect 23661 3139 23719 3145
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 24118 3136 24124 3188
rect 24176 3176 24182 3188
rect 24213 3179 24271 3185
rect 24213 3176 24225 3179
rect 24176 3148 24225 3176
rect 24176 3136 24182 3148
rect 24213 3145 24225 3148
rect 24259 3145 24271 3179
rect 24213 3139 24271 3145
rect 24581 3179 24639 3185
rect 24581 3145 24593 3179
rect 24627 3176 24639 3179
rect 24670 3176 24676 3188
rect 24627 3148 24676 3176
rect 24627 3145 24639 3148
rect 24581 3139 24639 3145
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 17368 3080 19288 3108
rect 19352 3080 21404 3108
rect 17368 3068 17374 3080
rect 18414 3040 18420 3052
rect 17236 3012 18420 3040
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3040 18935 3043
rect 18966 3040 18972 3052
rect 18923 3012 18972 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 11790 2972 11796 2984
rect 9263 2944 11796 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2972 12035 2975
rect 12023 2944 12434 2972
rect 12023 2941 12035 2944
rect 11977 2935 12035 2941
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 1854 2904 1860 2916
rect 1719 2876 1860 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 7834 2864 7840 2916
rect 7892 2904 7898 2916
rect 9033 2907 9091 2913
rect 7892 2876 8984 2904
rect 7892 2864 7898 2876
rect 4893 2839 4951 2845
rect 4893 2805 4905 2839
rect 4939 2836 4951 2839
rect 6638 2836 6644 2848
rect 4939 2808 6644 2836
rect 4939 2805 4951 2808
rect 4893 2799 4951 2805
rect 6638 2796 6644 2808
rect 6696 2836 6702 2848
rect 8846 2836 8852 2848
rect 6696 2808 8852 2836
rect 6696 2796 6702 2808
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 8956 2836 8984 2876
rect 9033 2873 9045 2907
rect 9079 2904 9091 2907
rect 9582 2904 9588 2916
rect 9079 2876 9588 2904
rect 9079 2873 9091 2876
rect 9033 2867 9091 2873
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 9677 2907 9735 2913
rect 9677 2873 9689 2907
rect 9723 2904 9735 2907
rect 12406 2904 12434 2944
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15896 2944 17325 2972
rect 15896 2932 15902 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19260 2972 19288 3080
rect 21542 3068 21548 3120
rect 21600 3108 21606 3120
rect 22186 3108 22192 3120
rect 21600 3080 22192 3108
rect 21600 3068 21606 3080
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 22278 3068 22284 3120
rect 22336 3068 22342 3120
rect 22830 3068 22836 3120
rect 22888 3108 22894 3120
rect 25041 3111 25099 3117
rect 25041 3108 25053 3111
rect 22888 3080 25053 3108
rect 22888 3068 22894 3080
rect 25041 3077 25053 3080
rect 25087 3077 25099 3111
rect 25041 3071 25099 3077
rect 19886 3000 19892 3052
rect 19944 3040 19950 3052
rect 20625 3043 20683 3049
rect 20625 3040 20637 3043
rect 19944 3012 20637 3040
rect 19944 3000 19950 3012
rect 20625 3009 20637 3012
rect 20671 3040 20683 3043
rect 21910 3040 21916 3052
rect 20671 3012 21916 3040
rect 20671 3009 20683 3012
rect 20625 3003 20683 3009
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 22002 3000 22008 3052
rect 22060 3040 22066 3052
rect 22097 3043 22155 3049
rect 22097 3040 22109 3043
rect 22060 3012 22109 3040
rect 22060 3000 22066 3012
rect 22097 3009 22109 3012
rect 22143 3040 22155 3043
rect 22143 3012 22416 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 22278 2972 22284 2984
rect 19260 2944 22284 2972
rect 19153 2935 19211 2941
rect 14458 2904 14464 2916
rect 9723 2876 11100 2904
rect 12406 2876 14464 2904
rect 9723 2873 9735 2876
rect 9677 2867 9735 2873
rect 9950 2836 9956 2848
rect 8956 2808 9956 2836
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10962 2796 10968 2848
rect 11020 2796 11026 2848
rect 11072 2836 11100 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 19168 2904 19196 2935
rect 22278 2932 22284 2944
rect 22336 2932 22342 2984
rect 22388 2972 22416 3012
rect 22646 3000 22652 3052
rect 22704 3040 22710 3052
rect 23569 3043 23627 3049
rect 23569 3040 23581 3043
rect 22704 3012 23581 3040
rect 22704 3000 22710 3012
rect 23569 3009 23581 3012
rect 23615 3009 23627 3043
rect 23569 3003 23627 3009
rect 24210 3000 24216 3052
rect 24268 3040 24274 3052
rect 24765 3043 24823 3049
rect 24765 3040 24777 3043
rect 24268 3012 24777 3040
rect 24268 3000 24274 3012
rect 24765 3009 24777 3012
rect 24811 3040 24823 3043
rect 25225 3043 25283 3049
rect 25225 3040 25237 3043
rect 24811 3012 25237 3040
rect 24811 3009 24823 3012
rect 24765 3003 24823 3009
rect 25225 3009 25237 3012
rect 25271 3009 25283 3043
rect 25225 3003 25283 3009
rect 24029 2975 24087 2981
rect 24029 2972 24041 2975
rect 22388 2944 24041 2972
rect 24029 2941 24041 2944
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 16632 2876 19196 2904
rect 16632 2864 16638 2876
rect 15010 2836 15016 2848
rect 11072 2808 15016 2836
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 17310 2836 17316 2848
rect 15160 2808 17316 2836
rect 15160 2796 15166 2808
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 17678 2796 17684 2848
rect 17736 2836 17742 2848
rect 19886 2836 19892 2848
rect 17736 2808 19892 2836
rect 17736 2796 17742 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 21542 2836 21548 2848
rect 20763 2808 21548 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 4614 2592 4620 2644
rect 4672 2592 4678 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 7558 2632 7564 2644
rect 7331 2604 7564 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 14918 2632 14924 2644
rect 8435 2604 14924 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 16114 2592 16120 2644
rect 16172 2632 16178 2644
rect 16172 2604 16574 2632
rect 16172 2592 16178 2604
rect 9766 2564 9772 2576
rect 2884 2536 9772 2564
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2593 2499 2651 2505
rect 2593 2496 2605 2499
rect 2363 2468 2605 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2593 2465 2605 2468
rect 2639 2496 2651 2499
rect 2774 2496 2780 2508
rect 2639 2468 2780 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 2884 2505 2912 2536
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 12158 2524 12164 2576
rect 12216 2564 12222 2576
rect 16301 2567 16359 2573
rect 16301 2564 16313 2567
rect 12216 2536 16313 2564
rect 12216 2524 12222 2536
rect 16301 2533 16313 2536
rect 16347 2533 16359 2567
rect 16546 2564 16574 2604
rect 18690 2592 18696 2644
rect 18748 2592 18754 2644
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 22002 2632 22008 2644
rect 20036 2604 22008 2632
rect 20036 2592 20042 2604
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22186 2564 22192 2576
rect 16546 2536 22192 2564
rect 16301 2527 16359 2533
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 5408 2468 5457 2496
rect 5408 2456 5414 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 13906 2496 13912 2508
rect 5445 2459 5503 2465
rect 12544 2468 13912 2496
rect 1854 2388 1860 2440
rect 1912 2388 1918 2440
rect 2958 2388 2964 2440
rect 3016 2428 3022 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3016 2400 3985 2428
rect 3016 2388 3022 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5215 2400 5580 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5552 2304 5580 2400
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8754 2428 8760 2440
rect 8619 2400 8760 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9306 2388 9312 2440
rect 9364 2388 9370 2440
rect 9953 2431 10011 2437
rect 9953 2397 9965 2431
rect 9999 2428 10011 2431
rect 11885 2431 11943 2437
rect 9999 2400 11100 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 10962 2320 10968 2372
rect 11020 2320 11026 2372
rect 11072 2360 11100 2400
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12158 2428 12164 2440
rect 11931 2400 12164 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12544 2437 12572 2468
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 14182 2456 14188 2508
rect 14240 2456 14246 2508
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 15930 2456 15936 2508
rect 15988 2496 15994 2508
rect 16117 2499 16175 2505
rect 16117 2496 16129 2499
rect 15988 2468 16129 2496
rect 15988 2456 15994 2468
rect 16117 2465 16129 2468
rect 16163 2465 16175 2499
rect 16117 2459 16175 2465
rect 17310 2456 17316 2508
rect 17368 2456 17374 2508
rect 18800 2468 19748 2496
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13780 2400 14473 2428
rect 13780 2388 13786 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 12434 2360 12440 2372
rect 11072 2332 12440 2360
rect 12434 2320 12440 2332
rect 12492 2320 12498 2372
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 1670 2252 1676 2304
rect 1728 2252 1734 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 6086 2292 6092 2304
rect 5592 2264 6092 2292
rect 5592 2252 5598 2264
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 7834 2292 7840 2304
rect 7791 2264 7840 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 9122 2252 9128 2304
rect 9180 2252 9186 2304
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 16022 2292 16028 2304
rect 11747 2264 16028 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 18800 2292 18828 2468
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19426 2428 19432 2440
rect 18923 2400 19432 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 19720 2428 19748 2468
rect 19886 2456 19892 2508
rect 19944 2456 19950 2508
rect 25225 2499 25283 2505
rect 25225 2496 25237 2499
rect 19996 2468 25237 2496
rect 19996 2428 20024 2468
rect 25225 2465 25237 2468
rect 25271 2465 25283 2499
rect 25225 2459 25283 2465
rect 19720 2400 20024 2428
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 21453 2431 21511 2437
rect 21453 2428 21465 2431
rect 20588 2400 21465 2428
rect 20588 2388 20594 2400
rect 21453 2397 21465 2400
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 22002 2388 22008 2440
rect 22060 2388 22066 2440
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 22336 2400 22937 2428
rect 22336 2388 22342 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 19242 2320 19248 2372
rect 19300 2360 19306 2372
rect 23845 2363 23903 2369
rect 23845 2360 23857 2363
rect 19300 2332 23857 2360
rect 19300 2320 19306 2332
rect 23845 2329 23857 2332
rect 23891 2329 23903 2363
rect 23845 2323 23903 2329
rect 16448 2264 18828 2292
rect 16448 2252 16454 2264
rect 21266 2252 21272 2304
rect 21324 2252 21330 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 1728 2060 2774 2088
rect 1728 2048 1734 2060
rect 2746 2020 2774 2060
rect 9122 2048 9128 2100
rect 9180 2088 9186 2100
rect 17586 2088 17592 2100
rect 9180 2060 17592 2088
rect 9180 2048 9186 2060
rect 17586 2048 17592 2060
rect 17644 2048 17650 2100
rect 19426 2048 19432 2100
rect 19484 2088 19490 2100
rect 24486 2088 24492 2100
rect 19484 2060 24492 2088
rect 19484 2048 19490 2060
rect 24486 2048 24492 2060
rect 24544 2048 24550 2100
rect 11514 2020 11520 2032
rect 2746 1992 11520 2020
rect 11514 1980 11520 1992
rect 11572 1980 11578 2032
rect 11054 1912 11060 1964
rect 11112 1952 11118 1964
rect 21266 1952 21272 1964
rect 11112 1924 21272 1952
rect 11112 1912 11118 1924
rect 21266 1912 21272 1924
rect 21324 1912 21330 1964
rect 3970 1844 3976 1896
rect 4028 1884 4034 1896
rect 6178 1884 6184 1896
rect 4028 1856 6184 1884
rect 4028 1844 4034 1856
rect 6178 1844 6184 1856
rect 6236 1844 6242 1896
rect 7834 1844 7840 1896
rect 7892 1884 7898 1896
rect 15654 1884 15660 1896
rect 7892 1856 15660 1884
rect 7892 1844 7898 1856
rect 15654 1844 15660 1856
rect 15712 1844 15718 1896
rect 8754 1776 8760 1828
rect 8812 1816 8818 1828
rect 10318 1816 10324 1828
rect 8812 1788 10324 1816
rect 8812 1776 8818 1788
rect 10318 1776 10324 1788
rect 10376 1776 10382 1828
rect 10962 1776 10968 1828
rect 11020 1816 11026 1828
rect 22094 1816 22100 1828
rect 11020 1788 22100 1816
rect 11020 1776 11026 1788
rect 22094 1776 22100 1788
rect 22152 1776 22158 1828
rect 9306 1708 9312 1760
rect 9364 1748 9370 1760
rect 11054 1748 11060 1760
rect 9364 1720 11060 1748
rect 9364 1708 9370 1720
rect 11054 1708 11060 1720
rect 11112 1708 11118 1760
rect 20254 1232 20260 1284
rect 20312 1272 20318 1284
rect 20806 1272 20812 1284
rect 20312 1244 20812 1272
rect 20312 1232 20318 1244
rect 20806 1232 20812 1244
rect 20864 1232 20870 1284
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 16212 54272 16264 54324
rect 8576 54204 8628 54256
rect 4068 54136 4120 54188
rect 4804 54179 4856 54188
rect 4804 54145 4813 54179
rect 4813 54145 4847 54179
rect 4847 54145 4856 54179
rect 4804 54136 4856 54145
rect 7380 54179 7432 54188
rect 7380 54145 7389 54179
rect 7389 54145 7423 54179
rect 7423 54145 7432 54179
rect 7380 54136 7432 54145
rect 9588 54179 9640 54188
rect 9588 54145 9597 54179
rect 9597 54145 9631 54179
rect 9631 54145 9640 54179
rect 9588 54136 9640 54145
rect 11704 54136 11756 54188
rect 14464 54179 14516 54188
rect 14464 54145 14473 54179
rect 14473 54145 14507 54179
rect 14507 54145 14516 54179
rect 14464 54136 14516 54145
rect 14832 54136 14884 54188
rect 16212 54136 16264 54188
rect 17960 54179 18012 54188
rect 17960 54145 17969 54179
rect 17969 54145 18003 54179
rect 18003 54145 18012 54179
rect 17960 54136 18012 54145
rect 2412 54068 2464 54120
rect 5172 54111 5224 54120
rect 5172 54077 5181 54111
rect 5181 54077 5215 54111
rect 5215 54077 5224 54111
rect 5172 54068 5224 54077
rect 7840 54111 7892 54120
rect 7840 54077 7849 54111
rect 7849 54077 7883 54111
rect 7883 54077 7892 54111
rect 7840 54068 7892 54077
rect 9312 54068 9364 54120
rect 12348 54068 12400 54120
rect 18972 54315 19024 54324
rect 18972 54281 18981 54315
rect 18981 54281 19015 54315
rect 19015 54281 19024 54315
rect 18972 54272 19024 54281
rect 20720 54179 20772 54188
rect 20720 54145 20729 54179
rect 20729 54145 20763 54179
rect 20763 54145 20772 54179
rect 20720 54136 20772 54145
rect 21732 54136 21784 54188
rect 25872 54136 25924 54188
rect 16764 54000 16816 54052
rect 13544 53932 13596 53984
rect 15568 53932 15620 53984
rect 17040 53932 17092 53984
rect 18604 53975 18656 53984
rect 18604 53941 18613 53975
rect 18613 53941 18647 53975
rect 18647 53941 18656 53975
rect 18604 53932 18656 53941
rect 18788 54000 18840 54052
rect 24676 53932 24728 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 13452 53728 13504 53780
rect 10692 53660 10744 53712
rect 1032 53592 1084 53644
rect 3792 53592 3844 53644
rect 6552 53592 6604 53644
rect 4160 53567 4212 53576
rect 4160 53533 4169 53567
rect 4169 53533 4203 53567
rect 4203 53533 4212 53567
rect 4160 53524 4212 53533
rect 7840 53524 7892 53576
rect 10692 53524 10744 53576
rect 14464 53728 14516 53780
rect 17868 53728 17920 53780
rect 23296 53592 23348 53644
rect 15568 53567 15620 53576
rect 15568 53533 15577 53567
rect 15577 53533 15611 53567
rect 15611 53533 15620 53567
rect 15568 53524 15620 53533
rect 17040 53567 17092 53576
rect 17040 53533 17049 53567
rect 17049 53533 17083 53567
rect 17083 53533 17092 53567
rect 17040 53524 17092 53533
rect 18604 53524 18656 53576
rect 22284 53567 22336 53576
rect 22284 53533 22293 53567
rect 22293 53533 22327 53567
rect 22327 53533 22336 53567
rect 22284 53524 22336 53533
rect 23388 53524 23440 53576
rect 24676 53567 24728 53576
rect 24676 53533 24685 53567
rect 24685 53533 24719 53567
rect 24719 53533 24728 53567
rect 24676 53524 24728 53533
rect 5540 53456 5592 53508
rect 21456 53456 21508 53508
rect 14740 53388 14792 53440
rect 15660 53388 15712 53440
rect 17684 53431 17736 53440
rect 17684 53397 17693 53431
rect 17693 53397 17727 53431
rect 17727 53397 17736 53431
rect 17684 53388 17736 53397
rect 19984 53388 20036 53440
rect 23940 53431 23992 53440
rect 23940 53397 23949 53431
rect 23949 53397 23983 53431
rect 23983 53397 23992 53431
rect 23940 53388 23992 53397
rect 24584 53388 24636 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 4068 53184 4120 53236
rect 23296 53227 23348 53236
rect 23296 53193 23305 53227
rect 23305 53193 23339 53227
rect 23339 53193 23348 53227
rect 23296 53184 23348 53193
rect 23388 53227 23440 53236
rect 23388 53193 23397 53227
rect 23397 53193 23431 53227
rect 23431 53193 23440 53227
rect 23388 53184 23440 53193
rect 24768 53184 24820 53236
rect 25320 53227 25372 53236
rect 25320 53193 25329 53227
rect 25329 53193 25363 53227
rect 25363 53193 25372 53227
rect 25320 53184 25372 53193
rect 7748 53048 7800 53100
rect 22284 52980 22336 53032
rect 24860 52980 24912 53032
rect 25504 52955 25556 52964
rect 25504 52921 25513 52955
rect 25513 52921 25547 52955
rect 25547 52921 25556 52955
rect 25504 52912 25556 52921
rect 23664 52844 23716 52896
rect 24676 52887 24728 52896
rect 24676 52853 24685 52887
rect 24685 52853 24719 52887
rect 24719 52853 24728 52887
rect 24676 52844 24728 52853
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 4160 52640 4212 52692
rect 24492 52683 24544 52692
rect 24492 52649 24501 52683
rect 24501 52649 24535 52683
rect 24535 52649 24544 52683
rect 24492 52640 24544 52649
rect 23848 52572 23900 52624
rect 9496 52436 9548 52488
rect 24492 52436 24544 52488
rect 25964 52436 26016 52488
rect 24952 52411 25004 52420
rect 24952 52377 24961 52411
rect 24961 52377 24995 52411
rect 24995 52377 25004 52411
rect 24952 52368 25004 52377
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 24952 52096 25004 52148
rect 24584 52003 24636 52012
rect 24584 51969 24593 52003
rect 24593 51969 24627 52003
rect 24627 51969 24636 52003
rect 24584 51960 24636 51969
rect 25504 51960 25556 52012
rect 24584 51756 24636 51808
rect 25228 51799 25280 51808
rect 25228 51765 25237 51799
rect 25237 51765 25271 51799
rect 25271 51765 25280 51799
rect 25228 51756 25280 51765
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 7380 51552 7432 51604
rect 7840 51484 7892 51536
rect 4804 51348 4856 51400
rect 8484 51391 8536 51400
rect 8484 51357 8493 51391
rect 8493 51357 8527 51391
rect 8527 51357 8536 51391
rect 8484 51348 8536 51357
rect 10508 51348 10560 51400
rect 10784 51280 10836 51332
rect 24952 51323 25004 51332
rect 24952 51289 24961 51323
rect 24961 51289 24995 51323
rect 24995 51289 25004 51323
rect 24952 51280 25004 51289
rect 25780 51280 25832 51332
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 25044 50872 25096 50924
rect 24952 50668 25004 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 5540 50464 5592 50516
rect 8392 50464 8444 50516
rect 9588 50507 9640 50516
rect 9588 50473 9597 50507
rect 9597 50473 9631 50507
rect 9631 50473 9640 50507
rect 9588 50464 9640 50473
rect 7748 50396 7800 50448
rect 8576 50328 8628 50380
rect 24584 50303 24636 50312
rect 24584 50269 24593 50303
rect 24593 50269 24627 50303
rect 24627 50269 24636 50303
rect 24584 50260 24636 50269
rect 9588 50192 9640 50244
rect 23388 50124 23440 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 19800 49852 19852 49904
rect 24216 49784 24268 49836
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 24216 49419 24268 49428
rect 24216 49385 24225 49419
rect 24225 49385 24259 49419
rect 24259 49385 24268 49419
rect 24216 49376 24268 49385
rect 24768 49376 24820 49428
rect 10692 49351 10744 49360
rect 10692 49317 10701 49351
rect 10701 49317 10735 49351
rect 10735 49317 10744 49351
rect 10692 49308 10744 49317
rect 11704 49351 11756 49360
rect 11704 49317 11713 49351
rect 11713 49317 11747 49351
rect 11747 49317 11756 49351
rect 11704 49308 11756 49317
rect 24860 49172 24912 49224
rect 10232 49104 10284 49156
rect 10876 49104 10928 49156
rect 25136 49036 25188 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 9128 48832 9180 48884
rect 24860 48832 24912 48884
rect 25136 48807 25188 48816
rect 25136 48773 25145 48807
rect 25145 48773 25179 48807
rect 25179 48773 25188 48807
rect 25136 48764 25188 48773
rect 8300 48628 8352 48680
rect 8392 48671 8444 48680
rect 8392 48637 8401 48671
rect 8401 48637 8435 48671
rect 8435 48637 8444 48671
rect 8392 48628 8444 48637
rect 9956 48560 10008 48612
rect 26148 48560 26200 48612
rect 9128 48492 9180 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 7748 48084 7800 48136
rect 23388 48127 23440 48136
rect 23388 48093 23397 48127
rect 23397 48093 23431 48127
rect 23431 48093 23440 48127
rect 23388 48084 23440 48093
rect 24860 48084 24912 48136
rect 13728 47948 13780 48000
rect 24032 47991 24084 48000
rect 24032 47957 24041 47991
rect 24041 47957 24075 47991
rect 24075 47957 24084 47991
rect 24032 47948 24084 47957
rect 25136 47948 25188 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9220 47744 9272 47796
rect 9496 47744 9548 47796
rect 24860 47744 24912 47796
rect 8576 47676 8628 47728
rect 10968 47676 11020 47728
rect 25136 47719 25188 47728
rect 25136 47685 25145 47719
rect 25145 47685 25179 47719
rect 25179 47685 25188 47719
rect 25136 47676 25188 47685
rect 16212 47540 16264 47592
rect 25228 47540 25280 47592
rect 25688 47472 25740 47524
rect 8300 47404 8352 47456
rect 9496 47447 9548 47456
rect 9496 47413 9505 47447
rect 9505 47413 9539 47447
rect 9539 47413 9548 47447
rect 9496 47404 9548 47413
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 26516 47132 26568 47184
rect 9220 46996 9272 47048
rect 25320 47039 25372 47048
rect 25320 47005 25329 47039
rect 25329 47005 25363 47039
rect 25363 47005 25372 47039
rect 25320 46996 25372 47005
rect 13636 46928 13688 46980
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 10784 46699 10836 46708
rect 10784 46665 10793 46699
rect 10793 46665 10827 46699
rect 10827 46665 10836 46699
rect 10784 46656 10836 46665
rect 10968 46656 11020 46708
rect 13636 46656 13688 46708
rect 14740 46631 14792 46640
rect 14740 46597 14749 46631
rect 14749 46597 14783 46631
rect 14783 46597 14792 46631
rect 14740 46588 14792 46597
rect 10784 46520 10836 46572
rect 25320 46563 25372 46572
rect 25320 46529 25329 46563
rect 25329 46529 25363 46563
rect 25363 46529 25372 46563
rect 25320 46520 25372 46529
rect 15752 46495 15804 46504
rect 15752 46461 15761 46495
rect 15761 46461 15795 46495
rect 15795 46461 15804 46495
rect 15752 46452 15804 46461
rect 10784 46384 10836 46436
rect 10416 46359 10468 46368
rect 10416 46325 10425 46359
rect 10425 46325 10459 46359
rect 10459 46325 10468 46359
rect 10416 46316 10468 46325
rect 15476 46316 15528 46368
rect 21180 46316 21232 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 8484 46155 8536 46164
rect 8484 46121 8493 46155
rect 8493 46121 8527 46155
rect 8527 46121 8536 46155
rect 8484 46112 8536 46121
rect 7748 45976 7800 46028
rect 15660 46019 15712 46028
rect 15660 45985 15669 46019
rect 15669 45985 15703 46019
rect 15703 45985 15712 46019
rect 15660 45976 15712 45985
rect 16488 46019 16540 46028
rect 16488 45985 16497 46019
rect 16497 45985 16531 46019
rect 16531 45985 16540 46019
rect 16488 45976 16540 45985
rect 7840 45908 7892 45960
rect 12808 45908 12860 45960
rect 25320 45951 25372 45960
rect 25320 45917 25329 45951
rect 25329 45917 25363 45951
rect 25363 45917 25372 45951
rect 25320 45908 25372 45917
rect 15476 45840 15528 45892
rect 14924 45772 14976 45824
rect 25044 45772 25096 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 10508 45500 10560 45552
rect 12808 45500 12860 45552
rect 13544 45543 13596 45552
rect 13544 45509 13553 45543
rect 13553 45509 13587 45543
rect 13587 45509 13596 45543
rect 13544 45500 13596 45509
rect 13728 45500 13780 45552
rect 25412 45432 25464 45484
rect 14556 45407 14608 45416
rect 14556 45373 14565 45407
rect 14565 45373 14599 45407
rect 14599 45373 14608 45407
rect 14556 45364 14608 45373
rect 25228 45228 25280 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 9496 45024 9548 45076
rect 16028 44956 16080 45008
rect 24952 44956 25004 45008
rect 9956 44888 10008 44940
rect 9128 44863 9180 44872
rect 9128 44829 9137 44863
rect 9137 44829 9171 44863
rect 9171 44829 9180 44863
rect 9128 44820 9180 44829
rect 9680 44752 9732 44804
rect 17684 44888 17736 44940
rect 11520 44752 11572 44804
rect 14924 44752 14976 44804
rect 17500 44795 17552 44804
rect 17500 44761 17509 44795
rect 17509 44761 17543 44795
rect 17543 44761 17552 44795
rect 17500 44752 17552 44761
rect 25320 44752 25372 44804
rect 10416 44684 10468 44736
rect 11704 44684 11756 44736
rect 25504 44684 25556 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 9588 44523 9640 44532
rect 9588 44489 9597 44523
rect 9597 44489 9631 44523
rect 9631 44489 9640 44523
rect 9588 44480 9640 44489
rect 13820 44480 13872 44532
rect 17500 44480 17552 44532
rect 25320 44523 25372 44532
rect 25320 44489 25329 44523
rect 25329 44489 25363 44523
rect 25363 44489 25372 44523
rect 25320 44480 25372 44489
rect 9220 44344 9272 44396
rect 10784 44344 10836 44396
rect 24676 44387 24728 44396
rect 24676 44353 24685 44387
rect 24685 44353 24719 44387
rect 24719 44353 24728 44387
rect 24676 44344 24728 44353
rect 9312 44276 9364 44328
rect 10508 44208 10560 44260
rect 10692 44183 10744 44192
rect 10692 44149 10701 44183
rect 10701 44149 10735 44183
rect 10735 44149 10744 44183
rect 10692 44140 10744 44149
rect 10968 44140 11020 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 24032 43800 24084 43852
rect 19524 43732 19576 43784
rect 21088 43664 21140 43716
rect 25320 43664 25372 43716
rect 21364 43596 21416 43648
rect 24860 43596 24912 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 25320 43435 25372 43444
rect 25320 43401 25329 43435
rect 25329 43401 25363 43435
rect 25363 43401 25372 43435
rect 25320 43392 25372 43401
rect 24952 43256 25004 43308
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 24860 42780 24912 42832
rect 10232 42755 10284 42764
rect 10232 42721 10241 42755
rect 10241 42721 10275 42755
rect 10275 42721 10284 42755
rect 10232 42712 10284 42721
rect 21272 42712 21324 42764
rect 8944 42644 8996 42696
rect 10600 42644 10652 42696
rect 24860 42644 24912 42696
rect 25136 42508 25188 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 9680 42304 9732 42356
rect 24860 42304 24912 42356
rect 11520 42236 11572 42288
rect 25136 42279 25188 42288
rect 25136 42245 25145 42279
rect 25145 42245 25179 42279
rect 25179 42245 25188 42279
rect 25136 42236 25188 42245
rect 9128 42100 9180 42152
rect 9680 42143 9732 42152
rect 9680 42109 9689 42143
rect 9689 42109 9723 42143
rect 9723 42109 9732 42143
rect 9680 42100 9732 42109
rect 10692 42100 10744 42152
rect 15844 42032 15896 42084
rect 24492 42032 24544 42084
rect 11520 42007 11572 42016
rect 11520 41973 11529 42007
rect 11529 41973 11563 42007
rect 11563 41973 11572 42007
rect 11520 41964 11572 41973
rect 11704 42007 11756 42016
rect 11704 41973 11713 42007
rect 11713 41973 11747 42007
rect 11747 41973 11756 42007
rect 11704 41964 11756 41973
rect 21732 41964 21784 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 10876 41803 10928 41812
rect 10876 41769 10885 41803
rect 10885 41769 10919 41803
rect 10919 41769 10928 41803
rect 10876 41760 10928 41769
rect 10968 41624 11020 41676
rect 10232 41599 10284 41608
rect 10232 41565 10241 41599
rect 10241 41565 10275 41599
rect 10275 41565 10284 41599
rect 10232 41556 10284 41565
rect 16856 41556 16908 41608
rect 21456 41556 21508 41608
rect 24860 41556 24912 41608
rect 25320 41463 25372 41472
rect 25320 41429 25329 41463
rect 25329 41429 25363 41463
rect 25363 41429 25372 41463
rect 25320 41420 25372 41429
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 24768 41259 24820 41268
rect 24768 41225 24777 41259
rect 24777 41225 24811 41259
rect 24811 41225 24820 41259
rect 24768 41216 24820 41225
rect 25320 41148 25372 41200
rect 24860 40876 24912 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 25320 40511 25372 40520
rect 25320 40477 25329 40511
rect 25329 40477 25363 40511
rect 25363 40477 25372 40511
rect 25320 40468 25372 40477
rect 25412 40332 25464 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 23296 40128 23348 40180
rect 25320 40035 25372 40044
rect 25320 40001 25329 40035
rect 25329 40001 25363 40035
rect 25363 40001 25372 40035
rect 25320 39992 25372 40001
rect 17040 39924 17092 39976
rect 23664 39924 23716 39976
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 10692 39584 10744 39636
rect 13820 39584 13872 39636
rect 25320 39423 25372 39432
rect 25320 39389 25329 39423
rect 25329 39389 25363 39423
rect 25363 39389 25372 39423
rect 25320 39380 25372 39389
rect 24124 39244 24176 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 24768 38700 24820 38752
rect 25044 38700 25096 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 16948 38496 17000 38548
rect 19984 38496 20036 38548
rect 25320 38224 25372 38276
rect 25872 38156 25924 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 7840 37952 7892 38004
rect 25320 37995 25372 38004
rect 25320 37961 25329 37995
rect 25329 37961 25363 37995
rect 25363 37961 25372 37995
rect 25320 37952 25372 37961
rect 9036 37884 9088 37936
rect 15752 37884 15804 37936
rect 8852 37859 8904 37868
rect 8852 37825 8861 37859
rect 8861 37825 8895 37859
rect 8895 37825 8904 37859
rect 8852 37816 8904 37825
rect 24860 37816 24912 37868
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 25596 37272 25648 37324
rect 25320 37136 25372 37188
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 25320 36907 25372 36916
rect 25320 36873 25329 36907
rect 25329 36873 25363 36907
rect 25363 36873 25372 36907
rect 25320 36864 25372 36873
rect 24952 36728 25004 36780
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 24768 36116 24820 36168
rect 24676 35980 24728 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 11704 35776 11756 35828
rect 21180 35819 21232 35828
rect 21180 35785 21189 35819
rect 21189 35785 21223 35819
rect 21223 35785 21232 35819
rect 21180 35776 21232 35785
rect 25136 35776 25188 35828
rect 11520 35751 11572 35760
rect 11520 35717 11529 35751
rect 11529 35717 11563 35751
rect 11563 35717 11572 35751
rect 11520 35708 11572 35717
rect 12348 35708 12400 35760
rect 22100 35708 22152 35760
rect 22008 35640 22060 35692
rect 24676 35683 24728 35692
rect 24676 35649 24685 35683
rect 24685 35649 24719 35683
rect 24719 35649 24728 35683
rect 24676 35640 24728 35649
rect 25320 35683 25372 35692
rect 25320 35649 25329 35683
rect 25329 35649 25363 35683
rect 25363 35649 25372 35683
rect 25320 35640 25372 35649
rect 10048 35572 10100 35624
rect 21180 35572 21232 35624
rect 22560 35615 22612 35624
rect 22560 35581 22569 35615
rect 22569 35581 22603 35615
rect 22603 35581 22612 35615
rect 22560 35572 22612 35581
rect 19064 35504 19116 35556
rect 9680 35436 9732 35488
rect 11796 35479 11848 35488
rect 11796 35445 11805 35479
rect 11805 35445 11839 35479
rect 11839 35445 11848 35479
rect 11796 35436 11848 35445
rect 20628 35504 20680 35556
rect 24584 35436 24636 35488
rect 26056 35436 26108 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 25320 35275 25372 35284
rect 25320 35241 25329 35275
rect 25329 35241 25363 35275
rect 25363 35241 25372 35275
rect 25320 35232 25372 35241
rect 22744 35096 22796 35148
rect 24860 35028 24912 35080
rect 22008 34892 22060 34944
rect 22192 34892 22244 34944
rect 25228 34960 25280 35012
rect 22468 34892 22520 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 21088 34688 21140 34740
rect 25228 34688 25280 34740
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 9312 34144 9364 34196
rect 23020 34144 23072 34196
rect 11796 34008 11848 34060
rect 19708 34008 19760 34060
rect 22284 34008 22336 34060
rect 9220 33940 9272 33992
rect 19432 33983 19484 33992
rect 19432 33949 19441 33983
rect 19441 33949 19475 33983
rect 19475 33949 19484 33983
rect 19432 33940 19484 33949
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 15384 33872 15436 33924
rect 19984 33872 20036 33924
rect 21088 33872 21140 33924
rect 22376 33872 22428 33924
rect 19248 33804 19300 33856
rect 21180 33847 21232 33856
rect 21180 33813 21189 33847
rect 21189 33813 21223 33847
rect 21223 33813 21232 33847
rect 21180 33804 21232 33813
rect 23204 33804 23256 33856
rect 24216 33804 24268 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 22560 33600 22612 33652
rect 23204 33600 23256 33652
rect 23572 33600 23624 33652
rect 21088 33532 21140 33584
rect 21916 33532 21968 33584
rect 19524 33507 19576 33516
rect 19524 33473 19533 33507
rect 19533 33473 19567 33507
rect 19567 33473 19576 33507
rect 19524 33464 19576 33473
rect 22284 33532 22336 33584
rect 22376 33532 22428 33584
rect 22376 33396 22428 33448
rect 23020 33396 23072 33448
rect 19248 33303 19300 33312
rect 19248 33269 19257 33303
rect 19257 33269 19291 33303
rect 19291 33269 19300 33303
rect 19248 33260 19300 33269
rect 19984 33260 20036 33312
rect 20536 33260 20588 33312
rect 23848 33260 23900 33312
rect 24768 33260 24820 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 16580 33056 16632 33108
rect 16120 32963 16172 32972
rect 16120 32929 16129 32963
rect 16129 32929 16163 32963
rect 16163 32929 16172 32963
rect 21364 33056 21416 33108
rect 21916 33099 21968 33108
rect 21916 33065 21925 33099
rect 21925 33065 21959 33099
rect 21959 33065 21968 33099
rect 21916 33056 21968 33065
rect 22376 33056 22428 33108
rect 22744 33056 22796 33108
rect 19892 32988 19944 33040
rect 21824 32988 21876 33040
rect 16120 32920 16172 32929
rect 16580 32852 16632 32904
rect 17316 32852 17368 32904
rect 17224 32784 17276 32836
rect 19432 32852 19484 32904
rect 17500 32784 17552 32836
rect 19892 32827 19944 32836
rect 19892 32793 19901 32827
rect 19901 32793 19935 32827
rect 19935 32793 19944 32827
rect 19892 32784 19944 32793
rect 12624 32716 12676 32768
rect 22284 32963 22336 32972
rect 22284 32929 22293 32963
rect 22293 32929 22327 32963
rect 22327 32929 22336 32963
rect 22284 32920 22336 32929
rect 25136 32920 25188 32972
rect 25228 32963 25280 32972
rect 25228 32929 25237 32963
rect 25237 32929 25271 32963
rect 25271 32929 25280 32963
rect 25228 32920 25280 32929
rect 25412 32852 25464 32904
rect 21916 32784 21968 32836
rect 23848 32784 23900 32836
rect 23480 32716 23532 32768
rect 24860 32716 24912 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 15384 32487 15436 32496
rect 15384 32453 15393 32487
rect 15393 32453 15427 32487
rect 15427 32453 15436 32487
rect 15384 32444 15436 32453
rect 17500 32512 17552 32564
rect 19248 32512 19300 32564
rect 17592 32444 17644 32496
rect 19616 32444 19668 32496
rect 25136 32512 25188 32564
rect 25412 32512 25464 32564
rect 21088 32444 21140 32496
rect 22284 32444 22336 32496
rect 21824 32376 21876 32428
rect 24032 32444 24084 32496
rect 13360 32308 13412 32360
rect 16764 32308 16816 32360
rect 17132 32308 17184 32360
rect 21180 32308 21232 32360
rect 25228 32308 25280 32360
rect 19432 32172 19484 32224
rect 19708 32172 19760 32224
rect 20904 32172 20956 32224
rect 21824 32172 21876 32224
rect 25964 32172 26016 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 9496 31968 9548 32020
rect 16488 31968 16540 32020
rect 18512 31968 18564 32020
rect 19248 31968 19300 32020
rect 24032 32011 24084 32020
rect 24032 31977 24041 32011
rect 24041 31977 24075 32011
rect 24075 31977 24084 32011
rect 24032 31968 24084 31977
rect 24860 31968 24912 32020
rect 25320 31968 25372 32020
rect 12532 31900 12584 31952
rect 20812 31900 20864 31952
rect 22744 31900 22796 31952
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 16672 31832 16724 31884
rect 17592 31832 17644 31884
rect 17684 31832 17736 31884
rect 19708 31875 19760 31884
rect 19708 31841 19717 31875
rect 19717 31841 19751 31875
rect 19751 31841 19760 31875
rect 19708 31832 19760 31841
rect 24124 31900 24176 31952
rect 25044 31900 25096 31952
rect 16764 31807 16816 31816
rect 16764 31773 16773 31807
rect 16773 31773 16807 31807
rect 16807 31773 16816 31807
rect 16764 31764 16816 31773
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 21088 31764 21140 31816
rect 23296 31832 23348 31884
rect 23020 31764 23072 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 19248 31696 19300 31748
rect 17132 31628 17184 31680
rect 20996 31628 21048 31680
rect 22008 31671 22060 31680
rect 22008 31637 22017 31671
rect 22017 31637 22051 31671
rect 22051 31637 22060 31671
rect 22008 31628 22060 31637
rect 22100 31628 22152 31680
rect 22560 31628 22612 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 16672 31467 16724 31476
rect 16672 31433 16681 31467
rect 16681 31433 16715 31467
rect 16715 31433 16724 31467
rect 16672 31424 16724 31433
rect 19708 31424 19760 31476
rect 25136 31424 25188 31476
rect 25504 31424 25556 31476
rect 26148 31424 26200 31476
rect 15016 31356 15068 31408
rect 19248 31356 19300 31408
rect 22652 31356 22704 31408
rect 23020 31356 23072 31408
rect 24032 31356 24084 31408
rect 16764 31288 16816 31340
rect 21916 31288 21968 31340
rect 22284 31288 22336 31340
rect 25504 31288 25556 31340
rect 13360 31263 13412 31272
rect 13360 31229 13369 31263
rect 13369 31229 13403 31263
rect 13403 31229 13412 31263
rect 13360 31220 13412 31229
rect 16120 31220 16172 31272
rect 17684 31263 17736 31272
rect 17684 31229 17693 31263
rect 17693 31229 17727 31263
rect 17727 31229 17736 31263
rect 17684 31220 17736 31229
rect 18696 31220 18748 31272
rect 22376 31220 22428 31272
rect 15016 31152 15068 31204
rect 13820 31084 13872 31136
rect 22008 31152 22060 31204
rect 22284 31152 22336 31204
rect 18420 31084 18472 31136
rect 19892 31084 19944 31136
rect 21916 31084 21968 31136
rect 22192 31084 22244 31136
rect 23480 31084 23532 31136
rect 25136 31127 25188 31136
rect 25136 31093 25145 31127
rect 25145 31093 25179 31127
rect 25179 31093 25188 31127
rect 25136 31084 25188 31093
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 10232 30880 10284 30932
rect 15384 30880 15436 30932
rect 18512 30923 18564 30932
rect 18512 30889 18521 30923
rect 18521 30889 18555 30923
rect 18555 30889 18564 30923
rect 18512 30880 18564 30889
rect 18696 30880 18748 30932
rect 19248 30880 19300 30932
rect 22652 30880 22704 30932
rect 25504 30923 25556 30932
rect 25504 30889 25513 30923
rect 25513 30889 25547 30923
rect 25547 30889 25556 30923
rect 25504 30880 25556 30889
rect 19432 30744 19484 30796
rect 8760 30676 8812 30728
rect 14096 30676 14148 30728
rect 15384 30676 15436 30728
rect 15108 30651 15160 30660
rect 15108 30617 15117 30651
rect 15117 30617 15151 30651
rect 15151 30617 15160 30651
rect 15108 30608 15160 30617
rect 18420 30608 18472 30660
rect 19248 30608 19300 30660
rect 20996 30651 21048 30660
rect 20996 30617 21005 30651
rect 21005 30617 21039 30651
rect 21039 30617 21048 30651
rect 20996 30608 21048 30617
rect 22376 30608 22428 30660
rect 18696 30540 18748 30592
rect 20076 30583 20128 30592
rect 20076 30549 20085 30583
rect 20085 30549 20119 30583
rect 20119 30549 20128 30583
rect 20076 30540 20128 30549
rect 22652 30608 22704 30660
rect 24032 30540 24084 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 13360 30336 13412 30388
rect 19248 30336 19300 30388
rect 20076 30336 20128 30388
rect 7656 30200 7708 30252
rect 12716 30268 12768 30320
rect 14096 30311 14148 30320
rect 14096 30277 14105 30311
rect 14105 30277 14139 30311
rect 14139 30277 14148 30311
rect 14096 30268 14148 30277
rect 20628 30268 20680 30320
rect 22468 30311 22520 30320
rect 22468 30277 22477 30311
rect 22477 30277 22511 30311
rect 22511 30277 22520 30311
rect 22468 30268 22520 30277
rect 23480 30268 23532 30320
rect 24032 30268 24084 30320
rect 16764 30200 16816 30252
rect 12072 30175 12124 30184
rect 12072 30141 12081 30175
rect 12081 30141 12115 30175
rect 12115 30141 12124 30175
rect 12072 30132 12124 30141
rect 12440 30132 12492 30184
rect 12716 30132 12768 30184
rect 13360 30132 13412 30184
rect 8944 30107 8996 30116
rect 8944 30073 8953 30107
rect 8953 30073 8987 30107
rect 8987 30073 8996 30107
rect 8944 30064 8996 30073
rect 16028 30175 16080 30184
rect 16028 30141 16037 30175
rect 16037 30141 16071 30175
rect 16071 30141 16080 30175
rect 16028 30132 16080 30141
rect 16488 30132 16540 30184
rect 17040 30064 17092 30116
rect 20536 30175 20588 30184
rect 20536 30141 20545 30175
rect 20545 30141 20579 30175
rect 20579 30141 20588 30175
rect 20536 30132 20588 30141
rect 22836 30132 22888 30184
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 23940 30132 23992 30184
rect 25228 30132 25280 30184
rect 11520 29996 11572 30048
rect 13636 29996 13688 30048
rect 15936 29996 15988 30048
rect 16672 30039 16724 30048
rect 16672 30005 16681 30039
rect 16681 30005 16715 30039
rect 16715 30005 16724 30039
rect 16672 29996 16724 30005
rect 16764 29996 16816 30048
rect 19248 29996 19300 30048
rect 20352 29996 20404 30048
rect 23756 29996 23808 30048
rect 25780 29996 25832 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 12072 29792 12124 29844
rect 13820 29792 13872 29844
rect 11428 29656 11480 29708
rect 13360 29656 13412 29708
rect 16028 29656 16080 29708
rect 15292 29588 15344 29640
rect 16488 29767 16540 29776
rect 16488 29733 16497 29767
rect 16497 29733 16531 29767
rect 16531 29733 16540 29767
rect 16488 29724 16540 29733
rect 18696 29792 18748 29844
rect 22836 29792 22888 29844
rect 23756 29724 23808 29776
rect 25688 29724 25740 29776
rect 19340 29656 19392 29708
rect 18420 29588 18472 29640
rect 11152 29520 11204 29572
rect 12716 29520 12768 29572
rect 16488 29520 16540 29572
rect 15016 29452 15068 29504
rect 15200 29495 15252 29504
rect 15200 29461 15209 29495
rect 15209 29461 15243 29495
rect 15243 29461 15252 29495
rect 15200 29452 15252 29461
rect 18880 29588 18932 29640
rect 24860 29656 24912 29708
rect 24584 29588 24636 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 24860 29520 24912 29572
rect 19156 29452 19208 29504
rect 19616 29452 19668 29504
rect 20536 29495 20588 29504
rect 20536 29461 20545 29495
rect 20545 29461 20579 29495
rect 20579 29461 20588 29495
rect 20536 29452 20588 29461
rect 22468 29452 22520 29504
rect 24584 29452 24636 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 8852 29248 8904 29300
rect 12440 29248 12492 29300
rect 12624 29291 12676 29300
rect 12624 29257 12633 29291
rect 12633 29257 12667 29291
rect 12667 29257 12676 29291
rect 12624 29248 12676 29257
rect 13820 29248 13872 29300
rect 13912 29248 13964 29300
rect 10416 29180 10468 29232
rect 10232 29112 10284 29164
rect 10048 29087 10100 29096
rect 10048 29053 10057 29087
rect 10057 29053 10091 29087
rect 10091 29053 10100 29087
rect 10048 29044 10100 29053
rect 11612 29044 11664 29096
rect 15016 29180 15068 29232
rect 13360 29155 13412 29164
rect 13360 29121 13369 29155
rect 13369 29121 13403 29155
rect 13403 29121 13412 29155
rect 13360 29112 13412 29121
rect 15200 29248 15252 29300
rect 16212 29248 16264 29300
rect 19156 29291 19208 29300
rect 19156 29257 19165 29291
rect 19165 29257 19199 29291
rect 19199 29257 19208 29291
rect 19156 29248 19208 29257
rect 20536 29248 20588 29300
rect 23848 29248 23900 29300
rect 25320 29248 25372 29300
rect 15936 29223 15988 29232
rect 15936 29189 15945 29223
rect 15945 29189 15979 29223
rect 15979 29189 15988 29223
rect 15936 29180 15988 29189
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 17316 29155 17368 29164
rect 17316 29121 17325 29155
rect 17325 29121 17359 29155
rect 17359 29121 17368 29155
rect 17316 29112 17368 29121
rect 13636 29044 13688 29096
rect 12256 28976 12308 29028
rect 15200 28976 15252 29028
rect 16580 28976 16632 29028
rect 19064 29180 19116 29232
rect 17500 29112 17552 29164
rect 18420 29112 18472 29164
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 20904 29044 20956 29096
rect 17500 28976 17552 29028
rect 19524 28976 19576 29028
rect 20536 28976 20588 29028
rect 21824 29019 21876 29028
rect 21824 28985 21833 29019
rect 21833 28985 21867 29019
rect 21867 28985 21876 29019
rect 26516 29112 26568 29164
rect 23388 29044 23440 29096
rect 23756 29044 23808 29096
rect 24952 29044 25004 29096
rect 21824 28976 21876 28985
rect 14096 28908 14148 28960
rect 15016 28908 15068 28960
rect 15936 28908 15988 28960
rect 18420 28908 18472 28960
rect 24124 28908 24176 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 10048 28704 10100 28756
rect 12072 28704 12124 28756
rect 14556 28704 14608 28756
rect 11428 28611 11480 28620
rect 11428 28577 11437 28611
rect 11437 28577 11471 28611
rect 11471 28577 11480 28611
rect 11428 28568 11480 28577
rect 14096 28568 14148 28620
rect 16488 28704 16540 28756
rect 18604 28704 18656 28756
rect 18880 28747 18932 28756
rect 18880 28713 18889 28747
rect 18889 28713 18923 28747
rect 18923 28713 18932 28747
rect 18880 28704 18932 28713
rect 23756 28704 23808 28756
rect 15936 28679 15988 28688
rect 15936 28645 15945 28679
rect 15945 28645 15979 28679
rect 15979 28645 15988 28679
rect 15936 28636 15988 28645
rect 21916 28636 21968 28688
rect 23204 28636 23256 28688
rect 15384 28611 15436 28620
rect 15384 28577 15393 28611
rect 15393 28577 15427 28611
rect 15427 28577 15436 28611
rect 15384 28568 15436 28577
rect 18972 28568 19024 28620
rect 20996 28568 21048 28620
rect 23664 28568 23716 28620
rect 24860 28568 24912 28620
rect 25412 28568 25464 28620
rect 15108 28500 15160 28552
rect 18420 28500 18472 28552
rect 19340 28500 19392 28552
rect 20628 28543 20680 28552
rect 20628 28509 20637 28543
rect 20637 28509 20671 28543
rect 20671 28509 20680 28543
rect 20628 28500 20680 28509
rect 23572 28500 23624 28552
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 9680 28432 9732 28484
rect 10968 28432 11020 28484
rect 11520 28364 11572 28416
rect 13544 28407 13596 28416
rect 13544 28373 13553 28407
rect 13553 28373 13587 28407
rect 13587 28373 13596 28407
rect 13544 28364 13596 28373
rect 14832 28407 14884 28416
rect 14832 28373 14841 28407
rect 14841 28373 14875 28407
rect 14875 28373 14884 28407
rect 14832 28364 14884 28373
rect 20812 28432 20864 28484
rect 20904 28475 20956 28484
rect 20904 28441 20913 28475
rect 20913 28441 20947 28475
rect 20947 28441 20956 28475
rect 20904 28432 20956 28441
rect 16028 28407 16080 28416
rect 16028 28373 16037 28407
rect 16037 28373 16071 28407
rect 16071 28373 16080 28407
rect 16028 28364 16080 28373
rect 19524 28364 19576 28416
rect 19708 28364 19760 28416
rect 22284 28364 22336 28416
rect 23204 28407 23256 28416
rect 23204 28373 23213 28407
rect 23213 28373 23247 28407
rect 23247 28373 23256 28407
rect 23204 28364 23256 28373
rect 23940 28407 23992 28416
rect 23940 28373 23949 28407
rect 23949 28373 23983 28407
rect 23983 28373 23992 28407
rect 23940 28364 23992 28373
rect 24400 28364 24452 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 13544 28160 13596 28212
rect 15016 28160 15068 28212
rect 15844 28160 15896 28212
rect 17132 28160 17184 28212
rect 11060 28092 11112 28144
rect 18512 28160 18564 28212
rect 18788 28160 18840 28212
rect 19708 28203 19760 28212
rect 19708 28169 19717 28203
rect 19717 28169 19751 28203
rect 19751 28169 19760 28203
rect 19708 28160 19760 28169
rect 24216 28160 24268 28212
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 12624 27956 12676 28008
rect 20628 28092 20680 28144
rect 22560 28092 22612 28144
rect 16304 28024 16356 28076
rect 18420 28024 18472 28076
rect 10784 27888 10836 27940
rect 10968 27863 11020 27872
rect 10968 27829 10977 27863
rect 10977 27829 11011 27863
rect 11011 27829 11020 27863
rect 10968 27820 11020 27829
rect 15384 27888 15436 27940
rect 13820 27820 13872 27872
rect 16304 27863 16356 27872
rect 16304 27829 16313 27863
rect 16313 27829 16347 27863
rect 16347 27829 16356 27863
rect 16304 27820 16356 27829
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 17408 27999 17460 28008
rect 17408 27965 17417 27999
rect 17417 27965 17451 27999
rect 17451 27965 17460 27999
rect 17408 27956 17460 27965
rect 18144 27956 18196 28008
rect 17684 27888 17736 27940
rect 21824 28024 21876 28076
rect 23388 28092 23440 28144
rect 23480 28135 23532 28144
rect 23480 28101 23489 28135
rect 23489 28101 23523 28135
rect 23523 28101 23532 28135
rect 23480 28092 23532 28101
rect 23940 28092 23992 28144
rect 20536 27888 20588 27940
rect 22560 27999 22612 28008
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 22560 27956 22612 27965
rect 17592 27820 17644 27872
rect 18512 27863 18564 27872
rect 18512 27829 18521 27863
rect 18521 27829 18555 27863
rect 18555 27829 18564 27863
rect 18512 27820 18564 27829
rect 20996 27820 21048 27872
rect 22376 27820 22428 27872
rect 23296 27820 23348 27872
rect 25228 27863 25280 27872
rect 25228 27829 25237 27863
rect 25237 27829 25271 27863
rect 25271 27829 25280 27863
rect 25228 27820 25280 27829
rect 25964 27820 26016 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 9036 27548 9088 27600
rect 3424 27480 3476 27532
rect 11428 27616 11480 27668
rect 12624 27659 12676 27668
rect 12624 27625 12633 27659
rect 12633 27625 12667 27659
rect 12667 27625 12676 27659
rect 12624 27616 12676 27625
rect 11796 27548 11848 27600
rect 13084 27548 13136 27600
rect 15108 27616 15160 27668
rect 16488 27659 16540 27668
rect 16488 27625 16497 27659
rect 16497 27625 16531 27659
rect 16531 27625 16540 27659
rect 16488 27616 16540 27625
rect 19984 27616 20036 27668
rect 23664 27616 23716 27668
rect 19432 27548 19484 27600
rect 23480 27548 23532 27600
rect 24768 27548 24820 27600
rect 10784 27523 10836 27532
rect 10784 27489 10793 27523
rect 10793 27489 10827 27523
rect 10827 27489 10836 27523
rect 10784 27480 10836 27489
rect 10876 27480 10928 27532
rect 11980 27480 12032 27532
rect 13360 27480 13412 27532
rect 14740 27480 14792 27532
rect 17776 27480 17828 27532
rect 23388 27480 23440 27532
rect 23848 27480 23900 27532
rect 25044 27523 25096 27532
rect 25044 27489 25053 27523
rect 25053 27489 25087 27523
rect 25087 27489 25096 27523
rect 25044 27480 25096 27489
rect 11888 27412 11940 27464
rect 12624 27412 12676 27464
rect 14832 27412 14884 27464
rect 16488 27412 16540 27464
rect 18144 27412 18196 27464
rect 23940 27412 23992 27464
rect 10876 27344 10928 27396
rect 13820 27344 13872 27396
rect 16028 27344 16080 27396
rect 12072 27276 12124 27328
rect 12164 27276 12216 27328
rect 12624 27276 12676 27328
rect 13728 27276 13780 27328
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 15660 27276 15712 27328
rect 16488 27276 16540 27328
rect 19892 27344 19944 27396
rect 22376 27387 22428 27396
rect 22376 27353 22385 27387
rect 22385 27353 22419 27387
rect 22419 27353 22428 27387
rect 22376 27344 22428 27353
rect 23664 27344 23716 27396
rect 19432 27276 19484 27328
rect 20076 27276 20128 27328
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 25044 27276 25096 27328
rect 25228 27276 25280 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 9036 26936 9088 26988
rect 9772 27072 9824 27124
rect 10876 27072 10928 27124
rect 11796 27072 11848 27124
rect 11980 27072 12032 27124
rect 15568 27072 15620 27124
rect 16856 27072 16908 27124
rect 10968 27004 11020 27056
rect 11888 27004 11940 27056
rect 13268 27004 13320 27056
rect 13636 27004 13688 27056
rect 16580 27004 16632 27056
rect 19248 27072 19300 27124
rect 22744 27072 22796 27124
rect 24768 27072 24820 27124
rect 7564 26868 7616 26920
rect 12164 26936 12216 26988
rect 12808 26936 12860 26988
rect 13084 26979 13136 26988
rect 13084 26945 13093 26979
rect 13093 26945 13127 26979
rect 13127 26945 13136 26979
rect 13084 26936 13136 26945
rect 15936 26936 15988 26988
rect 18788 27004 18840 27056
rect 22652 26936 22704 26988
rect 11152 26868 11204 26920
rect 9312 26800 9364 26852
rect 15752 26868 15804 26920
rect 22100 26868 22152 26920
rect 22560 26868 22612 26920
rect 23572 27004 23624 27056
rect 23940 27004 23992 27056
rect 23388 26868 23440 26920
rect 25228 26868 25280 26920
rect 11980 26732 12032 26784
rect 14924 26732 14976 26784
rect 18972 26732 19024 26784
rect 20076 26775 20128 26784
rect 20076 26741 20085 26775
rect 20085 26741 20119 26775
rect 20119 26741 20128 26775
rect 20076 26732 20128 26741
rect 21088 26732 21140 26784
rect 22376 26775 22428 26784
rect 22376 26741 22385 26775
rect 22385 26741 22419 26775
rect 22419 26741 22428 26775
rect 22376 26732 22428 26741
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 9404 26528 9456 26580
rect 11612 26528 11664 26580
rect 15752 26528 15804 26580
rect 20996 26528 21048 26580
rect 22100 26528 22152 26580
rect 9772 26392 9824 26444
rect 11060 26392 11112 26444
rect 11888 26460 11940 26512
rect 12716 26460 12768 26512
rect 14280 26460 14332 26512
rect 16028 26460 16080 26512
rect 16764 26460 16816 26512
rect 14832 26435 14884 26444
rect 14832 26401 14841 26435
rect 14841 26401 14875 26435
rect 14875 26401 14884 26435
rect 14832 26392 14884 26401
rect 15476 26392 15528 26444
rect 15936 26392 15988 26444
rect 11336 26324 11388 26376
rect 14740 26324 14792 26376
rect 16672 26367 16724 26376
rect 16672 26333 16681 26367
rect 16681 26333 16715 26367
rect 16715 26333 16724 26367
rect 16672 26324 16724 26333
rect 18788 26460 18840 26512
rect 22008 26460 22060 26512
rect 25044 26528 25096 26580
rect 22560 26460 22612 26512
rect 19432 26435 19484 26444
rect 19432 26401 19441 26435
rect 19441 26401 19475 26435
rect 19475 26401 19484 26435
rect 19432 26392 19484 26401
rect 20996 26392 21048 26444
rect 21640 26392 21692 26444
rect 22192 26392 22244 26444
rect 24860 26460 24912 26512
rect 17868 26324 17920 26376
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 25044 26392 25096 26444
rect 25504 26324 25556 26376
rect 8944 26256 8996 26308
rect 9404 26299 9456 26308
rect 9404 26265 9413 26299
rect 9413 26265 9447 26299
rect 9447 26265 9456 26299
rect 9404 26256 9456 26265
rect 15936 26256 15988 26308
rect 16304 26256 16356 26308
rect 16948 26256 17000 26308
rect 21088 26256 21140 26308
rect 14464 26188 14516 26240
rect 15016 26188 15068 26240
rect 15844 26188 15896 26240
rect 17224 26231 17276 26240
rect 17224 26197 17233 26231
rect 17233 26197 17267 26231
rect 17267 26197 17276 26231
rect 17224 26188 17276 26197
rect 18328 26188 18380 26240
rect 22284 26188 22336 26240
rect 22836 26256 22888 26308
rect 23020 26231 23072 26240
rect 23020 26197 23029 26231
rect 23029 26197 23063 26231
rect 23063 26197 23072 26231
rect 23020 26188 23072 26197
rect 25136 26256 25188 26308
rect 25964 26256 26016 26308
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 9496 26027 9548 26036
rect 9496 25993 9505 26027
rect 9505 25993 9539 26027
rect 9539 25993 9548 26027
rect 9496 25984 9548 25993
rect 12624 26027 12676 26036
rect 12624 25993 12633 26027
rect 12633 25993 12667 26027
rect 12667 25993 12676 26027
rect 12624 25984 12676 25993
rect 13912 25959 13964 25968
rect 13912 25925 13921 25959
rect 13921 25925 13955 25959
rect 13955 25925 13964 25959
rect 13912 25916 13964 25925
rect 15108 25916 15160 25968
rect 16856 26027 16908 26036
rect 16856 25993 16865 26027
rect 16865 25993 16899 26027
rect 16899 25993 16908 26027
rect 16856 25984 16908 25993
rect 17040 25984 17092 26036
rect 18328 25984 18380 26036
rect 18604 25984 18656 26036
rect 12624 25848 12676 25900
rect 19616 25916 19668 25968
rect 17132 25848 17184 25900
rect 22284 25984 22336 26036
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 23020 25984 23072 26036
rect 24952 25984 25004 26036
rect 4804 25780 4856 25832
rect 11152 25780 11204 25832
rect 14096 25823 14148 25832
rect 14096 25789 14105 25823
rect 14105 25789 14139 25823
rect 14139 25789 14148 25823
rect 14096 25780 14148 25789
rect 13452 25712 13504 25764
rect 11796 25644 11848 25696
rect 12440 25644 12492 25696
rect 13544 25687 13596 25696
rect 13544 25653 13553 25687
rect 13553 25653 13587 25687
rect 13587 25653 13596 25687
rect 13544 25644 13596 25653
rect 13820 25644 13872 25696
rect 15384 25823 15436 25832
rect 15384 25789 15393 25823
rect 15393 25789 15427 25823
rect 15427 25789 15436 25823
rect 15384 25780 15436 25789
rect 18696 25780 18748 25832
rect 26240 25916 26292 25968
rect 22008 25780 22060 25832
rect 23480 25891 23532 25900
rect 23480 25857 23489 25891
rect 23489 25857 23523 25891
rect 23523 25857 23532 25891
rect 23480 25848 23532 25857
rect 22744 25780 22796 25832
rect 22836 25780 22888 25832
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 17408 25687 17460 25696
rect 17408 25653 17417 25687
rect 17417 25653 17451 25687
rect 17451 25653 17460 25687
rect 17408 25644 17460 25653
rect 21548 25687 21600 25696
rect 21548 25653 21557 25687
rect 21557 25653 21591 25687
rect 21591 25653 21600 25687
rect 21548 25644 21600 25653
rect 21640 25644 21692 25696
rect 22100 25644 22152 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 11704 25440 11756 25492
rect 17960 25440 18012 25492
rect 18604 25440 18656 25492
rect 21088 25440 21140 25492
rect 22836 25440 22888 25492
rect 23480 25440 23532 25492
rect 12440 25372 12492 25424
rect 15384 25372 15436 25424
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 14740 25304 14792 25356
rect 14832 25347 14884 25356
rect 14832 25313 14841 25347
rect 14841 25313 14875 25347
rect 14875 25313 14884 25347
rect 14832 25304 14884 25313
rect 12716 25236 12768 25288
rect 13360 25236 13412 25288
rect 16856 25304 16908 25356
rect 15200 25236 15252 25288
rect 17592 25236 17644 25288
rect 18420 25236 18472 25288
rect 15292 25168 15344 25220
rect 18604 25168 18656 25220
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 20076 25168 20128 25220
rect 25320 25236 25372 25288
rect 12716 25100 12768 25152
rect 15384 25100 15436 25152
rect 15568 25100 15620 25152
rect 16304 25100 16356 25152
rect 18512 25100 18564 25152
rect 19892 25143 19944 25152
rect 19892 25109 19901 25143
rect 19901 25109 19935 25143
rect 19935 25109 19944 25143
rect 19892 25100 19944 25109
rect 23848 25211 23900 25220
rect 23848 25177 23857 25211
rect 23857 25177 23891 25211
rect 23891 25177 23900 25211
rect 23848 25168 23900 25177
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 7288 24760 7340 24812
rect 10140 24828 10192 24880
rect 11244 24896 11296 24948
rect 14832 24896 14884 24948
rect 15292 24896 15344 24948
rect 15476 24939 15528 24948
rect 15476 24905 15485 24939
rect 15485 24905 15519 24939
rect 15519 24905 15528 24939
rect 15476 24896 15528 24905
rect 17224 24939 17276 24948
rect 17224 24905 17233 24939
rect 17233 24905 17267 24939
rect 17267 24905 17276 24939
rect 17224 24896 17276 24905
rect 17868 24896 17920 24948
rect 22284 24896 22336 24948
rect 13544 24828 13596 24880
rect 18328 24828 18380 24880
rect 11152 24760 11204 24812
rect 12164 24803 12216 24812
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 12808 24760 12860 24812
rect 16396 24760 16448 24812
rect 11060 24692 11112 24744
rect 13912 24692 13964 24744
rect 14740 24735 14792 24744
rect 14740 24701 14749 24735
rect 14749 24701 14783 24735
rect 14783 24701 14792 24735
rect 14740 24692 14792 24701
rect 15108 24692 15160 24744
rect 11060 24556 11112 24608
rect 11244 24556 11296 24608
rect 15200 24624 15252 24676
rect 15384 24735 15436 24744
rect 15384 24701 15393 24735
rect 15393 24701 15427 24735
rect 15427 24701 15436 24735
rect 15384 24692 15436 24701
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 18696 24760 18748 24812
rect 22468 24871 22520 24880
rect 22468 24837 22477 24871
rect 22477 24837 22511 24871
rect 22511 24837 22520 24871
rect 22468 24828 22520 24837
rect 23940 24828 23992 24880
rect 19432 24760 19484 24812
rect 21088 24760 21140 24812
rect 22192 24760 22244 24812
rect 23480 24760 23532 24812
rect 18604 24735 18656 24744
rect 18604 24701 18613 24735
rect 18613 24701 18647 24735
rect 18647 24701 18656 24735
rect 18604 24692 18656 24701
rect 20444 24692 20496 24744
rect 19064 24624 19116 24676
rect 15936 24556 15988 24608
rect 17868 24556 17920 24608
rect 19340 24556 19392 24608
rect 23296 24692 23348 24744
rect 22836 24624 22888 24676
rect 23388 24624 23440 24676
rect 25044 24692 25096 24744
rect 25228 24692 25280 24744
rect 22652 24556 22704 24608
rect 23940 24556 23992 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 9496 24216 9548 24268
rect 12716 24352 12768 24404
rect 12900 24352 12952 24404
rect 20444 24352 20496 24404
rect 22652 24352 22704 24404
rect 11336 24327 11388 24336
rect 11336 24293 11345 24327
rect 11345 24293 11379 24327
rect 11379 24293 11388 24327
rect 11336 24284 11388 24293
rect 23388 24284 23440 24336
rect 11060 24216 11112 24268
rect 12348 24216 12400 24268
rect 18972 24216 19024 24268
rect 19432 24259 19484 24268
rect 19432 24225 19441 24259
rect 19441 24225 19475 24259
rect 19475 24225 19484 24259
rect 19432 24216 19484 24225
rect 22192 24216 22244 24268
rect 22284 24216 22336 24268
rect 22652 24216 22704 24268
rect 7840 24148 7892 24200
rect 17684 24191 17736 24200
rect 17684 24157 17693 24191
rect 17693 24157 17727 24191
rect 17727 24157 17736 24191
rect 17684 24148 17736 24157
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 25412 24148 25464 24200
rect 9864 24080 9916 24132
rect 9588 24012 9640 24064
rect 11336 24080 11388 24132
rect 11980 24080 12032 24132
rect 13544 24080 13596 24132
rect 18880 24080 18932 24132
rect 19708 24123 19760 24132
rect 19708 24089 19717 24123
rect 19717 24089 19751 24123
rect 19751 24089 19760 24123
rect 19708 24080 19760 24089
rect 21088 24080 21140 24132
rect 11060 24012 11112 24064
rect 13912 24012 13964 24064
rect 14096 24055 14148 24064
rect 14096 24021 14105 24055
rect 14105 24021 14139 24055
rect 14139 24021 14148 24055
rect 14096 24012 14148 24021
rect 18512 24012 18564 24064
rect 20536 24012 20588 24064
rect 22284 24012 22336 24064
rect 23572 24012 23624 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 9680 23808 9732 23860
rect 9588 23740 9640 23792
rect 7840 23672 7892 23724
rect 10416 23851 10468 23860
rect 10416 23817 10425 23851
rect 10425 23817 10459 23851
rect 10459 23817 10468 23851
rect 10416 23808 10468 23817
rect 13820 23808 13872 23860
rect 11152 23740 11204 23792
rect 11796 23740 11848 23792
rect 14280 23740 14332 23792
rect 14924 23851 14976 23860
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 16580 23808 16632 23860
rect 17316 23851 17368 23860
rect 17316 23817 17325 23851
rect 17325 23817 17359 23851
rect 17359 23817 17368 23851
rect 17316 23808 17368 23817
rect 18880 23851 18932 23860
rect 18880 23817 18889 23851
rect 18889 23817 18923 23851
rect 18923 23817 18932 23851
rect 18880 23808 18932 23817
rect 10692 23672 10744 23724
rect 10048 23604 10100 23656
rect 13728 23715 13780 23724
rect 13728 23681 13737 23715
rect 13737 23681 13771 23715
rect 13771 23681 13780 23715
rect 13728 23672 13780 23681
rect 14188 23672 14240 23724
rect 14924 23672 14976 23724
rect 16672 23672 16724 23724
rect 19248 23740 19300 23792
rect 11152 23536 11204 23588
rect 12900 23536 12952 23588
rect 13912 23604 13964 23656
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 19800 23808 19852 23860
rect 21916 23808 21968 23860
rect 23848 23808 23900 23860
rect 25044 23808 25096 23860
rect 25320 23808 25372 23860
rect 19708 23740 19760 23792
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 19984 23672 20036 23724
rect 15476 23536 15528 23588
rect 19708 23647 19760 23656
rect 19708 23613 19717 23647
rect 19717 23613 19751 23647
rect 19751 23613 19760 23647
rect 19708 23604 19760 23613
rect 22744 23740 22796 23792
rect 23204 23740 23256 23792
rect 23940 23740 23992 23792
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 22192 23672 22244 23724
rect 20996 23647 21048 23656
rect 20996 23613 21005 23647
rect 21005 23613 21039 23647
rect 21039 23613 21048 23647
rect 20996 23604 21048 23613
rect 22652 23672 22704 23724
rect 22836 23604 22888 23656
rect 23572 23604 23624 23656
rect 21180 23536 21232 23588
rect 9588 23468 9640 23520
rect 10140 23468 10192 23520
rect 12808 23468 12860 23520
rect 17316 23468 17368 23520
rect 19892 23468 19944 23520
rect 20260 23468 20312 23520
rect 22284 23468 22336 23520
rect 23940 23468 23992 23520
rect 25320 23511 25372 23520
rect 25320 23477 25329 23511
rect 25329 23477 25363 23511
rect 25363 23477 25372 23511
rect 25320 23468 25372 23477
rect 25964 23468 26016 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 10600 23264 10652 23316
rect 9588 23196 9640 23248
rect 6184 23128 6236 23180
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 11796 23171 11848 23180
rect 11796 23137 11805 23171
rect 11805 23137 11839 23171
rect 11839 23137 11848 23171
rect 11796 23128 11848 23137
rect 12532 23196 12584 23248
rect 14280 23060 14332 23112
rect 14372 23103 14424 23112
rect 14372 23069 14381 23103
rect 14381 23069 14415 23103
rect 14415 23069 14424 23103
rect 14372 23060 14424 23069
rect 15660 23060 15712 23112
rect 13268 22992 13320 23044
rect 14924 22992 14976 23044
rect 17224 23264 17276 23316
rect 25780 23264 25832 23316
rect 18328 23196 18380 23248
rect 18420 23196 18472 23248
rect 18696 23128 18748 23180
rect 19708 23128 19760 23180
rect 20444 23128 20496 23180
rect 20812 23128 20864 23180
rect 25412 23128 25464 23180
rect 18236 23103 18288 23112
rect 18236 23069 18245 23103
rect 18245 23069 18279 23103
rect 18279 23069 18288 23103
rect 18236 23060 18288 23069
rect 18788 23060 18840 23112
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 21640 23060 21692 23112
rect 16856 22992 16908 23044
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 25688 23060 25740 23112
rect 24860 22992 24912 23044
rect 25320 22992 25372 23044
rect 10600 22924 10652 22976
rect 10876 22924 10928 22976
rect 12072 22924 12124 22976
rect 16580 22924 16632 22976
rect 19064 22924 19116 22976
rect 22100 22924 22152 22976
rect 23480 22924 23532 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 10140 22763 10192 22772
rect 10140 22729 10149 22763
rect 10149 22729 10183 22763
rect 10183 22729 10192 22763
rect 10140 22720 10192 22729
rect 11336 22720 11388 22772
rect 14372 22720 14424 22772
rect 14924 22720 14976 22772
rect 16856 22763 16908 22772
rect 16856 22729 16865 22763
rect 16865 22729 16899 22763
rect 16899 22729 16908 22763
rect 16856 22720 16908 22729
rect 18788 22763 18840 22772
rect 18788 22729 18797 22763
rect 18797 22729 18831 22763
rect 18831 22729 18840 22763
rect 18788 22720 18840 22729
rect 19064 22720 19116 22772
rect 19616 22720 19668 22772
rect 23388 22720 23440 22772
rect 7840 22584 7892 22636
rect 9496 22584 9548 22636
rect 14096 22652 14148 22704
rect 14648 22652 14700 22704
rect 21456 22652 21508 22704
rect 25136 22695 25188 22704
rect 25136 22661 25145 22695
rect 25145 22661 25179 22695
rect 25179 22661 25188 22695
rect 25136 22652 25188 22661
rect 12348 22627 12400 22636
rect 12348 22593 12357 22627
rect 12357 22593 12391 22627
rect 12391 22593 12400 22627
rect 12348 22584 12400 22593
rect 15292 22584 15344 22636
rect 19064 22584 19116 22636
rect 19708 22584 19760 22636
rect 11244 22516 11296 22568
rect 13360 22516 13412 22568
rect 18788 22516 18840 22568
rect 18972 22516 19024 22568
rect 6920 22380 6972 22432
rect 11796 22448 11848 22500
rect 21548 22584 21600 22636
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 23848 22584 23900 22636
rect 19984 22516 20036 22568
rect 23296 22559 23348 22568
rect 23296 22525 23305 22559
rect 23305 22525 23339 22559
rect 23339 22525 23348 22559
rect 23296 22516 23348 22525
rect 13268 22380 13320 22432
rect 14096 22423 14148 22432
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 14096 22380 14148 22389
rect 14648 22423 14700 22432
rect 14648 22389 14657 22423
rect 14657 22389 14691 22423
rect 14691 22389 14700 22423
rect 14648 22380 14700 22389
rect 16120 22380 16172 22432
rect 17040 22380 17092 22432
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 11060 22176 11112 22228
rect 8668 22040 8720 22092
rect 11520 22108 11572 22160
rect 10416 21972 10468 22024
rect 11796 21904 11848 21956
rect 9220 21836 9272 21888
rect 10140 21836 10192 21888
rect 10416 21879 10468 21888
rect 10416 21845 10425 21879
rect 10425 21845 10459 21879
rect 10459 21845 10468 21879
rect 10416 21836 10468 21845
rect 10784 21836 10836 21888
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 16212 22176 16264 22228
rect 12808 22108 12860 22160
rect 15568 22108 15620 22160
rect 14096 21972 14148 22024
rect 16764 22040 16816 22092
rect 23112 22176 23164 22228
rect 23388 22176 23440 22228
rect 18604 22040 18656 22092
rect 20536 22108 20588 22160
rect 25228 22176 25280 22228
rect 22192 22040 22244 22092
rect 23020 22040 23072 22092
rect 24860 22040 24912 22092
rect 17500 21972 17552 22024
rect 23204 21972 23256 22024
rect 15292 21904 15344 21956
rect 12348 21879 12400 21888
rect 12348 21845 12357 21879
rect 12357 21845 12391 21879
rect 12391 21845 12400 21879
rect 12348 21836 12400 21845
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 16212 21836 16264 21888
rect 17132 21836 17184 21888
rect 21364 21904 21416 21956
rect 22284 21904 22336 21956
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20076 21836 20128 21845
rect 20168 21879 20220 21888
rect 20168 21845 20177 21879
rect 20177 21845 20211 21879
rect 20211 21845 20220 21879
rect 20168 21836 20220 21845
rect 23296 21836 23348 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 10232 21632 10284 21684
rect 10968 21632 11020 21684
rect 11060 21632 11112 21684
rect 11796 21632 11848 21684
rect 12716 21632 12768 21684
rect 8576 21564 8628 21616
rect 9496 21564 9548 21616
rect 12164 21564 12216 21616
rect 14648 21564 14700 21616
rect 15660 21632 15712 21684
rect 19064 21632 19116 21684
rect 20076 21632 20128 21684
rect 22560 21632 22612 21684
rect 22744 21632 22796 21684
rect 23112 21632 23164 21684
rect 14832 21564 14884 21616
rect 9956 21496 10008 21548
rect 10692 21496 10744 21548
rect 8392 21428 8444 21480
rect 8852 21428 8904 21480
rect 12440 21496 12492 21548
rect 15752 21496 15804 21548
rect 18788 21564 18840 21616
rect 20168 21564 20220 21616
rect 23204 21564 23256 21616
rect 24032 21564 24084 21616
rect 22008 21496 22060 21548
rect 22468 21496 22520 21548
rect 23020 21496 23072 21548
rect 9312 21360 9364 21412
rect 14096 21428 14148 21480
rect 15108 21428 15160 21480
rect 19984 21428 20036 21480
rect 10784 21360 10836 21412
rect 7748 21292 7800 21344
rect 8300 21292 8352 21344
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 10968 21292 11020 21344
rect 15476 21360 15528 21412
rect 20996 21360 21048 21412
rect 22284 21360 22336 21412
rect 22468 21360 22520 21412
rect 14004 21292 14056 21344
rect 15292 21292 15344 21344
rect 18696 21335 18748 21344
rect 18696 21301 18705 21335
rect 18705 21301 18739 21335
rect 18739 21301 18748 21335
rect 18696 21292 18748 21301
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 21916 21292 21968 21344
rect 25412 21428 25464 21480
rect 23572 21292 23624 21344
rect 24032 21292 24084 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 8484 21088 8536 21140
rect 12348 21088 12400 21140
rect 13360 21088 13412 21140
rect 16212 21088 16264 21140
rect 18696 21088 18748 21140
rect 24768 21088 24820 21140
rect 20076 21020 20128 21072
rect 9956 20995 10008 21004
rect 9956 20961 9965 20995
rect 9965 20961 9999 20995
rect 9999 20961 10008 20995
rect 9956 20952 10008 20961
rect 10968 20952 11020 21004
rect 12624 20952 12676 21004
rect 16764 20952 16816 21004
rect 19616 20952 19668 21004
rect 22008 20995 22060 21004
rect 22008 20961 22017 20995
rect 22017 20961 22051 20995
rect 22051 20961 22060 20995
rect 22008 20952 22060 20961
rect 10692 20927 10744 20936
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 25044 21020 25096 21072
rect 24860 20952 24912 21004
rect 24216 20884 24268 20936
rect 25504 20884 25556 20936
rect 8576 20816 8628 20868
rect 10876 20816 10928 20868
rect 8852 20748 8904 20800
rect 15752 20816 15804 20868
rect 14556 20748 14608 20800
rect 15660 20748 15712 20800
rect 19248 20816 19300 20868
rect 24952 20859 25004 20868
rect 24952 20825 24961 20859
rect 24961 20825 24995 20859
rect 24995 20825 25004 20859
rect 24952 20816 25004 20825
rect 25320 20816 25372 20868
rect 17224 20748 17276 20800
rect 17500 20748 17552 20800
rect 18788 20791 18840 20800
rect 18788 20757 18797 20791
rect 18797 20757 18831 20791
rect 18831 20757 18840 20791
rect 18788 20748 18840 20757
rect 21456 20791 21508 20800
rect 21456 20757 21465 20791
rect 21465 20757 21499 20791
rect 21499 20757 21508 20791
rect 21456 20748 21508 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 10140 20544 10192 20596
rect 12532 20544 12584 20596
rect 15936 20544 15988 20596
rect 8300 20476 8352 20528
rect 8576 20476 8628 20528
rect 14556 20476 14608 20528
rect 12440 20408 12492 20460
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 19432 20544 19484 20596
rect 21456 20544 21508 20596
rect 22836 20544 22888 20596
rect 24032 20544 24084 20596
rect 25412 20544 25464 20596
rect 17132 20519 17184 20528
rect 17132 20485 17141 20519
rect 17141 20485 17175 20519
rect 17175 20485 17184 20519
rect 17132 20476 17184 20485
rect 18788 20476 18840 20528
rect 18880 20476 18932 20528
rect 19156 20408 19208 20460
rect 20352 20408 20404 20460
rect 21180 20476 21232 20528
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 7748 20383 7800 20392
rect 7748 20349 7757 20383
rect 7757 20349 7791 20383
rect 7791 20349 7800 20383
rect 7748 20340 7800 20349
rect 8392 20340 8444 20392
rect 9312 20340 9364 20392
rect 9772 20383 9824 20392
rect 9772 20349 9781 20383
rect 9781 20349 9815 20383
rect 9815 20349 9824 20383
rect 9772 20340 9824 20349
rect 10232 20340 10284 20392
rect 13452 20340 13504 20392
rect 15108 20340 15160 20392
rect 17500 20340 17552 20392
rect 18604 20383 18656 20392
rect 18604 20349 18613 20383
rect 18613 20349 18647 20383
rect 18647 20349 18656 20383
rect 18604 20340 18656 20349
rect 22560 20340 22612 20392
rect 23572 20383 23624 20392
rect 23572 20349 23581 20383
rect 23581 20349 23615 20383
rect 23615 20349 23624 20383
rect 23572 20340 23624 20349
rect 25136 20340 25188 20392
rect 10140 20247 10192 20256
rect 10140 20213 10149 20247
rect 10149 20213 10183 20247
rect 10183 20213 10192 20247
rect 10140 20204 10192 20213
rect 14464 20247 14516 20256
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 19156 20272 19208 20324
rect 21548 20272 21600 20324
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19340 20204 19392 20256
rect 22468 20247 22520 20256
rect 22468 20213 22477 20247
rect 22477 20213 22511 20247
rect 22511 20213 22520 20247
rect 22468 20204 22520 20213
rect 23940 20204 23992 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 8576 20000 8628 20052
rect 14188 20000 14240 20052
rect 15568 20000 15620 20052
rect 15752 20000 15804 20052
rect 17224 20000 17276 20052
rect 15844 19932 15896 19984
rect 17040 19932 17092 19984
rect 17132 19932 17184 19984
rect 7748 19796 7800 19848
rect 9036 19796 9088 19848
rect 10692 19864 10744 19916
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 12440 19864 12492 19916
rect 14648 19864 14700 19916
rect 17224 19864 17276 19916
rect 17868 19864 17920 19916
rect 15660 19796 15712 19848
rect 8668 19728 8720 19780
rect 9496 19728 9548 19780
rect 10140 19728 10192 19780
rect 11612 19728 11664 19780
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 12532 19660 12584 19712
rect 22192 20000 22244 20052
rect 23664 20000 23716 20052
rect 24216 20000 24268 20052
rect 25320 20043 25372 20052
rect 25320 20009 25329 20043
rect 25329 20009 25363 20043
rect 25363 20009 25372 20043
rect 25320 20000 25372 20009
rect 21640 19975 21692 19984
rect 21640 19941 21649 19975
rect 21649 19941 21683 19975
rect 21683 19941 21692 19975
rect 21640 19932 21692 19941
rect 20168 19864 20220 19916
rect 19708 19796 19760 19848
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 17040 19728 17092 19780
rect 19800 19728 19852 19780
rect 19892 19728 19944 19780
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 18788 19660 18840 19712
rect 22468 19728 22520 19780
rect 24216 19660 24268 19712
rect 24584 19703 24636 19712
rect 24584 19669 24593 19703
rect 24593 19669 24627 19703
rect 24627 19669 24636 19703
rect 24584 19660 24636 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 10140 19456 10192 19508
rect 11152 19456 11204 19508
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 11796 19456 11848 19508
rect 8576 19388 8628 19440
rect 9220 19388 9272 19440
rect 15476 19456 15528 19508
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 6920 19252 6972 19304
rect 10140 19320 10192 19372
rect 12440 19320 12492 19372
rect 14556 19320 14608 19372
rect 16396 19320 16448 19372
rect 17224 19499 17276 19508
rect 17224 19465 17233 19499
rect 17233 19465 17267 19499
rect 17267 19465 17276 19499
rect 17224 19456 17276 19465
rect 17316 19499 17368 19508
rect 17316 19465 17325 19499
rect 17325 19465 17359 19499
rect 17359 19465 17368 19499
rect 17316 19456 17368 19465
rect 17408 19456 17460 19508
rect 18696 19456 18748 19508
rect 19524 19456 19576 19508
rect 20720 19456 20772 19508
rect 23480 19456 23532 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 22192 19388 22244 19440
rect 8484 19184 8536 19236
rect 14464 19252 14516 19304
rect 9404 19184 9456 19236
rect 10968 19184 11020 19236
rect 15752 19184 15804 19236
rect 17776 19252 17828 19304
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 19892 19320 19944 19372
rect 20352 19320 20404 19372
rect 23572 19388 23624 19440
rect 23664 19431 23716 19440
rect 23664 19397 23673 19431
rect 23673 19397 23707 19431
rect 23707 19397 23716 19431
rect 23664 19388 23716 19397
rect 24216 19388 24268 19440
rect 19984 19252 20036 19304
rect 21640 19252 21692 19304
rect 22744 19295 22796 19304
rect 22744 19261 22753 19295
rect 22753 19261 22787 19295
rect 22787 19261 22796 19295
rect 22744 19252 22796 19261
rect 17592 19184 17644 19236
rect 21180 19184 21232 19236
rect 21456 19184 21508 19236
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 9312 19116 9364 19168
rect 10324 19116 10376 19168
rect 11612 19116 11664 19168
rect 14096 19116 14148 19168
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 15108 19116 15160 19168
rect 18788 19116 18840 19168
rect 21824 19159 21876 19168
rect 21824 19125 21833 19159
rect 21833 19125 21867 19159
rect 21867 19125 21876 19159
rect 21824 19116 21876 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 8576 18912 8628 18964
rect 10048 18955 10100 18964
rect 10048 18921 10057 18955
rect 10057 18921 10091 18955
rect 10091 18921 10100 18955
rect 10048 18912 10100 18921
rect 8300 18776 8352 18828
rect 11244 18912 11296 18964
rect 12532 18912 12584 18964
rect 12716 18955 12768 18964
rect 12716 18921 12725 18955
rect 12725 18921 12759 18955
rect 12759 18921 12768 18955
rect 12716 18912 12768 18921
rect 10968 18844 11020 18896
rect 10876 18776 10928 18828
rect 16672 18776 16724 18828
rect 17592 18912 17644 18964
rect 21640 18844 21692 18896
rect 17592 18776 17644 18828
rect 18604 18776 18656 18828
rect 23388 18776 23440 18828
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 8576 18708 8628 18760
rect 8760 18708 8812 18760
rect 9128 18708 9180 18760
rect 8300 18640 8352 18692
rect 11244 18640 11296 18692
rect 12072 18640 12124 18692
rect 8576 18572 8628 18624
rect 8852 18572 8904 18624
rect 11428 18572 11480 18624
rect 13820 18708 13872 18760
rect 17776 18708 17828 18760
rect 12624 18640 12676 18692
rect 18972 18640 19024 18692
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 24584 18708 24636 18760
rect 24400 18640 24452 18692
rect 24492 18640 24544 18692
rect 24952 18640 25004 18692
rect 12808 18572 12860 18624
rect 13912 18572 13964 18624
rect 14280 18615 14332 18624
rect 14280 18581 14289 18615
rect 14289 18581 14323 18615
rect 14323 18581 14332 18615
rect 14280 18572 14332 18581
rect 17040 18572 17092 18624
rect 18328 18572 18380 18624
rect 19892 18572 19944 18624
rect 22100 18572 22152 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 9404 18368 9456 18420
rect 10784 18368 10836 18420
rect 11152 18368 11204 18420
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 11520 18368 11572 18420
rect 12440 18368 12492 18420
rect 8300 18300 8352 18352
rect 8760 18300 8812 18352
rect 9312 18300 9364 18352
rect 13820 18411 13872 18420
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 16856 18368 16908 18420
rect 26148 18368 26200 18420
rect 6644 18164 6696 18216
rect 8116 18164 8168 18216
rect 18880 18300 18932 18352
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 16764 18232 16816 18284
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 22376 18300 22428 18352
rect 24860 18300 24912 18352
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 13912 18164 13964 18216
rect 9036 18096 9088 18148
rect 9588 18096 9640 18148
rect 11796 18096 11848 18148
rect 9772 18028 9824 18080
rect 13728 18028 13780 18080
rect 17500 18164 17552 18216
rect 24676 18207 24728 18216
rect 24676 18173 24685 18207
rect 24685 18173 24719 18207
rect 24719 18173 24728 18207
rect 24676 18164 24728 18173
rect 16856 18096 16908 18148
rect 25228 18096 25280 18148
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 18880 18071 18932 18080
rect 18880 18037 18889 18071
rect 18889 18037 18923 18071
rect 18923 18037 18932 18071
rect 18880 18028 18932 18037
rect 21088 18071 21140 18080
rect 21088 18037 21097 18071
rect 21097 18037 21131 18071
rect 21131 18037 21140 18071
rect 21088 18028 21140 18037
rect 22744 18028 22796 18080
rect 24124 18028 24176 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 7656 17824 7708 17876
rect 12072 17824 12124 17876
rect 13912 17824 13964 17876
rect 17960 17824 18012 17876
rect 18696 17824 18748 17876
rect 18880 17824 18932 17876
rect 9772 17756 9824 17808
rect 15200 17756 15252 17808
rect 16948 17756 17000 17808
rect 17868 17756 17920 17808
rect 7840 17688 7892 17740
rect 13360 17688 13412 17740
rect 16028 17688 16080 17740
rect 17500 17688 17552 17740
rect 19432 17688 19484 17740
rect 19800 17688 19852 17740
rect 9588 17620 9640 17672
rect 11152 17620 11204 17672
rect 11336 17620 11388 17672
rect 11796 17663 11848 17672
rect 11796 17629 11805 17663
rect 11805 17629 11839 17663
rect 11839 17629 11848 17663
rect 11796 17620 11848 17629
rect 14280 17620 14332 17672
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 17776 17663 17828 17672
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 19708 17620 19760 17672
rect 26056 17824 26108 17876
rect 24860 17688 24912 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 24584 17620 24636 17672
rect 8760 17552 8812 17604
rect 12440 17552 12492 17604
rect 17684 17552 17736 17604
rect 17868 17595 17920 17604
rect 17868 17561 17877 17595
rect 17877 17561 17911 17595
rect 17911 17561 17920 17595
rect 17868 17552 17920 17561
rect 19248 17552 19300 17604
rect 19800 17552 19852 17604
rect 20260 17552 20312 17604
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 8300 17527 8352 17536
rect 8300 17493 8309 17527
rect 8309 17493 8343 17527
rect 8343 17493 8352 17527
rect 8300 17484 8352 17493
rect 9404 17484 9456 17536
rect 12072 17484 12124 17536
rect 13176 17484 13228 17536
rect 15476 17527 15528 17536
rect 15476 17493 15485 17527
rect 15485 17493 15519 17527
rect 15519 17493 15528 17527
rect 15476 17484 15528 17493
rect 15568 17484 15620 17536
rect 15752 17484 15804 17536
rect 16304 17484 16356 17536
rect 17408 17527 17460 17536
rect 17408 17493 17417 17527
rect 17417 17493 17451 17527
rect 17451 17493 17460 17527
rect 17408 17484 17460 17493
rect 22192 17595 22244 17604
rect 22192 17561 22201 17595
rect 22201 17561 22235 17595
rect 22235 17561 22244 17595
rect 22192 17552 22244 17561
rect 25044 17552 25096 17604
rect 22836 17484 22888 17536
rect 24676 17484 24728 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 7196 17280 7248 17332
rect 8392 17280 8444 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11336 17280 11388 17332
rect 12440 17280 12492 17332
rect 13176 17323 13228 17332
rect 13176 17289 13185 17323
rect 13185 17289 13219 17323
rect 13219 17289 13228 17323
rect 13176 17280 13228 17289
rect 9588 17212 9640 17264
rect 7288 17076 7340 17128
rect 8576 17144 8628 17196
rect 8944 17144 8996 17196
rect 11336 17144 11388 17196
rect 12440 17144 12492 17196
rect 12808 17144 12860 17196
rect 16396 17280 16448 17332
rect 16764 17280 16816 17332
rect 20352 17323 20404 17332
rect 20352 17289 20361 17323
rect 20361 17289 20395 17323
rect 20395 17289 20404 17323
rect 20352 17280 20404 17289
rect 22744 17323 22796 17332
rect 22744 17289 22753 17323
rect 22753 17289 22787 17323
rect 22787 17289 22796 17323
rect 22744 17280 22796 17289
rect 16120 17212 16172 17264
rect 17132 17212 17184 17264
rect 18420 17212 18472 17264
rect 23756 17255 23808 17264
rect 23756 17221 23765 17255
rect 23765 17221 23799 17255
rect 23799 17221 23808 17255
rect 23756 17212 23808 17221
rect 24216 17212 24268 17264
rect 19984 17144 20036 17196
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 3332 16940 3384 16992
rect 9404 17076 9456 17128
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 11152 17076 11204 17128
rect 12072 16983 12124 16992
rect 12072 16949 12081 16983
rect 12081 16949 12115 16983
rect 12115 16949 12124 16983
rect 12072 16940 12124 16949
rect 13452 17119 13504 17128
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 15568 17076 15620 17128
rect 16304 17119 16356 17128
rect 16304 17085 16313 17119
rect 16313 17085 16347 17119
rect 16347 17085 16356 17119
rect 16304 17076 16356 17085
rect 17868 17076 17920 17128
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 22836 17076 22888 17128
rect 13636 17008 13688 17060
rect 15936 17008 15988 17060
rect 12716 16940 12768 16992
rect 15384 16940 15436 16992
rect 16304 16940 16356 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 18420 16940 18472 16992
rect 18696 16940 18748 16992
rect 20996 16940 21048 16992
rect 21824 16940 21876 16992
rect 22376 16940 22428 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 11244 16779 11296 16788
rect 11244 16745 11253 16779
rect 11253 16745 11287 16779
rect 11287 16745 11296 16779
rect 11244 16736 11296 16745
rect 2412 16600 2464 16652
rect 8852 16668 8904 16720
rect 8300 16600 8352 16652
rect 9496 16600 9548 16652
rect 11612 16668 11664 16720
rect 11244 16600 11296 16652
rect 11704 16600 11756 16652
rect 12532 16600 12584 16652
rect 12808 16600 12860 16652
rect 14556 16736 14608 16788
rect 13544 16668 13596 16720
rect 15844 16736 15896 16788
rect 16120 16736 16172 16788
rect 18420 16736 18472 16788
rect 19984 16779 20036 16788
rect 19984 16745 19993 16779
rect 19993 16745 20027 16779
rect 20027 16745 20036 16779
rect 19984 16736 20036 16745
rect 20996 16736 21048 16788
rect 22928 16736 22980 16788
rect 24216 16736 24268 16788
rect 24584 16779 24636 16788
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 16212 16600 16264 16652
rect 16396 16600 16448 16652
rect 17868 16668 17920 16720
rect 22560 16668 22612 16720
rect 23572 16668 23624 16720
rect 13452 16532 13504 16584
rect 13636 16532 13688 16584
rect 15660 16532 15712 16584
rect 10416 16464 10468 16516
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 14096 16464 14148 16516
rect 13636 16396 13688 16448
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 17224 16507 17276 16516
rect 17224 16473 17233 16507
rect 17233 16473 17267 16507
rect 17267 16473 17276 16507
rect 17224 16464 17276 16473
rect 17776 16464 17828 16516
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 15476 16396 15528 16448
rect 16212 16439 16264 16448
rect 16212 16405 16221 16439
rect 16221 16405 16255 16439
rect 16255 16405 16264 16439
rect 16212 16396 16264 16405
rect 19432 16396 19484 16448
rect 20168 16532 20220 16584
rect 22560 16532 22612 16584
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 20628 16464 20680 16516
rect 20996 16464 21048 16516
rect 21916 16396 21968 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 8484 16192 8536 16244
rect 8576 16124 8628 16176
rect 9128 16192 9180 16244
rect 9312 16192 9364 16244
rect 11612 16192 11664 16244
rect 13544 16192 13596 16244
rect 15016 16192 15068 16244
rect 15660 16192 15712 16244
rect 17224 16192 17276 16244
rect 21364 16192 21416 16244
rect 11796 16167 11848 16176
rect 11796 16133 11805 16167
rect 11805 16133 11839 16167
rect 11839 16133 11848 16167
rect 11796 16124 11848 16133
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 8392 15988 8444 16040
rect 9588 15988 9640 16040
rect 12164 15963 12216 15972
rect 12164 15929 12173 15963
rect 12173 15929 12207 15963
rect 12207 15929 12216 15963
rect 12164 15920 12216 15929
rect 12256 15920 12308 15972
rect 14004 16124 14056 16176
rect 14096 16124 14148 16176
rect 14280 16056 14332 16108
rect 14740 16056 14792 16108
rect 13820 15988 13872 16040
rect 14464 15988 14516 16040
rect 17224 16099 17276 16108
rect 17224 16065 17233 16099
rect 17233 16065 17267 16099
rect 17267 16065 17276 16099
rect 17224 16056 17276 16065
rect 18512 16056 18564 16108
rect 19800 16124 19852 16176
rect 20168 16124 20220 16176
rect 17776 15988 17828 16040
rect 19432 16056 19484 16108
rect 20812 16056 20864 16108
rect 20536 15988 20588 16040
rect 21916 16056 21968 16108
rect 22284 16124 22336 16176
rect 23296 16192 23348 16244
rect 22928 16124 22980 16176
rect 15476 15920 15528 15972
rect 16672 15920 16724 15972
rect 15384 15852 15436 15904
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 16212 15852 16264 15861
rect 17132 15852 17184 15904
rect 17868 15895 17920 15904
rect 17868 15861 17877 15895
rect 17877 15861 17911 15895
rect 17911 15861 17920 15895
rect 17868 15852 17920 15861
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 21916 15920 21968 15972
rect 24584 15988 24636 16040
rect 23480 15920 23532 15972
rect 22652 15852 22704 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 9220 15648 9272 15700
rect 9312 15648 9364 15700
rect 11060 15648 11112 15700
rect 15476 15691 15528 15700
rect 15476 15657 15485 15691
rect 15485 15657 15519 15691
rect 15519 15657 15528 15691
rect 15476 15648 15528 15657
rect 5172 15580 5224 15632
rect 12072 15580 12124 15632
rect 14280 15580 14332 15632
rect 18696 15648 18748 15700
rect 20720 15648 20772 15700
rect 24400 15648 24452 15700
rect 9588 15512 9640 15564
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12256 15512 12308 15521
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 18604 15512 18656 15564
rect 20168 15512 20220 15564
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 22652 15512 22704 15564
rect 24676 15512 24728 15564
rect 5448 15444 5500 15496
rect 13544 15444 13596 15496
rect 21640 15444 21692 15496
rect 9220 15376 9272 15428
rect 12532 15376 12584 15428
rect 19616 15376 19668 15428
rect 10048 15308 10100 15360
rect 12716 15308 12768 15360
rect 13820 15308 13872 15360
rect 14188 15308 14240 15360
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 17684 15308 17736 15360
rect 18420 15351 18472 15360
rect 18420 15317 18429 15351
rect 18429 15317 18463 15351
rect 18463 15317 18472 15351
rect 18420 15308 18472 15317
rect 20996 15376 21048 15428
rect 21456 15376 21508 15428
rect 22652 15376 22704 15428
rect 20352 15308 20404 15360
rect 20628 15308 20680 15360
rect 21916 15308 21968 15360
rect 23572 15308 23624 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 10140 15147 10192 15156
rect 10140 15113 10149 15147
rect 10149 15113 10183 15147
rect 10183 15113 10192 15147
rect 10140 15104 10192 15113
rect 10232 15104 10284 15156
rect 11336 15147 11388 15156
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 12072 15104 12124 15156
rect 12808 15104 12860 15156
rect 14280 15104 14332 15156
rect 15752 15104 15804 15156
rect 17224 15104 17276 15156
rect 20076 15147 20128 15156
rect 20076 15113 20085 15147
rect 20085 15113 20119 15147
rect 20119 15113 20128 15147
rect 20076 15104 20128 15113
rect 8576 15036 8628 15088
rect 18788 15036 18840 15088
rect 22836 15104 22888 15156
rect 9588 14968 9640 15020
rect 8484 14900 8536 14952
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 11612 14968 11664 15020
rect 11796 14968 11848 15020
rect 14464 14968 14516 15020
rect 15200 14968 15252 15020
rect 18604 14968 18656 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 23204 15036 23256 15088
rect 23296 15079 23348 15088
rect 23296 15045 23305 15079
rect 23305 15045 23339 15079
rect 23339 15045 23348 15079
rect 23296 15036 23348 15045
rect 21456 14968 21508 15020
rect 22008 14968 22060 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 11428 14832 11480 14884
rect 15660 14900 15712 14952
rect 16856 14900 16908 14952
rect 20628 14900 20680 14952
rect 24768 14943 24820 14952
rect 24768 14909 24777 14943
rect 24777 14909 24811 14943
rect 24811 14909 24820 14943
rect 24768 14900 24820 14909
rect 14648 14832 14700 14884
rect 18972 14832 19024 14884
rect 24676 14832 24728 14884
rect 8300 14764 8352 14816
rect 11152 14764 11204 14816
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 12808 14764 12860 14816
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 16948 14764 17000 14816
rect 21456 14764 21508 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 7840 14560 7892 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 8300 14424 8352 14476
rect 8576 14356 8628 14408
rect 9036 14288 9088 14340
rect 9864 14560 9916 14612
rect 11796 14560 11848 14612
rect 12624 14560 12676 14612
rect 15752 14560 15804 14612
rect 16580 14560 16632 14612
rect 20168 14560 20220 14612
rect 9680 14424 9732 14476
rect 11704 14424 11756 14476
rect 12164 14424 12216 14476
rect 14740 14467 14792 14476
rect 9588 14356 9640 14408
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 15568 14492 15620 14544
rect 14924 14424 14976 14476
rect 17592 14492 17644 14544
rect 19340 14492 19392 14544
rect 19708 14492 19760 14544
rect 20444 14492 20496 14544
rect 22468 14492 22520 14544
rect 21548 14424 21600 14476
rect 22100 14467 22152 14476
rect 22100 14433 22109 14467
rect 22109 14433 22143 14467
rect 22143 14433 22152 14467
rect 22100 14424 22152 14433
rect 24860 14424 24912 14476
rect 11152 14220 11204 14272
rect 11244 14220 11296 14272
rect 16580 14356 16632 14408
rect 16672 14356 16724 14408
rect 20260 14356 20312 14408
rect 21824 14356 21876 14408
rect 23940 14356 23992 14408
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 13912 14288 13964 14340
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 13544 14263 13596 14272
rect 13544 14229 13553 14263
rect 13553 14229 13587 14263
rect 13587 14229 13596 14263
rect 13544 14220 13596 14229
rect 14372 14220 14424 14272
rect 19616 14220 19668 14272
rect 19800 14220 19852 14272
rect 21824 14263 21876 14272
rect 21824 14229 21833 14263
rect 21833 14229 21867 14263
rect 21867 14229 21876 14263
rect 21824 14220 21876 14229
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 8300 14016 8352 14068
rect 9588 14016 9640 14068
rect 9772 14016 9824 14068
rect 13544 14016 13596 14068
rect 16672 14016 16724 14068
rect 16764 14016 16816 14068
rect 17316 14016 17368 14068
rect 7932 13948 7984 14000
rect 8576 13948 8628 14000
rect 10232 13991 10284 14000
rect 10232 13957 10241 13991
rect 10241 13957 10275 13991
rect 10275 13957 10284 13991
rect 10232 13948 10284 13957
rect 12440 13948 12492 14000
rect 13820 13948 13872 14000
rect 16120 13948 16172 14000
rect 23388 14016 23440 14068
rect 9588 13880 9640 13932
rect 15660 13880 15712 13932
rect 18420 13948 18472 14000
rect 19524 13991 19576 14000
rect 19524 13957 19533 13991
rect 19533 13957 19567 13991
rect 19567 13957 19576 13991
rect 19524 13948 19576 13957
rect 19708 13948 19760 14000
rect 19616 13880 19668 13932
rect 21364 13880 21416 13932
rect 22652 13948 22704 14000
rect 22836 13948 22888 14000
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 9864 13812 9916 13864
rect 11060 13812 11112 13864
rect 12256 13812 12308 13864
rect 12900 13744 12952 13796
rect 13452 13812 13504 13864
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17500 13812 17552 13864
rect 15844 13744 15896 13796
rect 11888 13676 11940 13728
rect 12164 13676 12216 13728
rect 14096 13719 14148 13728
rect 14096 13685 14126 13719
rect 14126 13685 14148 13719
rect 14096 13676 14148 13685
rect 18880 13812 18932 13864
rect 21640 13812 21692 13864
rect 22560 13812 22612 13864
rect 22652 13812 22704 13864
rect 22284 13744 22336 13796
rect 23204 13812 23256 13864
rect 18972 13719 19024 13728
rect 18972 13685 18981 13719
rect 18981 13685 19015 13719
rect 19015 13685 19024 13719
rect 18972 13676 19024 13685
rect 23572 13676 23624 13728
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 8392 13472 8444 13524
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 8760 13472 8812 13524
rect 13636 13472 13688 13524
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 17316 13472 17368 13524
rect 17960 13472 18012 13524
rect 18420 13472 18472 13524
rect 21088 13472 21140 13524
rect 23940 13472 23992 13524
rect 9036 13404 9088 13456
rect 9312 13404 9364 13456
rect 6460 13336 6512 13388
rect 12900 13404 12952 13456
rect 15292 13404 15344 13456
rect 11704 13336 11756 13388
rect 13452 13379 13504 13388
rect 13452 13345 13461 13379
rect 13461 13345 13495 13379
rect 13495 13345 13504 13379
rect 13452 13336 13504 13345
rect 13544 13336 13596 13388
rect 15200 13336 15252 13388
rect 15476 13336 15528 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 16120 13336 16172 13388
rect 21456 13404 21508 13456
rect 12440 13268 12492 13320
rect 8576 13200 8628 13252
rect 9128 13200 9180 13252
rect 9036 13132 9088 13184
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 11152 13200 11204 13252
rect 17316 13268 17368 13320
rect 17500 13268 17552 13320
rect 20720 13336 20772 13388
rect 17960 13268 18012 13320
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 25044 13336 25096 13388
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 12072 13132 12124 13184
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 14740 13132 14792 13184
rect 15384 13132 15436 13184
rect 17132 13132 17184 13184
rect 20260 13243 20312 13252
rect 20260 13209 20269 13243
rect 20269 13209 20303 13243
rect 20303 13209 20312 13243
rect 20260 13200 20312 13209
rect 18696 13132 18748 13184
rect 21272 13200 21324 13252
rect 23388 13200 23440 13252
rect 20996 13132 21048 13184
rect 22376 13132 22428 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 7748 12928 7800 12980
rect 9220 12928 9272 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 9772 12928 9824 12980
rect 10048 12928 10100 12980
rect 11060 12928 11112 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 12532 12928 12584 12980
rect 13452 12928 13504 12980
rect 14924 12928 14976 12980
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 6920 12860 6972 12912
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7104 12767 7156 12776
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 7656 12860 7708 12912
rect 12348 12860 12400 12912
rect 15568 12860 15620 12912
rect 17408 12928 17460 12980
rect 17776 12928 17828 12980
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 21272 12928 21324 12980
rect 21456 12928 21508 12980
rect 22008 12971 22060 12980
rect 22008 12937 22017 12971
rect 22017 12937 22051 12971
rect 22051 12937 22060 12971
rect 22008 12928 22060 12937
rect 22836 12971 22888 12980
rect 22836 12937 22845 12971
rect 22845 12937 22879 12971
rect 22879 12937 22888 12971
rect 22836 12928 22888 12937
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 7840 12724 7892 12776
rect 8668 12724 8720 12776
rect 9036 12724 9088 12776
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 11888 12792 11940 12844
rect 12532 12724 12584 12776
rect 12900 12724 12952 12776
rect 13636 12792 13688 12844
rect 14556 12792 14608 12844
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 18328 12792 18380 12844
rect 18512 12860 18564 12912
rect 14096 12724 14148 12776
rect 15200 12724 15252 12776
rect 15844 12724 15896 12776
rect 18880 12724 18932 12776
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 20904 12860 20956 12912
rect 20996 12792 21048 12844
rect 22100 12860 22152 12912
rect 23296 12860 23348 12912
rect 20536 12724 20588 12776
rect 22008 12792 22060 12844
rect 11152 12656 11204 12708
rect 11336 12588 11388 12640
rect 11796 12656 11848 12708
rect 19708 12656 19760 12708
rect 12348 12588 12400 12640
rect 14740 12588 14792 12640
rect 15476 12588 15528 12640
rect 17316 12588 17368 12640
rect 18696 12588 18748 12640
rect 20812 12656 20864 12708
rect 22652 12724 22704 12776
rect 22560 12656 22612 12708
rect 22376 12588 22428 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 9496 12384 9548 12436
rect 10508 12384 10560 12436
rect 11888 12384 11940 12436
rect 12164 12384 12216 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 13820 12384 13872 12436
rect 17316 12384 17368 12436
rect 18788 12384 18840 12436
rect 20076 12384 20128 12436
rect 20168 12384 20220 12436
rect 21732 12384 21784 12436
rect 24124 12384 24176 12436
rect 11060 12316 11112 12368
rect 7012 12248 7064 12300
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 9036 12248 9088 12300
rect 9312 12248 9364 12300
rect 14004 12316 14056 12368
rect 14556 12316 14608 12368
rect 19248 12316 19300 12368
rect 22836 12316 22888 12368
rect 7472 12180 7524 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12164 12248 12216 12300
rect 13728 12248 13780 12300
rect 14924 12248 14976 12300
rect 15844 12248 15896 12300
rect 19156 12248 19208 12300
rect 11520 12112 11572 12164
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 18788 12180 18840 12232
rect 20260 12248 20312 12300
rect 20168 12180 20220 12232
rect 22008 12248 22060 12300
rect 23296 12248 23348 12300
rect 22836 12223 22888 12232
rect 22836 12189 22845 12223
rect 22845 12189 22879 12223
rect 22879 12189 22888 12223
rect 22836 12180 22888 12189
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 13636 12112 13688 12164
rect 8484 12044 8536 12096
rect 9404 12044 9456 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11428 12044 11480 12096
rect 12348 12044 12400 12096
rect 16488 12112 16540 12164
rect 16856 12112 16908 12164
rect 14004 12044 14056 12096
rect 14556 12044 14608 12096
rect 15292 12044 15344 12096
rect 16304 12044 16356 12096
rect 18420 12044 18472 12096
rect 18696 12112 18748 12164
rect 19432 12112 19484 12164
rect 20720 12155 20772 12164
rect 20720 12121 20729 12155
rect 20729 12121 20763 12155
rect 20763 12121 20772 12155
rect 20720 12112 20772 12121
rect 24952 12112 25004 12164
rect 18880 12044 18932 12096
rect 19248 12044 19300 12096
rect 19800 12044 19852 12096
rect 20352 12044 20404 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 5356 11840 5408 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9680 11840 9732 11892
rect 10232 11815 10284 11824
rect 10232 11781 10241 11815
rect 10241 11781 10275 11815
rect 10275 11781 10284 11815
rect 10232 11772 10284 11781
rect 12716 11840 12768 11892
rect 13544 11840 13596 11892
rect 14188 11840 14240 11892
rect 16948 11840 17000 11892
rect 17040 11840 17092 11892
rect 9128 11704 9180 11756
rect 9404 11704 9456 11756
rect 11060 11636 11112 11688
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12808 11772 12860 11824
rect 14372 11772 14424 11824
rect 15016 11772 15068 11824
rect 15200 11772 15252 11824
rect 17684 11772 17736 11824
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 22008 11840 22060 11892
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 12624 11636 12676 11688
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 12348 11568 12400 11620
rect 12716 11568 12768 11620
rect 19984 11772 20036 11824
rect 20076 11815 20128 11824
rect 20076 11781 20085 11815
rect 20085 11781 20119 11815
rect 20119 11781 20128 11815
rect 20076 11772 20128 11781
rect 20628 11772 20680 11824
rect 21732 11772 21784 11824
rect 24860 11772 24912 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 20536 11704 20588 11756
rect 23940 11704 23992 11756
rect 24952 11704 25004 11756
rect 16028 11636 16080 11688
rect 16672 11636 16724 11688
rect 17776 11636 17828 11688
rect 19800 11636 19852 11688
rect 19984 11636 20036 11688
rect 20904 11636 20956 11688
rect 24216 11636 24268 11688
rect 20168 11568 20220 11620
rect 20352 11568 20404 11620
rect 22284 11568 22336 11620
rect 8300 11500 8352 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10140 11500 10192 11552
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 15016 11500 15068 11552
rect 15476 11500 15528 11552
rect 15660 11500 15712 11552
rect 16028 11500 16080 11552
rect 19340 11500 19392 11552
rect 19800 11500 19852 11552
rect 20628 11500 20680 11552
rect 22008 11500 22060 11552
rect 25780 11500 25832 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 7196 11296 7248 11348
rect 10600 11296 10652 11348
rect 11244 11228 11296 11280
rect 12808 11228 12860 11280
rect 12900 11228 12952 11280
rect 13544 11228 13596 11280
rect 11888 11160 11940 11212
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 11060 11092 11112 11144
rect 13636 11160 13688 11212
rect 15384 11296 15436 11348
rect 15660 11296 15712 11348
rect 16672 11271 16724 11280
rect 16672 11237 16681 11271
rect 16681 11237 16715 11271
rect 16715 11237 16724 11271
rect 16672 11228 16724 11237
rect 16948 11160 17000 11212
rect 17776 11203 17828 11212
rect 17776 11169 17785 11203
rect 17785 11169 17819 11203
rect 17819 11169 17828 11203
rect 17776 11160 17828 11169
rect 16764 11092 16816 11144
rect 4160 11024 4212 11076
rect 7104 11024 7156 11076
rect 10140 11024 10192 11076
rect 12900 11024 12952 11076
rect 15108 11024 15160 11076
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 16488 11024 16540 11076
rect 9680 10956 9732 11008
rect 10876 10999 10928 11008
rect 10876 10965 10885 10999
rect 10885 10965 10919 10999
rect 10919 10965 10928 10999
rect 10876 10956 10928 10965
rect 11244 10956 11296 11008
rect 12256 10956 12308 11008
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 14372 10956 14424 11008
rect 17868 10956 17920 11008
rect 20168 11296 20220 11348
rect 20628 11296 20680 11348
rect 22468 11296 22520 11348
rect 22836 11296 22888 11348
rect 19524 11228 19576 11280
rect 21824 11228 21876 11280
rect 22008 11228 22060 11280
rect 22284 11271 22336 11280
rect 22284 11237 22293 11271
rect 22293 11237 22327 11271
rect 22327 11237 22336 11271
rect 22284 11228 22336 11237
rect 25596 11228 25648 11280
rect 19432 11160 19484 11212
rect 19156 11092 19208 11144
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 20996 11160 21048 11212
rect 21916 11160 21968 11212
rect 20628 11092 20680 11144
rect 23296 11092 23348 11144
rect 19984 10956 20036 11008
rect 20352 11024 20404 11076
rect 21272 11024 21324 11076
rect 22284 11024 22336 11076
rect 23388 11024 23440 11076
rect 21456 10956 21508 11008
rect 24032 10956 24084 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 12164 10752 12216 10804
rect 7104 10412 7156 10464
rect 8208 10684 8260 10736
rect 10140 10616 10192 10668
rect 12808 10795 12860 10804
rect 12808 10761 12817 10795
rect 12817 10761 12851 10795
rect 12851 10761 12860 10795
rect 12808 10752 12860 10761
rect 13912 10752 13964 10804
rect 14372 10752 14424 10804
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 16764 10752 16816 10804
rect 14280 10684 14332 10736
rect 14832 10684 14884 10736
rect 8300 10412 8352 10464
rect 9128 10412 9180 10464
rect 9588 10412 9640 10464
rect 12808 10548 12860 10600
rect 10876 10480 10928 10532
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 15384 10548 15436 10600
rect 16488 10548 16540 10600
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17592 10727 17644 10736
rect 17592 10693 17601 10727
rect 17601 10693 17635 10727
rect 17635 10693 17644 10727
rect 17592 10684 17644 10693
rect 22008 10752 22060 10804
rect 23204 10752 23256 10804
rect 19524 10684 19576 10736
rect 20076 10684 20128 10736
rect 21088 10727 21140 10736
rect 21088 10693 21097 10727
rect 21097 10693 21131 10727
rect 21131 10693 21140 10727
rect 21088 10684 21140 10693
rect 21180 10727 21232 10736
rect 21180 10693 21189 10727
rect 21189 10693 21223 10727
rect 21223 10693 21232 10727
rect 21180 10684 21232 10693
rect 22560 10684 22612 10736
rect 23848 10684 23900 10736
rect 18328 10548 18380 10600
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12440 10412 12492 10464
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 15384 10412 15436 10464
rect 18788 10480 18840 10532
rect 19340 10548 19392 10600
rect 20168 10591 20220 10600
rect 20168 10557 20177 10591
rect 20177 10557 20211 10591
rect 20211 10557 20220 10591
rect 20168 10548 20220 10557
rect 20720 10548 20772 10600
rect 21272 10591 21324 10600
rect 21272 10557 21281 10591
rect 21281 10557 21315 10591
rect 21315 10557 21324 10591
rect 21272 10548 21324 10557
rect 22652 10616 22704 10668
rect 22744 10548 22796 10600
rect 17316 10412 17368 10464
rect 18420 10412 18472 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 21364 10480 21416 10532
rect 23388 10412 23440 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 8208 10208 8260 10260
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 12072 10208 12124 10260
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 14924 10208 14976 10260
rect 20444 10208 20496 10260
rect 21272 10208 21324 10260
rect 9588 10072 9640 10124
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12440 10140 12492 10192
rect 17040 10140 17092 10192
rect 17868 10140 17920 10192
rect 20352 10140 20404 10192
rect 21824 10140 21876 10192
rect 24308 10208 24360 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 22560 10140 22612 10192
rect 23848 10183 23900 10192
rect 23848 10149 23857 10183
rect 23857 10149 23891 10183
rect 23891 10149 23900 10183
rect 23848 10140 23900 10149
rect 24124 10140 24176 10192
rect 12808 10004 12860 10056
rect 13636 10072 13688 10124
rect 14464 10072 14516 10124
rect 15844 10072 15896 10124
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 17776 10072 17828 10124
rect 17960 10072 18012 10124
rect 18328 10072 18380 10124
rect 18788 10072 18840 10124
rect 19524 10072 19576 10124
rect 9496 9936 9548 9988
rect 10968 9936 11020 9988
rect 11520 9936 11572 9988
rect 13912 9936 13964 9988
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 13360 9868 13412 9920
rect 13544 9868 13596 9920
rect 14740 9868 14792 9920
rect 16120 9979 16172 9988
rect 16120 9945 16129 9979
rect 16129 9945 16163 9979
rect 16163 9945 16172 9979
rect 16120 9936 16172 9945
rect 16856 9979 16908 9988
rect 16856 9945 16865 9979
rect 16865 9945 16899 9979
rect 16899 9945 16908 9979
rect 16856 9936 16908 9945
rect 16764 9868 16816 9920
rect 18236 9868 18288 9920
rect 18880 10004 18932 10056
rect 22376 10072 22428 10124
rect 23388 10115 23440 10124
rect 23388 10081 23397 10115
rect 23397 10081 23431 10115
rect 23431 10081 23440 10115
rect 23388 10072 23440 10081
rect 19892 9936 19944 9988
rect 20720 9936 20772 9988
rect 22560 9936 22612 9988
rect 22744 10004 22796 10056
rect 24676 10004 24728 10056
rect 18696 9868 18748 9920
rect 19156 9868 19208 9920
rect 19340 9868 19392 9920
rect 19984 9911 20036 9920
rect 19984 9877 19993 9911
rect 19993 9877 20027 9911
rect 20027 9877 20036 9911
rect 19984 9868 20036 9877
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 20444 9868 20496 9920
rect 21824 9868 21876 9920
rect 22100 9868 22152 9920
rect 24676 9868 24728 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 11520 9596 11572 9648
rect 13452 9664 13504 9716
rect 13912 9707 13964 9716
rect 13912 9673 13921 9707
rect 13921 9673 13955 9707
rect 13955 9673 13964 9707
rect 13912 9664 13964 9673
rect 14556 9664 14608 9716
rect 17868 9664 17920 9716
rect 18512 9664 18564 9716
rect 15292 9596 15344 9648
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 14004 9528 14056 9580
rect 18972 9664 19024 9716
rect 19248 9596 19300 9648
rect 12716 9460 12768 9512
rect 14096 9460 14148 9512
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 15108 9435 15160 9444
rect 15108 9401 15117 9435
rect 15117 9401 15151 9435
rect 15151 9401 15160 9435
rect 15108 9392 15160 9401
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 13820 9324 13872 9376
rect 15384 9324 15436 9376
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 16948 9460 17000 9512
rect 18236 9460 18288 9512
rect 18880 9460 18932 9512
rect 19524 9664 19576 9716
rect 20168 9664 20220 9716
rect 21088 9664 21140 9716
rect 21824 9664 21876 9716
rect 22008 9664 22060 9716
rect 22284 9664 22336 9716
rect 20076 9571 20128 9580
rect 20076 9537 20085 9571
rect 20085 9537 20119 9571
rect 20119 9537 20128 9571
rect 20076 9528 20128 9537
rect 20168 9392 20220 9444
rect 20720 9460 20772 9512
rect 21180 9460 21232 9512
rect 21824 9460 21876 9512
rect 21916 9460 21968 9512
rect 22100 9460 22152 9512
rect 22652 9503 22704 9512
rect 22652 9469 22661 9503
rect 22661 9469 22695 9503
rect 22695 9469 22704 9503
rect 22652 9460 22704 9469
rect 23388 9460 23440 9512
rect 24400 9528 24452 9580
rect 24124 9460 24176 9512
rect 18696 9324 18748 9376
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 19248 9324 19300 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 19892 9324 19944 9376
rect 21640 9324 21692 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 12072 9120 12124 9172
rect 15016 9120 15068 9172
rect 19064 9120 19116 9172
rect 10692 9052 10744 9104
rect 13728 9052 13780 9104
rect 11060 8984 11112 9036
rect 11704 8984 11756 9036
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 14464 8984 14516 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 15844 8916 15896 8968
rect 19432 9052 19484 9104
rect 21180 9120 21232 9172
rect 22836 9120 22888 9172
rect 23296 9120 23348 9172
rect 23940 9120 23992 9172
rect 21548 9052 21600 9104
rect 18236 8984 18288 9036
rect 19248 8984 19300 9036
rect 20260 8984 20312 9036
rect 20352 8984 20404 9036
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 9680 8848 9732 8900
rect 11336 8848 11388 8900
rect 12532 8848 12584 8900
rect 12900 8848 12952 8900
rect 14004 8848 14056 8900
rect 14924 8848 14976 8900
rect 15384 8848 15436 8900
rect 15568 8848 15620 8900
rect 10968 8780 11020 8832
rect 14464 8780 14516 8832
rect 14556 8780 14608 8832
rect 15108 8780 15160 8832
rect 19524 8916 19576 8968
rect 22560 8916 22612 8968
rect 19432 8848 19484 8900
rect 21640 8848 21692 8900
rect 22468 8848 22520 8900
rect 24952 8848 25004 8900
rect 21180 8780 21232 8832
rect 21732 8780 21784 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 9864 8576 9916 8628
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 13820 8508 13872 8560
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 11612 8440 11664 8492
rect 15016 8440 15068 8492
rect 15752 8508 15804 8560
rect 17592 8508 17644 8560
rect 18696 8508 18748 8560
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 13360 8372 13412 8424
rect 3792 8304 3844 8356
rect 4804 8304 4856 8356
rect 5264 8304 5316 8356
rect 11152 8304 11204 8356
rect 12532 8304 12584 8356
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 14004 8304 14056 8356
rect 14648 8304 14700 8356
rect 17592 8415 17644 8424
rect 17592 8381 17601 8415
rect 17601 8381 17635 8415
rect 17635 8381 17644 8415
rect 17592 8372 17644 8381
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 19708 8440 19760 8492
rect 18512 8372 18564 8424
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 19984 8304 20036 8356
rect 22836 8508 22888 8560
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22468 8372 22520 8424
rect 24584 8372 24636 8424
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 23848 8304 23900 8356
rect 17592 8236 17644 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 11980 8032 12032 8084
rect 12716 8032 12768 8084
rect 13728 8032 13780 8084
rect 14832 8032 14884 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 17868 8032 17920 8084
rect 19156 8032 19208 8084
rect 20720 8032 20772 8084
rect 8392 7964 8444 8016
rect 11612 7939 11664 7948
rect 11612 7905 11621 7939
rect 11621 7905 11655 7939
rect 11655 7905 11664 7939
rect 11612 7896 11664 7905
rect 11888 7896 11940 7948
rect 15200 7964 15252 8016
rect 13728 7896 13780 7948
rect 14924 7896 14976 7948
rect 15476 7896 15528 7948
rect 15752 7896 15804 7948
rect 11704 7828 11756 7880
rect 12440 7828 12492 7880
rect 12624 7828 12676 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 16120 7828 16172 7880
rect 21272 7896 21324 7948
rect 21916 7896 21968 7948
rect 22100 7939 22152 7948
rect 22100 7905 22109 7939
rect 22109 7905 22143 7939
rect 22143 7905 22152 7939
rect 22100 7896 22152 7905
rect 23388 8032 23440 8084
rect 23940 7964 23992 8016
rect 18604 7828 18656 7880
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 20628 7828 20680 7880
rect 12808 7760 12860 7812
rect 11612 7692 11664 7744
rect 12624 7692 12676 7744
rect 12900 7692 12952 7744
rect 14280 7692 14332 7744
rect 17224 7760 17276 7812
rect 15476 7692 15528 7744
rect 15660 7692 15712 7744
rect 16028 7692 16080 7744
rect 16856 7735 16908 7744
rect 16856 7701 16865 7735
rect 16865 7701 16899 7735
rect 16899 7701 16908 7735
rect 16856 7692 16908 7701
rect 19708 7803 19760 7812
rect 19708 7769 19717 7803
rect 19717 7769 19751 7803
rect 19751 7769 19760 7803
rect 19708 7760 19760 7769
rect 21456 7803 21508 7812
rect 21456 7769 21465 7803
rect 21465 7769 21499 7803
rect 21499 7769 21508 7803
rect 21456 7760 21508 7769
rect 24124 7828 24176 7880
rect 21364 7692 21416 7744
rect 22376 7803 22428 7812
rect 22376 7769 22385 7803
rect 22385 7769 22419 7803
rect 22419 7769 22428 7803
rect 22376 7760 22428 7769
rect 23756 7692 23808 7744
rect 24124 7735 24176 7744
rect 24124 7701 24133 7735
rect 24133 7701 24167 7735
rect 24167 7701 24176 7735
rect 24124 7692 24176 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 9128 7488 9180 7540
rect 9588 7420 9640 7472
rect 11336 7488 11388 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12348 7488 12400 7540
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 13636 7488 13688 7540
rect 17224 7531 17276 7540
rect 17224 7497 17233 7531
rect 17233 7497 17267 7531
rect 17267 7497 17276 7531
rect 17224 7488 17276 7497
rect 17408 7488 17460 7540
rect 17868 7488 17920 7540
rect 14280 7420 14332 7472
rect 14740 7420 14792 7472
rect 16580 7420 16632 7472
rect 16856 7420 16908 7472
rect 11336 7352 11388 7404
rect 11520 7352 11572 7404
rect 19616 7488 19668 7540
rect 20260 7488 20312 7540
rect 21916 7488 21968 7540
rect 22928 7488 22980 7540
rect 23388 7488 23440 7540
rect 24860 7420 24912 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 19892 7352 19944 7404
rect 20352 7352 20404 7404
rect 20444 7352 20496 7404
rect 23480 7352 23532 7404
rect 23940 7395 23992 7404
rect 23940 7361 23949 7395
rect 23949 7361 23983 7395
rect 23983 7361 23992 7395
rect 23940 7352 23992 7361
rect 10968 7284 11020 7336
rect 11152 7284 11204 7336
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 16672 7284 16724 7336
rect 17684 7284 17736 7336
rect 18880 7284 18932 7336
rect 19248 7284 19300 7336
rect 20720 7284 20772 7336
rect 16396 7216 16448 7268
rect 16488 7216 16540 7268
rect 18420 7216 18472 7268
rect 15108 7148 15160 7200
rect 17776 7148 17828 7200
rect 18512 7148 18564 7200
rect 18788 7191 18840 7200
rect 18788 7157 18818 7191
rect 18818 7157 18840 7191
rect 18788 7148 18840 7157
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 21088 7216 21140 7268
rect 21364 7284 21416 7336
rect 24768 7216 24820 7268
rect 21364 7148 21416 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 11520 6944 11572 6996
rect 13912 6944 13964 6996
rect 14740 6944 14792 6996
rect 15660 6944 15712 6996
rect 16028 6944 16080 6996
rect 20444 6944 20496 6996
rect 21456 6944 21508 6996
rect 22560 6944 22612 6996
rect 12900 6876 12952 6928
rect 16488 6876 16540 6928
rect 19524 6876 19576 6928
rect 19892 6876 19944 6928
rect 21272 6876 21324 6928
rect 22652 6876 22704 6928
rect 23664 6876 23716 6928
rect 11060 6808 11112 6860
rect 12716 6808 12768 6860
rect 14372 6851 14424 6860
rect 14372 6817 14381 6851
rect 14381 6817 14415 6851
rect 14415 6817 14424 6851
rect 14372 6808 14424 6817
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 16580 6808 16632 6860
rect 20352 6808 20404 6860
rect 22376 6808 22428 6860
rect 16304 6740 16356 6792
rect 16948 6740 17000 6792
rect 18788 6740 18840 6792
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 20904 6740 20956 6792
rect 11336 6672 11388 6724
rect 11520 6672 11572 6724
rect 12624 6672 12676 6724
rect 4068 6604 4120 6656
rect 7564 6604 7616 6656
rect 13452 6604 13504 6656
rect 16488 6715 16540 6724
rect 16488 6681 16497 6715
rect 16497 6681 16531 6715
rect 16531 6681 16540 6715
rect 16488 6672 16540 6681
rect 17684 6672 17736 6724
rect 17868 6672 17920 6724
rect 14740 6604 14792 6656
rect 23940 6740 23992 6792
rect 24860 6672 24912 6724
rect 19340 6604 19392 6656
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 19800 6647 19852 6656
rect 19800 6613 19809 6647
rect 19809 6613 19843 6647
rect 19843 6613 19852 6647
rect 19800 6604 19852 6613
rect 21088 6604 21140 6656
rect 23756 6604 23808 6656
rect 24492 6604 24544 6656
rect 24676 6604 24728 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 11152 6400 11204 6452
rect 12808 6400 12860 6452
rect 19340 6400 19392 6452
rect 20260 6400 20312 6452
rect 12716 6375 12768 6384
rect 12716 6341 12725 6375
rect 12725 6341 12759 6375
rect 12759 6341 12768 6375
rect 12716 6332 12768 6341
rect 13636 6332 13688 6384
rect 6552 6264 6604 6316
rect 11152 6264 11204 6316
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 11336 6196 11388 6248
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 4252 6060 4304 6112
rect 7840 6060 7892 6112
rect 9680 6060 9732 6112
rect 13452 6196 13504 6248
rect 14004 6332 14056 6384
rect 15384 6264 15436 6316
rect 16672 6264 16724 6316
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 16304 6196 16356 6248
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 17960 6307 18012 6316
rect 17960 6273 17969 6307
rect 17969 6273 18003 6307
rect 18003 6273 18012 6307
rect 17960 6264 18012 6273
rect 13728 6128 13780 6180
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 17868 6196 17920 6248
rect 20904 6332 20956 6384
rect 21272 6332 21324 6384
rect 21732 6332 21784 6384
rect 23664 6400 23716 6452
rect 23756 6443 23808 6452
rect 23756 6409 23765 6443
rect 23765 6409 23799 6443
rect 23799 6409 23808 6443
rect 23756 6400 23808 6409
rect 24124 6332 24176 6384
rect 24308 6375 24360 6384
rect 24308 6341 24317 6375
rect 24317 6341 24351 6375
rect 24351 6341 24360 6375
rect 24308 6332 24360 6341
rect 20352 6264 20404 6316
rect 21916 6264 21968 6316
rect 24676 6264 24728 6316
rect 20628 6196 20680 6248
rect 21732 6196 21784 6248
rect 23020 6196 23072 6248
rect 16488 6060 16540 6112
rect 21456 6060 21508 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 11336 5856 11388 5908
rect 14004 5856 14056 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 13728 5788 13780 5840
rect 10784 5720 10836 5772
rect 9588 5652 9640 5704
rect 11520 5720 11572 5772
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 17776 5856 17828 5908
rect 19800 5788 19852 5840
rect 15384 5763 15436 5772
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 13544 5652 13596 5704
rect 15108 5652 15160 5704
rect 16948 5720 17000 5772
rect 18328 5720 18380 5772
rect 18880 5720 18932 5772
rect 19156 5720 19208 5772
rect 20260 5856 20312 5908
rect 20444 5788 20496 5840
rect 24124 5899 24176 5908
rect 24124 5865 24133 5899
rect 24133 5865 24167 5899
rect 24167 5865 24176 5899
rect 24124 5856 24176 5865
rect 24308 5856 24360 5908
rect 24952 5788 25004 5840
rect 20996 5652 21048 5704
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 24584 5652 24636 5704
rect 10416 5516 10468 5568
rect 15200 5627 15252 5636
rect 15200 5593 15209 5627
rect 15209 5593 15243 5627
rect 15243 5593 15252 5627
rect 15200 5584 15252 5593
rect 16488 5584 16540 5636
rect 16672 5584 16724 5636
rect 19248 5584 19300 5636
rect 20628 5584 20680 5636
rect 23388 5584 23440 5636
rect 23480 5627 23532 5636
rect 23480 5593 23489 5627
rect 23489 5593 23523 5627
rect 23523 5593 23532 5627
rect 23480 5584 23532 5593
rect 12440 5516 12492 5568
rect 18328 5516 18380 5568
rect 19340 5516 19392 5568
rect 21916 5516 21968 5568
rect 23112 5559 23164 5568
rect 23112 5525 23121 5559
rect 23121 5525 23155 5559
rect 23155 5525 23164 5559
rect 23112 5516 23164 5525
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 13636 5312 13688 5364
rect 14280 5312 14332 5364
rect 17408 5312 17460 5364
rect 18880 5312 18932 5364
rect 13360 5244 13412 5296
rect 13912 5244 13964 5296
rect 14740 5244 14792 5296
rect 19432 5244 19484 5296
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 21548 5312 21600 5364
rect 21916 5312 21968 5364
rect 11060 5176 11112 5228
rect 11428 5108 11480 5160
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 13084 5176 13136 5228
rect 15844 5176 15896 5228
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 6092 5015 6144 5024
rect 6092 4981 6101 5015
rect 6101 4981 6135 5015
rect 6135 4981 6144 5015
rect 6092 4972 6144 4981
rect 6460 4972 6512 5024
rect 11520 4972 11572 5024
rect 14004 5108 14056 5160
rect 15660 5108 15712 5160
rect 17776 5176 17828 5228
rect 13912 4972 13964 5024
rect 14188 4972 14240 5024
rect 19340 5040 19392 5092
rect 16672 4972 16724 5024
rect 18880 4972 18932 5024
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 22192 5219 22244 5228
rect 22192 5185 22201 5219
rect 22201 5185 22235 5219
rect 22235 5185 22244 5219
rect 22192 5176 22244 5185
rect 21272 5108 21324 5160
rect 21364 5108 21416 5160
rect 25044 5176 25096 5228
rect 19616 5040 19668 5092
rect 20904 5040 20956 5092
rect 22100 4972 22152 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 12072 4768 12124 4820
rect 14188 4768 14240 4820
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 9588 4632 9640 4684
rect 12808 4700 12860 4752
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 11244 4632 11296 4684
rect 14004 4632 14056 4684
rect 17224 4768 17276 4820
rect 18880 4768 18932 4820
rect 16580 4700 16632 4752
rect 19800 4768 19852 4820
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 24400 4768 24452 4820
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 15384 4675 15436 4684
rect 15384 4641 15393 4675
rect 15393 4641 15427 4675
rect 15427 4641 15436 4675
rect 15384 4632 15436 4641
rect 19524 4675 19576 4684
rect 19524 4641 19533 4675
rect 19533 4641 19567 4675
rect 19567 4641 19576 4675
rect 19524 4632 19576 4641
rect 6460 4564 6512 4616
rect 6644 4564 6696 4616
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 12624 4564 12676 4616
rect 14188 4607 14240 4616
rect 14188 4573 14197 4607
rect 14197 4573 14231 4607
rect 14231 4573 14240 4607
rect 14188 4564 14240 4573
rect 14924 4564 14976 4616
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 13176 4496 13228 4548
rect 13268 4539 13320 4548
rect 13268 4505 13277 4539
rect 13277 4505 13311 4539
rect 13311 4505 13320 4539
rect 13268 4496 13320 4505
rect 7380 4428 7432 4480
rect 7748 4471 7800 4480
rect 7748 4437 7757 4471
rect 7757 4437 7791 4471
rect 7791 4437 7800 4471
rect 7748 4428 7800 4437
rect 7840 4428 7892 4480
rect 8300 4471 8352 4480
rect 8300 4437 8309 4471
rect 8309 4437 8343 4471
rect 8343 4437 8352 4471
rect 8300 4428 8352 4437
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 8760 4428 8812 4437
rect 12440 4428 12492 4480
rect 15660 4496 15712 4548
rect 15844 4496 15896 4548
rect 19524 4496 19576 4548
rect 22008 4564 22060 4616
rect 13452 4428 13504 4480
rect 17868 4428 17920 4480
rect 21548 4496 21600 4548
rect 21088 4428 21140 4480
rect 21916 4428 21968 4480
rect 23664 4539 23716 4548
rect 23664 4505 23673 4539
rect 23673 4505 23707 4539
rect 23707 4505 23716 4539
rect 23664 4496 23716 4505
rect 24308 4496 24360 4548
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 7196 4267 7248 4276
rect 7196 4233 7205 4267
rect 7205 4233 7239 4267
rect 7239 4233 7248 4267
rect 7196 4224 7248 4233
rect 10048 4224 10100 4276
rect 1492 4088 1544 4140
rect 2780 4020 2832 4072
rect 4068 4088 4120 4140
rect 5908 4088 5960 4140
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 7012 4088 7064 4140
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 7564 4088 7616 4140
rect 8300 4088 8352 4140
rect 9220 4088 9272 4140
rect 3700 4020 3752 4072
rect 2504 3884 2556 3936
rect 2780 3884 2832 3936
rect 4160 3995 4212 4004
rect 4160 3961 4169 3995
rect 4169 3961 4203 3995
rect 4203 3961 4212 3995
rect 4160 3952 4212 3961
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 4068 3884 4120 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 6552 3995 6604 4004
rect 6552 3961 6561 3995
rect 6561 3961 6595 3995
rect 6595 3961 6604 3995
rect 6552 3952 6604 3961
rect 9680 4020 9732 4072
rect 9956 4020 10008 4072
rect 10048 4020 10100 4072
rect 11336 4224 11388 4276
rect 13268 4224 13320 4276
rect 13176 4156 13228 4208
rect 13820 4156 13872 4208
rect 14280 4156 14332 4208
rect 21548 4267 21600 4276
rect 21548 4233 21557 4267
rect 21557 4233 21591 4267
rect 21591 4233 21600 4267
rect 21548 4224 21600 4233
rect 21640 4224 21692 4276
rect 22008 4224 22060 4276
rect 22100 4267 22152 4276
rect 22100 4233 22109 4267
rect 22109 4233 22143 4267
rect 22143 4233 22152 4267
rect 22100 4224 22152 4233
rect 22744 4267 22796 4276
rect 22744 4233 22753 4267
rect 22753 4233 22787 4267
rect 22787 4233 22796 4267
rect 22744 4224 22796 4233
rect 11428 4088 11480 4140
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 15844 4088 15896 4140
rect 16396 4088 16448 4140
rect 17592 4088 17644 4140
rect 20168 4156 20220 4208
rect 21916 4156 21968 4208
rect 23296 4156 23348 4208
rect 18512 4088 18564 4140
rect 19064 4088 19116 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 23480 4088 23532 4140
rect 24032 4088 24084 4140
rect 24308 4088 24360 4140
rect 8852 3952 8904 4004
rect 12532 4020 12584 4072
rect 15384 3952 15436 4004
rect 16212 4020 16264 4072
rect 17408 4020 17460 4072
rect 20720 4020 20772 4072
rect 21272 4020 21324 4072
rect 17776 3952 17828 4004
rect 18696 3952 18748 4004
rect 20260 3952 20312 4004
rect 20352 3952 20404 4004
rect 10048 3884 10100 3936
rect 10140 3884 10192 3936
rect 10692 3884 10744 3936
rect 11704 3884 11756 3936
rect 12532 3884 12584 3936
rect 19064 3884 19116 3936
rect 20536 3927 20588 3936
rect 20536 3893 20545 3927
rect 20545 3893 20579 3927
rect 20579 3893 20588 3927
rect 20536 3884 20588 3893
rect 24032 3927 24084 3936
rect 24032 3893 24041 3927
rect 24041 3893 24075 3927
rect 24075 3893 24084 3927
rect 24032 3884 24084 3893
rect 24584 3884 24636 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 1768 3680 1820 3732
rect 3332 3680 3384 3732
rect 4252 3723 4304 3732
rect 4252 3689 4261 3723
rect 4261 3689 4295 3723
rect 4295 3689 4304 3723
rect 4252 3680 4304 3689
rect 7012 3723 7064 3732
rect 7012 3689 7021 3723
rect 7021 3689 7055 3723
rect 7055 3689 7064 3723
rect 7012 3680 7064 3689
rect 7472 3723 7524 3732
rect 7472 3689 7481 3723
rect 7481 3689 7515 3723
rect 7515 3689 7524 3723
rect 7472 3680 7524 3689
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 9864 3680 9916 3732
rect 10416 3723 10468 3732
rect 10416 3689 10425 3723
rect 10425 3689 10459 3723
rect 10459 3689 10468 3723
rect 10416 3680 10468 3689
rect 2504 3612 2556 3664
rect 3424 3612 3476 3664
rect 4620 3612 4672 3664
rect 5816 3612 5868 3664
rect 11152 3680 11204 3732
rect 20076 3680 20128 3732
rect 20260 3680 20312 3732
rect 4804 3544 4856 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 7012 3544 7064 3596
rect 2228 3476 2280 3528
rect 2688 3476 2740 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 5540 3476 5592 3528
rect 6276 3476 6328 3528
rect 3424 3408 3476 3460
rect 8484 3476 8536 3528
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 9588 3476 9640 3528
rect 10140 3476 10192 3528
rect 18604 3612 18656 3664
rect 18880 3612 18932 3664
rect 21916 3680 21968 3732
rect 23480 3680 23532 3732
rect 12532 3544 12584 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 18696 3544 18748 3596
rect 19064 3544 19116 3596
rect 23204 3612 23256 3664
rect 9404 3408 9456 3460
rect 14188 3476 14240 3528
rect 15936 3476 15988 3528
rect 17316 3476 17368 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 19524 3476 19576 3528
rect 14556 3408 14608 3460
rect 20720 3476 20772 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 22376 3408 22428 3460
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 9312 3340 9364 3392
rect 11152 3340 11204 3392
rect 18236 3340 18288 3392
rect 18328 3340 18380 3392
rect 19524 3340 19576 3392
rect 21364 3340 21416 3392
rect 22100 3340 22152 3392
rect 22836 3340 22888 3392
rect 24584 3340 24636 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 6000 3136 6052 3188
rect 9404 3179 9456 3188
rect 9404 3145 9413 3179
rect 9413 3145 9447 3179
rect 9447 3145 9456 3179
rect 9404 3136 9456 3145
rect 9956 3136 10008 3188
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 3332 3000 3384 3052
rect 3516 3000 3568 3052
rect 5356 3000 5408 3052
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 7748 3000 7800 3052
rect 10968 3068 11020 3120
rect 11244 3068 11296 3120
rect 2596 2932 2648 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7656 2932 7708 2984
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11428 3000 11480 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 14188 3068 14240 3120
rect 16304 3068 16356 3120
rect 14648 3000 14700 3052
rect 17132 3000 17184 3052
rect 17500 3136 17552 3188
rect 17316 3068 17368 3120
rect 20904 3136 20956 3188
rect 23848 3136 23900 3188
rect 24124 3136 24176 3188
rect 24676 3136 24728 3188
rect 18420 3000 18472 3052
rect 18972 3000 19024 3052
rect 11796 2932 11848 2984
rect 1860 2864 1912 2916
rect 7840 2864 7892 2916
rect 6644 2796 6696 2848
rect 8852 2796 8904 2848
rect 9588 2864 9640 2916
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 21548 3068 21600 3120
rect 22192 3068 22244 3120
rect 22284 3111 22336 3120
rect 22284 3077 22293 3111
rect 22293 3077 22327 3111
rect 22327 3077 22336 3111
rect 22284 3068 22336 3077
rect 22836 3111 22888 3120
rect 22836 3077 22845 3111
rect 22845 3077 22879 3111
rect 22879 3077 22888 3111
rect 22836 3068 22888 3077
rect 19892 3000 19944 3052
rect 21916 3000 21968 3052
rect 22008 3000 22060 3052
rect 9956 2796 10008 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 14464 2864 14516 2916
rect 16580 2864 16632 2916
rect 22284 2932 22336 2984
rect 22652 3000 22704 3052
rect 24216 3000 24268 3052
rect 15016 2796 15068 2848
rect 15108 2796 15160 2848
rect 17316 2796 17368 2848
rect 17684 2796 17736 2848
rect 19892 2796 19944 2848
rect 21548 2796 21600 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 4620 2635 4672 2644
rect 4620 2601 4629 2635
rect 4629 2601 4663 2635
rect 4663 2601 4672 2635
rect 4620 2592 4672 2601
rect 7564 2592 7616 2644
rect 14924 2592 14976 2644
rect 16120 2592 16172 2644
rect 2780 2456 2832 2508
rect 9772 2524 9824 2576
rect 12164 2524 12216 2576
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 19984 2592 20036 2644
rect 22008 2592 22060 2644
rect 22192 2524 22244 2576
rect 5356 2456 5408 2508
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 2964 2388 3016 2440
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 8760 2388 8812 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 10968 2363 11020 2372
rect 10968 2329 10977 2363
rect 10977 2329 11011 2363
rect 11011 2329 11020 2363
rect 10968 2320 11020 2329
rect 12164 2388 12216 2440
rect 13912 2456 13964 2508
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 14372 2456 14424 2508
rect 15936 2456 15988 2508
rect 17316 2499 17368 2508
rect 17316 2465 17325 2499
rect 17325 2465 17359 2499
rect 17359 2465 17368 2499
rect 17316 2456 17368 2465
rect 13728 2388 13780 2440
rect 16764 2388 16816 2440
rect 12440 2320 12492 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 1676 2295 1728 2304
rect 1676 2261 1685 2295
rect 1685 2261 1719 2295
rect 1719 2261 1728 2295
rect 1676 2252 1728 2261
rect 5540 2252 5592 2304
rect 6092 2252 6144 2304
rect 7840 2252 7892 2304
rect 9128 2295 9180 2304
rect 9128 2261 9137 2295
rect 9137 2261 9171 2295
rect 9171 2261 9180 2295
rect 9128 2252 9180 2261
rect 16028 2252 16080 2304
rect 16396 2252 16448 2304
rect 19432 2388 19484 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 20536 2388 20588 2440
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 22284 2388 22336 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 19248 2320 19300 2372
rect 21272 2295 21324 2304
rect 21272 2261 21281 2295
rect 21281 2261 21315 2295
rect 21315 2261 21324 2295
rect 21272 2252 21324 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 1676 2048 1728 2100
rect 9128 2048 9180 2100
rect 17592 2048 17644 2100
rect 19432 2048 19484 2100
rect 24492 2048 24544 2100
rect 11520 1980 11572 2032
rect 11060 1912 11112 1964
rect 21272 1912 21324 1964
rect 3976 1844 4028 1896
rect 6184 1844 6236 1896
rect 7840 1844 7892 1896
rect 15660 1844 15712 1896
rect 8760 1776 8812 1828
rect 10324 1776 10376 1828
rect 10968 1776 11020 1828
rect 22100 1776 22152 1828
rect 9312 1708 9364 1760
rect 11060 1708 11112 1760
rect 20260 1232 20312 1284
rect 20812 1232 20864 1284
<< metal2 >>
rect 1030 56200 1086 57000
rect 2410 56200 2466 57000
rect 3790 56200 3846 57000
rect 5170 56200 5226 57000
rect 6550 56200 6606 57000
rect 7930 56200 7986 57000
rect 9310 56200 9366 57000
rect 10690 56200 10746 57000
rect 12070 56200 12126 57000
rect 12176 56222 12388 56250
rect 1044 53650 1072 56200
rect 2424 54126 2452 56200
rect 2412 54120 2464 54126
rect 2412 54062 2464 54068
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 3804 53650 3832 56200
rect 4068 54188 4120 54194
rect 4068 54130 4120 54136
rect 4804 54188 4856 54194
rect 4804 54130 4856 54136
rect 1032 53644 1084 53650
rect 1032 53586 1084 53592
rect 3792 53644 3844 53650
rect 3792 53586 3844 53592
rect 4080 53242 4108 54130
rect 4160 53576 4212 53582
rect 4160 53518 4212 53524
rect 4068 53236 4120 53242
rect 4068 53178 4120 53184
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 4172 52698 4200 53518
rect 4160 52692 4212 52698
rect 4160 52634 4212 52640
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 4816 51406 4844 54130
rect 5184 54126 5212 56200
rect 5172 54120 5224 54126
rect 5172 54062 5224 54068
rect 6564 53650 6592 56200
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 7380 54188 7432 54194
rect 7380 54130 7432 54136
rect 6552 53644 6604 53650
rect 6552 53586 6604 53592
rect 5540 53508 5592 53514
rect 5540 53450 5592 53456
rect 4804 51400 4856 51406
rect 4804 51342 4856 51348
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 5552 50522 5580 53450
rect 7392 51610 7420 54130
rect 7852 54126 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8576 54256 8628 54262
rect 8576 54198 8628 54204
rect 7840 54120 7892 54126
rect 7840 54062 7892 54068
rect 7840 53576 7892 53582
rect 7840 53518 7892 53524
rect 7748 53100 7800 53106
rect 7748 53042 7800 53048
rect 7380 51604 7432 51610
rect 7380 51546 7432 51552
rect 5540 50516 5592 50522
rect 5540 50458 5592 50464
rect 7760 50454 7788 53042
rect 7852 51542 7880 53518
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7840 51536 7892 51542
rect 7840 51478 7892 51484
rect 8484 51400 8536 51406
rect 8484 51342 8536 51348
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 8392 50516 8444 50522
rect 8392 50458 8444 50464
rect 7748 50448 7800 50454
rect 7748 50390 7800 50396
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 7760 48142 7788 50390
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 8404 48686 8432 50458
rect 8300 48680 8352 48686
rect 8300 48622 8352 48628
rect 8392 48680 8444 48686
rect 8392 48622 8444 48628
rect 7748 48136 7800 48142
rect 7748 48078 7800 48084
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 7760 46034 7788 48078
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 8312 47462 8340 48622
rect 8300 47456 8352 47462
rect 8300 47398 8352 47404
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 8496 46170 8524 51342
rect 8588 50386 8616 54198
rect 9324 54126 9352 56200
rect 9588 54188 9640 54194
rect 9588 54130 9640 54136
rect 9312 54120 9364 54126
rect 9312 54062 9364 54068
rect 9496 52488 9548 52494
rect 9496 52430 9548 52436
rect 8576 50380 8628 50386
rect 8576 50322 8628 50328
rect 8588 47734 8616 50322
rect 9128 48884 9180 48890
rect 9128 48826 9180 48832
rect 9140 48550 9168 48826
rect 9128 48544 9180 48550
rect 9128 48486 9180 48492
rect 8576 47728 8628 47734
rect 8576 47670 8628 47676
rect 8484 46164 8536 46170
rect 8484 46106 8536 46112
rect 7748 46028 7800 46034
rect 7748 45970 7800 45976
rect 7840 45960 7892 45966
rect 7840 45902 7892 45908
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 7852 38010 7880 45902
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 9140 44878 9168 48486
rect 9508 47802 9536 52430
rect 9600 50522 9628 54130
rect 10704 53718 10732 56200
rect 12084 56114 12112 56200
rect 12176 56114 12204 56222
rect 12084 56086 12204 56114
rect 11704 54188 11756 54194
rect 11704 54130 11756 54136
rect 10692 53712 10744 53718
rect 10692 53654 10744 53660
rect 10692 53576 10744 53582
rect 10692 53518 10744 53524
rect 10508 51400 10560 51406
rect 10508 51342 10560 51348
rect 9588 50516 9640 50522
rect 9588 50458 9640 50464
rect 9588 50244 9640 50250
rect 9588 50186 9640 50192
rect 9220 47796 9272 47802
rect 9220 47738 9272 47744
rect 9496 47796 9548 47802
rect 9496 47738 9548 47744
rect 9232 47054 9260 47738
rect 9496 47456 9548 47462
rect 9496 47398 9548 47404
rect 9220 47048 9272 47054
rect 9220 46990 9272 46996
rect 9128 44872 9180 44878
rect 9128 44814 9180 44820
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8944 42696 8996 42702
rect 8944 42638 8996 42644
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7840 38004 7892 38010
rect 7840 37946 7892 37952
rect 8852 37868 8904 37874
rect 8852 37810 8904 37816
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 3424 27532 3476 27538
rect 3424 27474 3476 27480
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1504 3398 1532 4082
rect 1780 3738 1808 4558
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 800 1532 3334
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1872 2446 1900 2858
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 1688 2106 1716 2246
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1872 800 1900 2382
rect 2240 800 2268 3470
rect 2424 3058 2452 16594
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2780 4072 2832 4078
rect 2832 4032 2912 4060
rect 2780 4014 2832 4020
rect 2504 3936 2556 3942
rect 2780 3936 2832 3942
rect 2504 3878 2556 3884
rect 2700 3884 2780 3890
rect 2700 3878 2832 3884
rect 2516 3670 2544 3878
rect 2700 3862 2820 3878
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2700 3534 2728 3862
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2608 800 2636 2926
rect 2884 2530 2912 4032
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3344 3738 3372 16934
rect 3436 8809 3464 27474
rect 7564 26920 7616 26926
rect 7564 26862 7616 26868
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3422 8800 3478 8809
rect 3422 8735 3478 8744
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 4185 3832 8298
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6497 4108 6598
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 3790 4176 3846 4185
rect 3790 4111 3846 4120
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3436 3466 3464 3606
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3528 3058 3556 3878
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2780 2508 2832 2514
rect 2884 2502 3004 2530
rect 2780 2450 2832 2456
rect 2792 1306 2820 2450
rect 2976 2446 3004 2502
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2792 1278 3004 1306
rect 2976 800 3004 1278
rect 3344 800 3372 2994
rect 3712 800 3740 4014
rect 4080 3942 4108 4082
rect 4172 4010 4200 11018
rect 4816 8362 4844 25774
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 1896 4028 1902
rect 3974 1864 3976 1873
rect 4028 1864 4030 1873
rect 3974 1799 4030 1808
rect 4080 800 4108 3878
rect 4264 3738 4292 6054
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4448 800 4476 3470
rect 4632 2650 4660 3606
rect 5184 3602 5212 15574
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4816 800 4844 3538
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5184 800 5212 2926
rect 5276 2774 5304 8298
rect 5368 3058 5396 11834
rect 5460 3058 5488 15438
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5552 3534 5580 3878
rect 5828 3670 5856 3878
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5276 2746 5396 2774
rect 5368 2514 5396 2746
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5552 800 5580 2246
rect 5920 800 5948 4082
rect 6012 3194 6040 4082
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6104 2310 6132 4966
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 6196 1902 6224 23122
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6932 19310 6960 22374
rect 6552 19304 6604 19310
rect 6920 19304 6972 19310
rect 6604 19252 6684 19258
rect 6552 19246 6684 19252
rect 6920 19246 6972 19252
rect 6564 19230 6684 19246
rect 6656 18766 6684 19230
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6656 18222 6684 18702
rect 6644 18216 6696 18222
rect 6564 18164 6644 18170
rect 6564 18158 6696 18164
rect 6564 18142 6684 18158
rect 6564 16114 6592 18142
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 13394 6500 14418
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6932 12918 6960 19246
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17338 7236 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7300 17134 7328 24754
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 12306 7052 12786
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7116 11082 7144 12718
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4622 6500 4966
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6564 4010 6592 6258
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6184 1896 6236 1902
rect 6184 1838 6236 1844
rect 6288 800 6316 3470
rect 6656 3058 6684 4558
rect 7116 4554 7144 10406
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7208 4282 7236 11290
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7392 4146 7420 4422
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7024 3738 7052 4082
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6644 3052 6696 3058
rect 6564 3012 6644 3040
rect 6564 1034 6592 3012
rect 6644 2994 6696 3000
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6656 2446 6684 2790
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6564 1006 6684 1034
rect 6656 800 6684 1006
rect 7024 800 7052 3538
rect 7392 800 7420 4082
rect 7484 3738 7512 12174
rect 7576 6662 7604 26862
rect 7668 17882 7696 30194
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7852 23730 7880 24142
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7852 22642 7880 23666
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7852 22094 7880 22578
rect 7760 22066 7880 22094
rect 8668 22092 8720 22098
rect 7760 21350 7788 22066
rect 8668 22034 8720 22040
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8576 21616 8628 21622
rect 8576 21558 8628 21564
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 7760 20398 7788 21286
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 20534 8340 21286
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8404 20398 8432 21422
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 7760 19854 7788 20334
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8496 19360 8524 21082
rect 8588 20874 8616 21558
rect 8680 21350 8708 22034
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8588 20534 8616 20810
rect 8576 20528 8628 20534
rect 8576 20470 8628 20476
rect 8588 20058 8616 20470
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8588 19446 8616 19994
rect 8668 19780 8720 19786
rect 8668 19722 8720 19728
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8404 19332 8524 19360
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 18834 8340 19110
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8312 18358 8340 18634
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 17898 8156 18158
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7760 17870 8156 17898
rect 7760 12986 7788 17870
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7852 14618 7880 17682
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 16658 8340 17478
rect 8404 17338 8432 19332
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8496 16250 8524 19178
rect 8588 18970 8616 19382
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8588 18766 8616 18906
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8576 18624 8628 18630
rect 8680 18612 8708 19722
rect 8772 19514 8800 30670
rect 8864 29306 8892 37810
rect 8956 30122 8984 42638
rect 9140 42158 9168 44814
rect 9232 44402 9260 46990
rect 9508 45082 9536 47398
rect 9496 45076 9548 45082
rect 9496 45018 9548 45024
rect 9600 44538 9628 50186
rect 10232 49156 10284 49162
rect 10232 49098 10284 49104
rect 9956 48612 10008 48618
rect 9956 48554 10008 48560
rect 9968 44946 9996 48554
rect 9956 44940 10008 44946
rect 9956 44882 10008 44888
rect 9680 44804 9732 44810
rect 9680 44746 9732 44752
rect 9588 44532 9640 44538
rect 9588 44474 9640 44480
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9312 44328 9364 44334
rect 9312 44270 9364 44276
rect 9128 42152 9180 42158
rect 9128 42094 9180 42100
rect 9036 37936 9088 37942
rect 9036 37878 9088 37884
rect 8944 30116 8996 30122
rect 8944 30058 8996 30064
rect 8852 29300 8904 29306
rect 8852 29242 8904 29248
rect 9048 27606 9076 37878
rect 9324 34202 9352 44270
rect 9692 42362 9720 44746
rect 10244 42770 10272 49098
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 44742 10456 46310
rect 10520 45558 10548 51342
rect 10704 49366 10732 53518
rect 10784 51332 10836 51338
rect 10784 51274 10836 51280
rect 10692 49360 10744 49366
rect 10692 49302 10744 49308
rect 10796 46714 10824 51274
rect 11716 49366 11744 54130
rect 12360 54126 12388 56222
rect 13450 56200 13506 57000
rect 14830 56200 14886 57000
rect 16210 56200 16266 57000
rect 17590 56200 17646 57000
rect 17696 56222 17908 56250
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 13464 53786 13492 56200
rect 14844 54194 14872 56200
rect 16224 54330 16252 56200
rect 17604 56114 17632 56200
rect 17696 56114 17724 56222
rect 17604 56086 17724 56114
rect 16212 54324 16264 54330
rect 16212 54266 16264 54272
rect 16224 54194 16252 54266
rect 17880 54210 17908 56222
rect 18970 56200 19026 57000
rect 20350 56200 20406 57000
rect 20456 56222 20668 56250
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18984 54330 19012 56200
rect 20364 56114 20392 56200
rect 20456 56114 20484 56222
rect 20364 56086 20484 56114
rect 20640 55214 20668 56222
rect 21730 56200 21786 57000
rect 23110 56200 23166 57000
rect 24490 56200 24546 57000
rect 25870 56200 25926 57000
rect 20640 55186 20760 55214
rect 18972 54324 19024 54330
rect 18972 54266 19024 54272
rect 17880 54194 18000 54210
rect 20732 54194 20760 55186
rect 21744 54194 21772 56200
rect 23124 55214 23152 56200
rect 23386 56128 23442 56137
rect 23386 56063 23442 56072
rect 23124 55186 23336 55214
rect 14464 54188 14516 54194
rect 14464 54130 14516 54136
rect 14832 54188 14884 54194
rect 14832 54130 14884 54136
rect 16212 54188 16264 54194
rect 16212 54130 16264 54136
rect 17880 54188 18012 54194
rect 17880 54182 17960 54188
rect 13544 53984 13596 53990
rect 13544 53926 13596 53932
rect 13452 53780 13504 53786
rect 13452 53722 13504 53728
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 11704 49360 11756 49366
rect 11704 49302 11756 49308
rect 10876 49156 10928 49162
rect 10876 49098 10928 49104
rect 10784 46708 10836 46714
rect 10784 46650 10836 46656
rect 10796 46594 10824 46650
rect 10612 46578 10824 46594
rect 10612 46572 10836 46578
rect 10612 46566 10784 46572
rect 10508 45552 10560 45558
rect 10508 45494 10560 45500
rect 10416 44736 10468 44742
rect 10416 44678 10468 44684
rect 10520 44266 10548 45494
rect 10508 44260 10560 44266
rect 10508 44202 10560 44208
rect 10232 42764 10284 42770
rect 10232 42706 10284 42712
rect 10612 42702 10640 46566
rect 10784 46514 10836 46520
rect 10784 46436 10836 46442
rect 10784 46378 10836 46384
rect 10796 44402 10824 46378
rect 10784 44396 10836 44402
rect 10784 44338 10836 44344
rect 10692 44192 10744 44198
rect 10692 44134 10744 44140
rect 10600 42696 10652 42702
rect 10600 42638 10652 42644
rect 9680 42356 9732 42362
rect 9680 42298 9732 42304
rect 10704 42158 10732 44134
rect 9680 42152 9732 42158
rect 9680 42094 9732 42100
rect 10692 42152 10744 42158
rect 10692 42094 10744 42100
rect 9692 35494 9720 42094
rect 10888 41818 10916 49098
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 10968 47728 11020 47734
rect 10968 47670 11020 47676
rect 10980 46714 11008 47670
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 10968 46708 11020 46714
rect 10968 46650 11020 46656
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 12808 45960 12860 45966
rect 12808 45902 12860 45908
rect 12820 45558 12848 45902
rect 13556 45558 13584 53926
rect 14476 53786 14504 54130
rect 16764 54052 16816 54058
rect 16764 53994 16816 54000
rect 15568 53984 15620 53990
rect 15568 53926 15620 53932
rect 14464 53780 14516 53786
rect 14464 53722 14516 53728
rect 15580 53582 15608 53926
rect 15568 53576 15620 53582
rect 15568 53518 15620 53524
rect 14740 53440 14792 53446
rect 14740 53382 14792 53388
rect 15660 53440 15712 53446
rect 15660 53382 15712 53388
rect 13728 48000 13780 48006
rect 13728 47942 13780 47948
rect 13636 46980 13688 46986
rect 13636 46922 13688 46928
rect 13648 46714 13676 46922
rect 13636 46708 13688 46714
rect 13636 46650 13688 46656
rect 13740 45558 13768 47942
rect 14752 46646 14780 53382
rect 14740 46640 14792 46646
rect 14740 46582 14792 46588
rect 15476 46368 15528 46374
rect 15476 46310 15528 46316
rect 15488 45898 15516 46310
rect 15672 46034 15700 53382
rect 16212 47592 16264 47598
rect 16212 47534 16264 47540
rect 15752 46504 15804 46510
rect 15752 46446 15804 46452
rect 15660 46028 15712 46034
rect 15660 45970 15712 45976
rect 15476 45892 15528 45898
rect 15476 45834 15528 45840
rect 14924 45824 14976 45830
rect 14924 45766 14976 45772
rect 12808 45552 12860 45558
rect 12808 45494 12860 45500
rect 13544 45552 13596 45558
rect 13544 45494 13596 45500
rect 13728 45552 13780 45558
rect 13728 45494 13780 45500
rect 14556 45416 14608 45422
rect 14556 45358 14608 45364
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 11520 44804 11572 44810
rect 11520 44746 11572 44752
rect 10968 44192 11020 44198
rect 10968 44134 11020 44140
rect 10876 41812 10928 41818
rect 10876 41754 10928 41760
rect 10980 41682 11008 44134
rect 11532 42294 11560 44746
rect 11704 44736 11756 44742
rect 11704 44678 11756 44684
rect 11520 42288 11572 42294
rect 11520 42230 11572 42236
rect 11532 42022 11560 42230
rect 11716 42022 11744 44678
rect 13820 44532 13872 44538
rect 13820 44474 13872 44480
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 11520 42016 11572 42022
rect 11520 41958 11572 41964
rect 11704 42016 11756 42022
rect 11704 41958 11756 41964
rect 10968 41676 11020 41682
rect 10968 41618 11020 41624
rect 10232 41608 10284 41614
rect 10232 41550 10284 41556
rect 10048 35624 10100 35630
rect 10048 35566 10100 35572
rect 9680 35488 9732 35494
rect 9680 35430 9732 35436
rect 9312 34196 9364 34202
rect 9312 34138 9364 34144
rect 9220 33992 9272 33998
rect 9220 33934 9272 33940
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 9048 26994 9076 27542
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8864 20806 8892 21422
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8628 18584 8708 18612
rect 8576 18566 8628 18572
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8588 16794 8616 17138
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7852 13954 7880 14554
rect 8312 14482 8340 14758
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8312 14074 8340 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7932 14000 7984 14006
rect 7852 13948 7932 13954
rect 7852 13942 7984 13948
rect 7852 13926 7972 13942
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7576 2650 7604 4082
rect 7668 2990 7696 12854
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7852 6118 7880 12718
rect 8220 12306 8248 12786
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8312 11558 8340 14010
rect 8404 13530 8432 15982
rect 8496 14958 8524 16186
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8588 15094 8616 16118
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8588 14618 8616 15030
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8588 14414 8616 14554
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8588 14006 8616 14350
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8588 13530 8616 13942
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8588 13258 8616 13466
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8680 12782 8708 18584
rect 8772 18358 8800 18702
rect 8864 18630 8892 20742
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 8772 13530 8800 17546
rect 8864 16726 8892 18566
rect 8956 17202 8984 26250
rect 9232 21894 9260 33934
rect 9496 32020 9548 32026
rect 9496 31962 9548 31968
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9324 21418 9352 26794
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9416 26314 9444 26522
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 9508 26042 9536 31962
rect 10060 29102 10088 35566
rect 10244 30938 10272 41550
rect 10692 39636 10744 39642
rect 10692 39578 10744 39584
rect 10704 31754 10732 39578
rect 11532 35766 11560 41958
rect 11716 35894 11744 41958
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 13832 39642 13860 44474
rect 13820 39636 13872 39642
rect 13820 39578 13872 39584
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 11716 35866 11836 35894
rect 11716 35834 11744 35866
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 11808 35494 11836 35866
rect 12348 35760 12400 35766
rect 12348 35702 12400 35708
rect 11796 35488 11848 35494
rect 11796 35430 11848 35436
rect 11808 34066 11836 35430
rect 11796 34060 11848 34066
rect 11796 34002 11848 34008
rect 10612 31726 10732 31754
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10416 29232 10468 29238
rect 10416 29174 10468 29180
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 10048 29096 10100 29102
rect 10048 29038 10100 29044
rect 10060 28762 10088 29038
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9496 24268 9548 24274
rect 9496 24210 9548 24216
rect 9508 23508 9536 24210
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9600 23798 9628 24006
rect 9692 23866 9720 28426
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9784 26450 9812 27066
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 10140 24880 10192 24886
rect 10140 24822 10192 24828
rect 9864 24132 9916 24138
rect 10152 24120 10180 24822
rect 9916 24092 10180 24120
rect 9864 24074 9916 24080
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9588 23792 9640 23798
rect 9588 23734 9640 23740
rect 9600 23526 9628 23734
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9416 23480 9536 23508
rect 9588 23520 9640 23526
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9048 18154 9076 19790
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 9140 16250 9168 18702
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9232 15706 9260 19382
rect 9324 19258 9352 20334
rect 9416 19666 9444 23480
rect 9588 23462 9640 23468
rect 9588 23248 9640 23254
rect 9588 23190 9640 23196
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9508 21622 9536 22578
rect 9496 21616 9548 21622
rect 9496 21558 9548 21564
rect 9600 19802 9628 23190
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9968 21010 9996 21490
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9508 19786 9628 19802
rect 9496 19780 9628 19786
rect 9548 19774 9628 19780
rect 9496 19722 9548 19728
rect 9416 19638 9536 19666
rect 9324 19242 9444 19258
rect 9324 19236 9456 19242
rect 9324 19230 9404 19236
rect 9404 19178 9456 19184
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9324 18358 9352 19110
rect 9416 18426 9444 19178
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9416 17338 9444 17478
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9508 17082 9536 19638
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9600 17678 9628 18090
rect 9784 18086 9812 20334
rect 10060 18970 10088 23598
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10152 22778 10180 23462
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10152 20602 10180 21830
rect 10244 21690 10272 29106
rect 10428 23866 10456 29174
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10612 23322 10640 31726
rect 12072 30184 12124 30190
rect 12360 30172 12388 35702
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12624 32768 12676 32774
rect 12624 32710 12676 32716
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 12440 30184 12492 30190
rect 12360 30144 12440 30172
rect 12072 30126 12124 30132
rect 12440 30126 12492 30132
rect 11520 30048 11572 30054
rect 11520 29990 11572 29996
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 11152 29572 11204 29578
rect 11152 29514 11204 29520
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 10784 27940 10836 27946
rect 10784 27882 10836 27888
rect 10796 27538 10824 27882
rect 10980 27878 11008 28426
rect 11060 28144 11112 28150
rect 11060 28086 11112 28092
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 10784 27532 10836 27538
rect 10784 27474 10836 27480
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 10888 27402 10916 27474
rect 10876 27396 10928 27402
rect 10876 27338 10928 27344
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10888 25362 10916 27066
rect 10980 27062 11008 27814
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 11072 26450 11100 28086
rect 11164 26926 11192 29514
rect 11440 28626 11468 29650
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11440 27674 11468 28562
rect 11532 28422 11560 29990
rect 12084 29850 12112 30126
rect 12544 30002 12572 31894
rect 12452 29974 12572 30002
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12452 29306 12480 29974
rect 12636 29306 12664 32710
rect 13360 32360 13412 32366
rect 13360 32302 13412 32308
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13372 31278 13400 32302
rect 13360 31272 13412 31278
rect 13360 31214 13412 31220
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 13372 30394 13400 31214
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 12728 30190 12756 30262
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 13360 30184 13412 30190
rect 13360 30126 13412 30132
rect 12728 29578 12756 30126
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13372 29714 13400 30126
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 12716 29572 12768 29578
rect 12716 29514 12768 29520
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 13372 29170 13400 29650
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13648 29102 13676 29990
rect 13832 29850 13860 31078
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 14108 30326 14136 30670
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 13832 29306 13860 29786
rect 13820 29300 13872 29306
rect 13820 29242 13872 29248
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 13924 29186 13952 29242
rect 13740 29158 13952 29186
rect 11612 29096 11664 29102
rect 11612 29038 11664 29044
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11428 27668 11480 27674
rect 11428 27610 11480 27616
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 11072 24750 11100 26386
rect 11164 25838 11192 26862
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11152 25832 11204 25838
rect 11152 25774 11204 25780
rect 11244 24948 11296 24954
rect 11244 24890 11296 24896
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11072 24274 11100 24550
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 11164 24154 11192 24754
rect 11256 24614 11284 24890
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11072 24126 11192 24154
rect 11072 24070 11100 24126
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10600 23316 10652 23322
rect 10600 23258 10652 23264
rect 10612 22982 10640 23258
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10428 21894 10456 21966
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10152 19786 10180 20198
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10152 19514 10180 19722
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17814 9812 18022
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9600 17270 9628 17614
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9588 17128 9640 17134
rect 9508 17076 9588 17082
rect 9508 17070 9640 17076
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9324 15706 9352 16186
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 9048 13462 9076 14282
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12782 9076 13126
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 9036 12300 9088 12306
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8220 10266 8248 10678
rect 8312 10470 8340 11494
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 7760 3058 7788 4422
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7760 800 7788 2994
rect 7852 2922 7880 4422
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8312 4146 8340 4422
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7852 2774 7880 2858
rect 7852 2746 7972 2774
rect 7944 2446 7972 2746
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7852 1902 7880 2246
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8312 1986 8340 4082
rect 8404 3738 8432 7958
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8496 3534 8524 12038
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8588 3534 8616 4422
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8588 2774 8616 3470
rect 8128 1958 8340 1986
rect 8496 2746 8616 2774
rect 7840 1896 7892 1902
rect 7840 1838 7892 1844
rect 8128 800 8156 1958
rect 8496 800 8524 2746
rect 8772 2446 8800 4422
rect 8864 4010 8892 12271
rect 9036 12242 9088 12248
rect 9048 11898 9076 12242
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9140 11762 9168 13194
rect 9232 12986 9260 15370
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 12306 9352 13398
rect 9416 12986 9444 17070
rect 9508 17054 9628 17070
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9416 12102 9444 12922
rect 9508 12442 9536 16594
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 15570 9628 15982
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15026 9628 15506
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 14482 9720 14894
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 14074 9628 14350
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9600 13938 9628 14010
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9692 13818 9720 14418
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9600 13790 9720 13818
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9416 11558 9444 11698
rect 9404 11552 9456 11558
rect 9600 11540 9628 13790
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 11898 9720 13126
rect 9784 12986 9812 14010
rect 9876 13870 9904 14554
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9968 12866 9996 16390
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 12986 10088 15302
rect 10152 15162 10180 19314
rect 10244 16454 10272 20334
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10244 14006 10272 15098
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9784 12838 9996 12866
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9404 11494 9456 11500
rect 9508 11512 9628 11540
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 10470 9168 11086
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9508 9994 9536 11512
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10130 9628 10406
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 9140 3738 9168 7482
rect 9600 7478 9628 10066
rect 9692 8906 9720 10950
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9600 5710 9628 7414
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 4690 9628 5646
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8772 1834 8800 2382
rect 8760 1828 8812 1834
rect 8760 1770 8812 1776
rect 8864 800 8892 2790
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 2106 9168 2246
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 9232 800 9260 4082
rect 9692 4078 9720 6054
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 2446 9352 3334
rect 9416 3194 9444 3402
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9600 2922 9628 3470
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9324 1766 9352 2382
rect 9312 1760 9364 1766
rect 9312 1702 9364 1708
rect 9600 800 9628 2858
rect 9784 2582 9812 12838
rect 10336 12434 10364 19110
rect 10428 16522 10456 21830
rect 10704 21554 10732 23666
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10796 21418 10824 21830
rect 10784 21412 10836 21418
rect 10784 21354 10836 21360
rect 10888 20992 10916 22918
rect 11072 22234 11100 24006
rect 11152 23792 11204 23798
rect 11152 23734 11204 23740
rect 11164 23594 11192 23734
rect 11152 23588 11204 23594
rect 11152 23530 11204 23536
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 11164 22094 11192 23530
rect 11256 22574 11284 24550
rect 11348 24342 11376 26318
rect 11336 24336 11388 24342
rect 11336 24278 11388 24284
rect 11348 24138 11376 24278
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11164 22066 11284 22094
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21690 11100 21830
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10980 21570 11008 21626
rect 10980 21542 11100 21570
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10980 21010 11008 21286
rect 10796 20964 10916 20992
rect 10968 21004 11020 21010
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10704 19922 10732 20878
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10796 18426 10824 20964
rect 10968 20946 11020 20952
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10888 19718 10916 20810
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 18834 10916 19654
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10980 18902 11008 19178
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 11072 15706 11100 21542
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 11164 18426 11192 19450
rect 11256 18970 11284 22066
rect 11348 19122 11376 22714
rect 11532 22166 11560 28358
rect 11624 26586 11652 29038
rect 12256 29028 12308 29034
rect 12256 28970 12308 28976
rect 12072 28756 12124 28762
rect 12072 28698 12124 28704
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11716 27690 11744 27950
rect 11716 27662 11836 27690
rect 11808 27606 11836 27662
rect 11796 27600 11848 27606
rect 11796 27542 11848 27548
rect 11808 27130 11836 27542
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 11900 27062 11928 27406
rect 11992 27130 12020 27474
rect 12084 27334 12112 28698
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 12164 27328 12216 27334
rect 12164 27270 12216 27276
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11612 26580 11664 26586
rect 11612 26522 11664 26528
rect 11900 26518 11928 26998
rect 12176 26994 12204 27270
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11888 26512 11940 26518
rect 11888 26454 11940 26460
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 11716 23186 11744 25434
rect 11808 23798 11836 25638
rect 11992 24138 12020 26726
rect 12164 24812 12216 24818
rect 12268 24800 12296 28970
rect 13740 28914 13768 29158
rect 13648 28886 13768 28914
rect 14096 28960 14148 28966
rect 14096 28902 14148 28908
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13556 28218 13584 28358
rect 13544 28212 13596 28218
rect 13544 28154 13596 28160
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12636 27674 12664 27950
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12636 27470 12664 27610
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12636 26042 12664 27270
rect 13096 26994 13124 27542
rect 13360 27532 13412 27538
rect 13280 27492 13360 27520
rect 13280 27062 13308 27492
rect 13360 27474 13412 27480
rect 13648 27062 13676 28886
rect 14108 28626 14136 28902
rect 14568 28762 14596 45358
rect 14936 44810 14964 45766
rect 14924 44804 14976 44810
rect 14924 44746 14976 44752
rect 15764 37942 15792 46446
rect 16028 45008 16080 45014
rect 16028 44950 16080 44956
rect 15844 42084 15896 42090
rect 15844 42026 15896 42032
rect 15752 37936 15804 37942
rect 15752 37878 15804 37884
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15396 32502 15424 33866
rect 15384 32496 15436 32502
rect 15384 32438 15436 32444
rect 15016 31408 15068 31414
rect 15016 31350 15068 31356
rect 15028 31210 15056 31350
rect 15016 31204 15068 31210
rect 15016 31146 15068 31152
rect 15396 30938 15424 32438
rect 15384 30932 15436 30938
rect 15384 30874 15436 30880
rect 15396 30734 15424 30874
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 15028 29238 15056 29446
rect 15016 29232 15068 29238
rect 15016 29174 15068 29180
rect 15028 28966 15056 29174
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 14556 28756 14608 28762
rect 14556 28698 14608 28704
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13832 27402 13860 27814
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13268 27056 13320 27062
rect 13268 26998 13320 27004
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 12716 26512 12768 26518
rect 12716 26454 12768 26460
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12452 25430 12480 25638
rect 12440 25424 12492 25430
rect 12440 25366 12492 25372
rect 12216 24772 12296 24800
rect 12164 24754 12216 24760
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 11980 24132 12032 24138
rect 11980 24074 12032 24080
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11808 22506 11836 23122
rect 11796 22500 11848 22506
rect 11796 22442 11848 22448
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 11808 21690 11836 21898
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11992 19922 12020 24074
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11624 19174 11652 19722
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11716 19514 11744 19654
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11612 19168 11664 19174
rect 11348 19094 11560 19122
rect 11612 19110 11664 19116
rect 11244 18964 11296 18970
rect 11296 18924 11376 18952
rect 11244 18906 11296 18912
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11256 18426 11284 18634
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11164 17678 11192 18362
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11164 17134 11192 17614
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11256 16794 11284 18362
rect 11348 17678 11376 18924
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11348 17202 11376 17274
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11256 16658 11284 16730
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11348 15162 11376 17138
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11440 15042 11468 18566
rect 11532 18426 11560 19094
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11808 18154 11836 19450
rect 12084 18698 12112 22918
rect 12360 22642 12388 24210
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12360 22114 12388 22578
rect 12360 22086 12480 22114
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11624 16250 11652 16662
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 11348 15014 11468 15042
rect 11612 15020 11664 15026
rect 10520 12442 10548 14962
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11164 14278 11192 14758
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 12986 11100 13806
rect 11164 13258 11192 14214
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10244 12406 10364 12434
rect 10508 12436 10560 12442
rect 10244 11830 10272 12406
rect 10508 12378 10560 12384
rect 11072 12374 11100 12718
rect 11164 12714 11192 13194
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11256 12434 11284 14214
rect 11348 12646 11376 15014
rect 11612 14962 11664 14968
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11164 12406 11284 12434
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 11082 10180 11494
rect 10612 11354 10640 12038
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10152 10674 10180 11018
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10704 9110 10732 12038
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11072 11150 11100 11630
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10538 10916 10950
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 9994 11008 10406
rect 11072 10266 11100 11086
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10692 9104 10744 9110
rect 10046 9072 10102 9081
rect 10692 9046 10744 9052
rect 10046 9007 10102 9016
rect 11060 9036 11112 9042
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9876 3738 9904 8570
rect 9954 7440 10010 7449
rect 9954 7375 10010 7384
rect 9968 4690 9996 7375
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10060 4282 10088 9007
rect 11060 8978 11112 8984
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 7342 11008 8774
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 5778 10824 7142
rect 10980 6254 11008 7278
rect 11072 6866 11100 8978
rect 11164 8362 11192 12406
rect 11440 12102 11468 14826
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11244 11552 11296 11558
rect 11440 11540 11468 12038
rect 11296 11512 11468 11540
rect 11244 11494 11296 11500
rect 11256 11286 11284 11494
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10470 11284 10950
rect 11532 10577 11560 12106
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10876 6248 10928 6254
rect 10874 6216 10876 6225
rect 10968 6248 11020 6254
rect 10928 6216 10930 6225
rect 10968 6190 11020 6196
rect 10874 6151 10930 6160
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9968 3194 9996 4014
rect 10060 3942 10088 4014
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3534 10180 3878
rect 10428 3738 10456 5510
rect 11072 5234 11100 6802
rect 11164 6458 11192 7278
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9968 800 9996 2790
rect 10324 1828 10376 1834
rect 10324 1770 10376 1776
rect 10336 800 10364 1770
rect 10704 800 10732 3878
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 10980 2854 11008 3062
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10980 1834 11008 2314
rect 11072 1970 11100 4558
rect 11164 3738 11192 6258
rect 11256 5794 11284 10406
rect 11624 10266 11652 14962
rect 11716 14482 11744 16594
rect 11808 16182 11836 17614
rect 12084 17542 12112 17818
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 12084 16998 12112 17478
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 12084 15638 12112 16934
rect 12176 15978 12204 21558
rect 12360 21146 12388 21830
rect 12452 21554 12480 22086
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12452 20466 12480 21490
rect 12544 20602 12572 23190
rect 12636 22094 12664 25842
rect 12728 25294 12756 26454
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12728 24410 12756 25094
rect 12820 24818 12848 26930
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13450 25800 13506 25809
rect 13450 25735 13452 25744
rect 13504 25735 13506 25744
rect 13452 25706 13504 25712
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13556 25401 13584 25638
rect 13542 25392 13598 25401
rect 13542 25327 13598 25336
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12912 23594 12940 24346
rect 12900 23588 12952 23594
rect 12900 23530 12952 23536
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12820 22166 12848 23462
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 13280 22438 13308 22986
rect 13372 22574 13400 25230
rect 13544 24880 13596 24886
rect 13544 24822 13596 24828
rect 13556 24138 13584 24822
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13740 23730 13768 27270
rect 13912 25968 13964 25974
rect 13912 25910 13964 25916
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13832 23866 13860 25638
rect 13924 24834 13952 25910
rect 14108 25838 14136 28562
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14740 27532 14792 27538
rect 14740 27474 14792 27480
rect 14280 26512 14332 26518
rect 14280 26454 14332 26460
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 13924 24806 14044 24834
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13924 24070 13952 24686
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13924 23662 13952 24006
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12636 22066 12756 22094
rect 12728 21842 12756 22066
rect 12636 21814 12756 21842
rect 12636 21010 12664 21814
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12452 19922 12480 20402
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12452 19378 12480 19858
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18426 12480 19314
rect 12544 18970 12572 19654
rect 12728 18970 12756 21626
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 21146 13400 22510
rect 14016 21350 14044 24806
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14108 22710 14136 24006
rect 14292 23798 14320 26454
rect 14752 26382 14780 27474
rect 14844 27470 14872 28358
rect 15028 28218 15056 28902
rect 15120 28558 15148 30602
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15212 29306 15240 29446
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15016 28212 15068 28218
rect 15016 28154 15068 28160
rect 15120 27674 15148 28494
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14832 26444 14884 26450
rect 14832 26386 14884 26392
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 22030 14136 22374
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21486 14136 21966
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12440 18420 12492 18426
rect 12492 18380 12572 18408
rect 12440 18362 12492 18368
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12452 17610 12480 18226
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12452 17338 12480 17546
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12256 15972 12308 15978
rect 12256 15914 12308 15920
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 12268 15570 12296 15914
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 14618 11836 14962
rect 12084 14822 12112 15098
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 13734 12204 14418
rect 12452 14396 12480 17138
rect 12544 16658 12572 18380
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 14498 12572 15370
rect 12636 14618 12664 18634
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 17202 12848 18566
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17746 13400 21082
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17338 13216 17478
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 13464 17134 13492 20334
rect 14200 20058 14228 23666
rect 14476 23202 14504 26182
rect 14752 25362 14780 26318
rect 14844 25362 14872 26386
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14752 24750 14780 25298
rect 14844 24954 14872 25298
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14936 23866 14964 26726
rect 15016 26240 15068 26246
rect 15016 26182 15068 26188
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14924 23724 14976 23730
rect 15028 23712 15056 26182
rect 15108 25968 15160 25974
rect 15212 25956 15240 28970
rect 15160 25928 15240 25956
rect 15108 25910 15160 25916
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 14976 23684 15056 23712
rect 14924 23666 14976 23672
rect 14292 23174 14504 23202
rect 14292 23118 14320 23174
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14384 22778 14412 23054
rect 14936 23050 14964 23666
rect 14924 23044 14976 23050
rect 14924 22986 14976 22992
rect 14936 22778 14964 22986
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 14648 22704 14700 22710
rect 14648 22646 14700 22652
rect 14660 22438 14688 22646
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14660 21622 14688 22374
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21622 14872 21830
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 15120 21486 15148 24686
rect 15212 24682 15240 25230
rect 15304 25226 15332 29582
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15396 27946 15424 28562
rect 15856 28218 15884 42026
rect 16040 30274 16068 44950
rect 16224 35894 16252 47534
rect 16488 46028 16540 46034
rect 16488 45970 16540 45976
rect 16224 35866 16344 35894
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16132 31890 16160 32914
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16132 31278 16160 31826
rect 16120 31272 16172 31278
rect 16120 31214 16172 31220
rect 16040 30246 16160 30274
rect 16028 30184 16080 30190
rect 16028 30126 16080 30132
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15948 29238 15976 29990
rect 16040 29714 16068 30126
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 16132 28994 16160 30246
rect 16212 29300 16264 29306
rect 16212 29242 16264 29248
rect 16040 28966 16160 28994
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15948 28694 15976 28902
rect 15936 28688 15988 28694
rect 15936 28630 15988 28636
rect 15844 28212 15896 28218
rect 15844 28154 15896 28160
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 15568 27328 15620 27334
rect 15566 27296 15568 27305
rect 15660 27328 15712 27334
rect 15620 27296 15622 27305
rect 15660 27270 15712 27276
rect 15566 27231 15622 27240
rect 15672 27146 15700 27270
rect 15580 27130 15700 27146
rect 15568 27124 15700 27130
rect 15620 27118 15700 27124
rect 15568 27066 15620 27072
rect 15752 26920 15804 26926
rect 15752 26862 15804 26868
rect 15764 26586 15792 26862
rect 15752 26580 15804 26586
rect 15752 26522 15804 26528
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15384 25832 15436 25838
rect 15384 25774 15436 25780
rect 15396 25430 15424 25774
rect 15384 25424 15436 25430
rect 15384 25366 15436 25372
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15304 24954 15332 25162
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15304 24857 15332 24890
rect 15290 24848 15346 24857
rect 15290 24783 15346 24792
rect 15396 24750 15424 25094
rect 15488 24954 15516 26386
rect 15856 26246 15884 28154
rect 15948 26994 15976 28630
rect 16040 28422 16068 28966
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 16040 27402 16068 28358
rect 16028 27396 16080 27402
rect 16028 27338 16080 27344
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15948 26450 15976 26930
rect 16028 26512 16080 26518
rect 16028 26454 16080 26460
rect 15936 26444 15988 26450
rect 15936 26386 15988 26392
rect 16040 26330 16068 26454
rect 15948 26314 16068 26330
rect 15936 26308 16068 26314
rect 15988 26302 16068 26308
rect 15936 26250 15988 26256
rect 15844 26240 15896 26246
rect 15844 26182 15896 26188
rect 16224 25650 16252 29242
rect 16316 28082 16344 35866
rect 16500 32026 16528 45970
rect 16776 35894 16804 53994
rect 17040 53984 17092 53990
rect 17040 53926 17092 53932
rect 17052 53582 17080 53926
rect 17880 53786 17908 54182
rect 17960 54130 18012 54136
rect 20720 54188 20772 54194
rect 20720 54130 20772 54136
rect 21732 54188 21784 54194
rect 21732 54130 21784 54136
rect 18788 54052 18840 54058
rect 18788 53994 18840 54000
rect 18604 53984 18656 53990
rect 18604 53926 18656 53932
rect 17868 53780 17920 53786
rect 17868 53722 17920 53728
rect 18616 53582 18644 53926
rect 17040 53576 17092 53582
rect 17040 53518 17092 53524
rect 18604 53576 18656 53582
rect 18604 53518 18656 53524
rect 17684 53440 17736 53446
rect 17684 53382 17736 53388
rect 17696 44946 17724 53382
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17684 44940 17736 44946
rect 17684 44882 17736 44888
rect 17500 44804 17552 44810
rect 17500 44746 17552 44752
rect 17512 44538 17540 44746
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17500 44532 17552 44538
rect 17500 44474 17552 44480
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 16856 41608 16908 41614
rect 16856 41550 16908 41556
rect 16592 35866 16804 35894
rect 16592 33114 16620 35866
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16592 32910 16620 33050
rect 16580 32904 16632 32910
rect 16580 32846 16632 32852
rect 16764 32360 16816 32366
rect 16764 32302 16816 32308
rect 16488 32020 16540 32026
rect 16488 31962 16540 31968
rect 16672 31884 16724 31890
rect 16672 31826 16724 31832
rect 16684 31482 16712 31826
rect 16776 31822 16804 32302
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16672 31476 16724 31482
rect 16672 31418 16724 31424
rect 16776 31346 16804 31758
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16868 30274 16896 41550
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17040 39976 17092 39982
rect 17040 39918 17092 39924
rect 16948 38548 17000 38554
rect 16948 38490 17000 38496
rect 16960 31754 16988 38490
rect 17052 35894 17080 39918
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 17052 35866 17172 35894
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 18800 35894 18828 53994
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23308 53650 23336 55186
rect 23296 53644 23348 53650
rect 23296 53586 23348 53592
rect 22284 53576 22336 53582
rect 22284 53518 22336 53524
rect 21456 53508 21508 53514
rect 21456 53450 21508 53456
rect 19984 53440 20036 53446
rect 19984 53382 20036 53388
rect 19800 49904 19852 49910
rect 19800 49846 19852 49852
rect 19524 43784 19576 43790
rect 19524 43726 19576 43732
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17144 32366 17172 35866
rect 18708 35866 18828 35894
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17316 32904 17368 32910
rect 17316 32846 17368 32852
rect 17224 32836 17276 32842
rect 17224 32778 17276 32784
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 16960 31726 17080 31754
rect 16776 30258 16896 30274
rect 16764 30252 16896 30258
rect 16816 30246 16896 30252
rect 16764 30194 16816 30200
rect 16488 30184 16540 30190
rect 16488 30126 16540 30132
rect 16500 29782 16528 30126
rect 16776 30054 16804 30194
rect 17052 30122 17080 31726
rect 17144 31686 17172 32302
rect 17132 31680 17184 31686
rect 17132 31622 17184 31628
rect 17040 30116 17092 30122
rect 17040 30058 17092 30064
rect 16672 30048 16724 30054
rect 16672 29990 16724 29996
rect 16764 30048 16816 30054
rect 16764 29990 16816 29996
rect 16488 29776 16540 29782
rect 16488 29718 16540 29724
rect 16500 29578 16528 29718
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 16500 28914 16528 29514
rect 16580 29028 16632 29034
rect 16580 28970 16632 28976
rect 16408 28886 16528 28914
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16316 27878 16344 28018
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16316 26314 16344 27814
rect 16304 26308 16356 26314
rect 16304 26250 16356 26256
rect 15764 25622 16252 25650
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15304 21962 15332 22578
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14568 20534 14596 20742
rect 14556 20528 14608 20534
rect 14556 20470 14608 20476
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14476 19310 14504 20198
rect 14568 19378 14596 20470
rect 15120 20398 15148 21422
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14568 19174 14596 19314
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13832 18426 13860 18702
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13924 18222 13952 18566
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 12716 16992 12768 16998
rect 12768 16940 12848 16946
rect 12716 16934 12848 16940
rect 12728 16918 12848 16934
rect 12820 16658 12848 16918
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12544 14470 12664 14498
rect 12452 14368 12572 14396
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11532 9674 11560 9930
rect 11348 9654 11560 9674
rect 11348 9648 11572 9654
rect 11348 9646 11520 9648
rect 11348 9382 11376 9646
rect 11520 9590 11572 9596
rect 11716 9586 11744 13330
rect 11900 12986 11928 13670
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11900 12850 11928 12922
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11808 12238 11836 12650
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11900 11218 11928 12378
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11978 11112 12034 11121
rect 11978 11047 12034 11056
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11426 9480 11482 9489
rect 11426 9415 11482 9424
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 8906 11376 9318
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11348 7546 11376 8842
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11348 7410 11376 7482
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11348 6254 11376 6666
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 5914 11376 6190
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11256 5766 11376 5794
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 3058 11192 3334
rect 11256 3126 11284 4626
rect 11348 4282 11376 5766
rect 11440 5166 11468 9415
rect 11716 9042 11744 9522
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11624 7954 11652 8434
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11716 7886 11744 8366
rect 11992 8090 12020 11047
rect 12084 10266 12112 13126
rect 12176 12442 12204 13126
rect 12268 12986 12296 13806
rect 12452 13326 12480 13942
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12544 12986 12572 14368
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 10810 12204 12242
rect 12268 11014 12296 12922
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12360 12646 12388 12854
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11762 12388 12038
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12440 11688 12492 11694
rect 12346 11656 12402 11665
rect 12440 11630 12492 11636
rect 12346 11591 12348 11600
rect 12400 11591 12402 11600
rect 12348 11562 12400 11568
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12176 10130 12204 10746
rect 12452 10470 12480 11630
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12440 10192 12492 10198
rect 12440 10134 12492 10140
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12084 9178 12112 9862
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12452 8650 12480 10134
rect 12544 8906 12572 12718
rect 12636 12442 12664 14470
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12728 11898 12756 15302
rect 12820 15162 12848 16594
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13464 16266 13492 16526
rect 13556 16402 13584 16662
rect 13648 16590 13676 17002
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13636 16448 13688 16454
rect 13556 16396 13636 16402
rect 13556 16390 13688 16396
rect 13556 16374 13676 16390
rect 13464 16250 13584 16266
rect 13464 16244 13596 16250
rect 13464 16238 13544 16244
rect 13544 16186 13596 16192
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13556 15502 13584 16186
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14600 12848 14758
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12820 14572 12940 14600
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12820 11830 12848 14214
rect 12912 13802 12940 14572
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 14074 13584 14214
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12912 12782 12940 13398
rect 13464 13394 13492 13806
rect 13648 13530 13676 16374
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 13358 11792 13414 11801
rect 13358 11727 13414 11736
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12360 8622 12480 8650
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11532 7002 11560 7346
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11532 6730 11560 6938
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11532 5778 11560 6666
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11532 5370 11560 5714
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11440 4146 11468 5102
rect 11532 5030 11560 5306
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11060 1964 11112 1970
rect 11060 1906 11112 1912
rect 10968 1828 11020 1834
rect 10968 1770 11020 1776
rect 11060 1760 11112 1766
rect 11060 1702 11112 1708
rect 11072 800 11100 1702
rect 11440 800 11468 2994
rect 11624 2774 11652 7686
rect 11900 7546 11928 7890
rect 12360 7546 12388 8622
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12452 5574 12480 7822
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12084 4826 12112 5102
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12254 4584 12310 4593
rect 12452 4570 12480 5510
rect 12544 5370 12572 8298
rect 12636 7886 12664 11630
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12728 9602 12756 11562
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12820 10810 12848 11222
rect 12912 11082 12940 11222
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12820 10062 12848 10542
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 13372 9926 13400 11727
rect 13464 11370 13492 12922
rect 13556 12345 13584 13330
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13542 12336 13598 12345
rect 13542 12271 13598 12280
rect 13648 12170 13676 12786
rect 13740 12306 13768 18022
rect 13924 17882 13952 18158
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 14108 16522 14136 19110
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 17678 14320 18566
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14568 16794 14596 19110
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14108 16182 14136 16458
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13832 15366 13860 15982
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13832 13530 13860 13942
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13832 12442 13860 13466
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13542 11928 13598 11937
rect 13542 11863 13544 11872
rect 13596 11863 13598 11872
rect 13544 11834 13596 11840
rect 13740 11694 13768 12242
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13464 11342 13768 11370
rect 13544 11280 13596 11286
rect 13542 11248 13544 11257
rect 13596 11248 13598 11257
rect 13542 11183 13598 11192
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13464 9722 13492 10406
rect 13648 10130 13676 11154
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 12728 9574 12848 9602
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 8090 12756 9454
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7546 12664 7686
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12728 6866 12756 8026
rect 12820 7970 12848 9574
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12912 8634 12940 8842
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12820 7942 12940 7970
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12636 4622 12664 6666
rect 12714 6488 12770 6497
rect 12820 6458 12848 7754
rect 12912 7750 12940 7942
rect 13372 7886 13400 8366
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12714 6423 12770 6432
rect 12808 6452 12860 6458
rect 12728 6390 12756 6423
rect 12808 6394 12860 6400
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12912 6202 12940 6870
rect 13450 6760 13506 6769
rect 13450 6695 13506 6704
rect 13464 6662 13492 6695
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13450 6352 13506 6361
rect 13450 6287 13506 6296
rect 13464 6254 13492 6287
rect 12992 6248 13044 6254
rect 12820 6174 12940 6202
rect 12990 6216 12992 6225
rect 13452 6248 13504 6254
rect 13044 6216 13046 6225
rect 12820 4758 12848 6174
rect 13452 6190 13504 6196
rect 12990 6151 13046 6160
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13556 5710 13584 9862
rect 13648 9042 13676 10066
rect 13740 9110 13768 11342
rect 13924 10810 13952 14282
rect 14016 12374 14044 16118
rect 14292 16114 14320 16390
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14292 15638 14320 16050
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 12782 14136 13670
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13924 9722 13952 9930
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14016 9586 14044 12038
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14108 9518 14136 12718
rect 14200 11898 14228 15302
rect 14292 15162 14320 15302
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14476 15026 14504 15982
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14384 11830 14412 14214
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14292 10742 14320 10950
rect 14384 10810 14412 10950
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14280 10736 14332 10742
rect 14280 10678 14332 10684
rect 14476 10606 14504 14962
rect 14660 14890 14688 19858
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 16250 15056 16390
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15366 14780 16050
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14752 14482 14780 15302
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12374 14596 12786
rect 14752 12646 14780 13126
rect 14936 12986 14964 14418
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14738 12472 14794 12481
rect 14738 12407 14794 12416
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14752 12238 14780 12407
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14740 12232 14792 12238
rect 14660 12192 14740 12220
rect 14556 12096 14608 12102
rect 14660 12084 14688 12192
rect 14740 12174 14792 12180
rect 14608 12056 14688 12084
rect 14556 12038 14608 12044
rect 14936 11694 14964 12242
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 14740 11688 14792 11694
rect 14660 11648 14740 11676
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14554 10568 14610 10577
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13832 8566 13860 9318
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13818 8392 13874 8401
rect 14016 8362 14044 8842
rect 13818 8327 13874 8336
rect 14004 8356 14056 8362
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13740 7954 13768 8026
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13648 6390 13676 7482
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13648 5370 13676 6326
rect 13740 6186 13768 6734
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13360 5296 13412 5302
rect 13082 5264 13138 5273
rect 13412 5244 13492 5250
rect 13360 5238 13492 5244
rect 13372 5222 13492 5238
rect 13082 5199 13084 5208
rect 13136 5199 13138 5208
rect 13084 5170 13136 5176
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12624 4616 12676 4622
rect 12452 4542 12572 4570
rect 12624 4558 12676 4564
rect 12254 4519 12310 4528
rect 12268 4146 12296 4519
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11716 3058 11744 3878
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11532 2746 11652 2774
rect 11532 2038 11560 2746
rect 11520 2032 11572 2038
rect 11520 1974 11572 1980
rect 11808 800 11836 2926
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12176 2446 12204 2518
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12176 800 12204 2382
rect 12452 2378 12480 4422
rect 12544 4078 12572 4542
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13268 4548 13320 4554
rect 13268 4490 13320 4496
rect 13188 4214 13216 4490
rect 13280 4282 13308 4490
rect 13464 4486 13492 5222
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12544 3602 12572 3878
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12544 800 12572 3538
rect 12820 1714 12848 3538
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 1686 12940 1714
rect 12912 800 12940 1686
rect 13280 800 13308 2314
rect 13648 800 13676 2926
rect 13740 2446 13768 5782
rect 13832 4214 13860 8327
rect 14004 8298 14056 8304
rect 14292 7750 14320 10542
rect 14554 10503 14610 10512
rect 14568 10266 14596 10503
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14476 9518 14504 10066
rect 14556 9716 14608 9722
rect 14660 9704 14688 11648
rect 14740 11630 14792 11636
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 15028 11558 15056 11766
rect 15120 11665 15148 19110
rect 15212 17814 15240 21830
rect 15488 21570 15516 23530
rect 15580 22166 15608 25094
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15672 23118 15700 23598
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15488 21542 15608 21570
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15212 14822 15240 14962
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15212 13394 15240 14758
rect 15304 13462 15332 21286
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15396 16998 15424 20402
rect 15488 19514 15516 21354
rect 15580 20058 15608 21542
rect 15672 20806 15700 21626
rect 15764 21554 15792 25622
rect 16302 25256 16358 25265
rect 16302 25191 16358 25200
rect 16316 25158 16344 25191
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16408 24818 16436 28886
rect 16488 28756 16540 28762
rect 16488 28698 16540 28704
rect 16500 27674 16528 28698
rect 16488 27668 16540 27674
rect 16488 27610 16540 27616
rect 16500 27470 16528 27610
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15580 17542 15608 19994
rect 15672 19854 15700 20742
rect 15764 20058 15792 20810
rect 15948 20602 15976 24550
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15764 19242 15792 19994
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15488 16454 15516 17478
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15200 13388 15252 13394
rect 15396 13376 15424 15846
rect 15488 15706 15516 15914
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15580 14550 15608 17070
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15672 16250 15700 16526
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15764 15450 15792 17478
rect 15856 16794 15884 19926
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15672 15422 15792 15450
rect 15672 14958 15700 15422
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15162 15792 15302
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 15580 13870 15608 14486
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15476 13388 15528 13394
rect 15396 13348 15476 13376
rect 15200 13330 15252 13336
rect 15476 13330 15528 13336
rect 15212 12782 15240 13330
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15106 11656 15162 11665
rect 15106 11591 15162 11600
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14608 9676 14688 9704
rect 14556 9658 14608 9664
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14384 8514 14412 9454
rect 14476 9042 14504 9454
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8838 14504 8978
rect 14568 8838 14596 9658
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14476 8634 14504 8774
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14384 8486 14504 8514
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7478 14320 7686
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13924 5302 13952 6938
rect 14370 6896 14426 6905
rect 14370 6831 14372 6840
rect 14424 6831 14426 6840
rect 14372 6802 14424 6808
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14016 5914 14044 6326
rect 14186 5944 14242 5953
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14108 5888 14186 5896
rect 14108 5868 14188 5888
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13924 4146 13952 4966
rect 14016 4690 14044 5102
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14108 4026 14136 5868
rect 14240 5879 14242 5888
rect 14188 5850 14240 5856
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4826 14228 4966
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 13924 3998 14136 4026
rect 13924 2514 13952 3998
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 14016 800 14044 3538
rect 14200 3534 14228 4558
rect 14292 4214 14320 5306
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14200 2514 14228 3062
rect 14476 2922 14504 8486
rect 14568 3466 14596 8774
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14660 3058 14688 8298
rect 14752 7970 14780 9862
rect 14844 8090 14872 10678
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14936 10062 14964 10202
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 15028 9908 15056 11494
rect 15212 11082 15240 11766
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 14936 9880 15056 9908
rect 14936 8906 14964 9880
rect 15120 9450 15148 11018
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 15028 8498 15056 9114
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15120 8378 15148 8774
rect 15028 8350 15148 8378
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14752 7942 14872 7970
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14752 7002 14780 7414
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 5914 14780 6598
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14740 5296 14792 5302
rect 14738 5264 14740 5273
rect 14792 5264 14794 5273
rect 14738 5199 14794 5208
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14384 800 14412 2450
rect 14752 800 14780 2926
rect 14844 2774 14872 7942
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14936 4622 14964 7890
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15028 2854 15056 8350
rect 15212 8022 15240 11018
rect 15304 10305 15332 12038
rect 15396 11354 15424 13126
rect 15488 12646 15516 13330
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10470 15424 10542
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15290 10296 15346 10305
rect 15290 10231 15346 10240
rect 15304 9654 15332 10231
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15304 9042 15332 9590
rect 15396 9382 15424 10406
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15396 7732 15424 8842
rect 15488 7954 15516 11494
rect 15580 10810 15608 12854
rect 15672 11558 15700 13874
rect 15764 13394 15792 14554
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15568 9512 15620 9518
rect 15672 9500 15700 11290
rect 15764 9518 15792 13330
rect 15856 12782 15884 13738
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 12306 15884 12718
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15856 10130 15884 12242
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15620 9472 15700 9500
rect 15752 9512 15804 9518
rect 15568 9454 15620 9460
rect 15752 9454 15804 9460
rect 15580 8906 15608 9454
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15476 7744 15528 7750
rect 15396 7704 15476 7732
rect 15476 7686 15528 7692
rect 15198 7304 15254 7313
rect 15198 7239 15254 7248
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 5710 15148 7142
rect 15212 6225 15240 7239
rect 15382 6352 15438 6361
rect 15382 6287 15384 6296
rect 15436 6287 15438 6296
rect 15384 6258 15436 6264
rect 15198 6216 15254 6225
rect 15198 6151 15254 6160
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 4690 15148 5646
rect 15212 5642 15240 6151
rect 15488 5817 15516 7686
rect 15474 5808 15530 5817
rect 15384 5772 15436 5778
rect 15474 5743 15530 5752
rect 15384 5714 15436 5720
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15396 4690 15424 5714
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15396 4010 15424 4626
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 14844 2746 14964 2774
rect 14936 2650 14964 2746
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15120 800 15148 2790
rect 15488 800 15516 3538
rect 15580 2774 15608 8842
rect 15764 8566 15792 9454
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15764 7954 15792 8502
rect 15856 8090 15884 8910
rect 15948 8650 15976 17002
rect 16040 12209 16068 17682
rect 16132 17678 16160 22374
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16224 21894 16252 22170
rect 16500 22094 16528 27270
rect 16592 27062 16620 28970
rect 16580 27056 16632 27062
rect 16580 26998 16632 27004
rect 16684 26382 16712 29990
rect 16776 26518 16804 29990
rect 17144 28218 17172 31622
rect 17236 29170 17264 32778
rect 17328 29186 17356 32846
rect 17500 32836 17552 32842
rect 17500 32778 17552 32784
rect 17512 32570 17540 32778
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 17500 32564 17552 32570
rect 17500 32506 17552 32512
rect 17592 32496 17644 32502
rect 17592 32438 17644 32444
rect 17604 31890 17632 32438
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 17592 31884 17644 31890
rect 17512 31844 17592 31872
rect 17512 31754 17540 31844
rect 17592 31826 17644 31832
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17512 31726 17632 31754
rect 17328 29170 17540 29186
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17316 29164 17552 29170
rect 17368 29158 17500 29164
rect 17316 29106 17368 29112
rect 17500 29106 17552 29112
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27130 16896 27814
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16764 26512 16816 26518
rect 16764 26454 16816 26460
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16592 22982 16620 23802
rect 16684 23730 16712 26318
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 16868 25362 16896 25978
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16868 22778 16896 22986
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16408 22066 16528 22094
rect 16764 22092 16816 22098
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 21146 16252 21830
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16132 16794 16160 17206
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16132 14006 16160 16730
rect 16224 16658 16252 21082
rect 16408 19378 16436 22066
rect 16764 22034 16816 22040
rect 16776 21010 16804 22034
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 17134 16344 17478
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16224 15910 16252 16390
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16132 13546 16160 13942
rect 16132 13518 16252 13546
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16132 12986 16160 13330
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16026 12200 16082 12209
rect 16026 12135 16082 12144
rect 16040 11937 16068 12135
rect 16026 11928 16082 11937
rect 16026 11863 16082 11872
rect 16040 11694 16068 11863
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 11257 16068 11494
rect 16026 11248 16082 11257
rect 16026 11183 16082 11192
rect 16224 11064 16252 13518
rect 16316 12102 16344 16934
rect 16408 16658 16436 17274
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16408 15570 16436 16594
rect 16684 15978 16712 18770
rect 16776 18290 16804 20946
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16868 18329 16896 18362
rect 16854 18320 16910 18329
rect 16764 18284 16816 18290
rect 16854 18255 16910 18264
rect 16764 18226 16816 18232
rect 16776 17338 16804 18226
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16868 14958 16896 18090
rect 16960 17814 16988 26250
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 17052 22438 17080 25978
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17144 25809 17172 25842
rect 17130 25800 17186 25809
rect 17130 25735 17186 25744
rect 17236 24954 17264 26182
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17328 23866 17356 29106
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17420 28014 17448 29038
rect 17500 29028 17552 29034
rect 17500 28970 17552 28976
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17408 25696 17460 25702
rect 17406 25664 17408 25673
rect 17460 25664 17462 25673
rect 17406 25599 17462 25608
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17236 22817 17264 23258
rect 17222 22808 17278 22817
rect 17222 22743 17278 22752
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17144 20534 17172 21830
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17144 19990 17172 20470
rect 17236 20058 17264 20742
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17052 19786 17080 19926
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17236 19514 17264 19858
rect 17328 19514 17356 23462
rect 17512 22094 17540 28970
rect 17604 27878 17632 31726
rect 17696 31278 17724 31826
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 17696 29458 17724 31214
rect 18420 31136 18472 31142
rect 18420 31078 18472 31084
rect 18432 30666 18460 31078
rect 18524 30938 18552 31962
rect 18708 31754 18736 35866
rect 19064 35556 19116 35562
rect 19064 35498 19116 35504
rect 18616 31726 18736 31754
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 18420 30660 18472 30666
rect 18420 30602 18472 30608
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18432 29646 18460 30602
rect 18420 29640 18472 29646
rect 18420 29582 18472 29588
rect 17696 29430 17816 29458
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17590 25392 17646 25401
rect 17590 25327 17646 25336
rect 17604 25294 17632 25327
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17696 24206 17724 27882
rect 17788 27538 17816 29430
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18432 29170 18460 29582
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 18432 28966 18460 29106
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 28558 18460 28902
rect 18616 28762 18644 31726
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30938 18736 31214
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18696 30592 18748 30598
rect 18696 30534 18748 30540
rect 18708 29850 18736 30534
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18420 28552 18472 28558
rect 18472 28512 18552 28540
rect 18420 28494 18472 28500
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 18524 28218 18552 28512
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 18156 27470 18184 27950
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 17880 25378 17908 26318
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26042 18368 26182
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17788 25350 17908 25378
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17512 22066 17632 22094
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 20806 17540 21966
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16592 14414 16620 14554
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16684 14074 16712 14350
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16776 12434 16804 14010
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16592 12406 16804 12434
rect 16592 12186 16620 12406
rect 16500 12170 16620 12186
rect 16868 12170 16896 13806
rect 16488 12164 16620 12170
rect 16540 12158 16620 12164
rect 16488 12106 16540 12112
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16488 11076 16540 11082
rect 16224 11036 16488 11064
rect 16488 11018 16540 11024
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16118 10024 16174 10033
rect 16118 9959 16120 9968
rect 16172 9959 16174 9968
rect 16120 9930 16172 9936
rect 16500 9042 16528 10542
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 15948 8622 16252 8650
rect 15934 8528 15990 8537
rect 15934 8463 15990 8472
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 7002 15700 7686
rect 15660 6996 15712 7002
rect 15712 6956 15884 6984
rect 15660 6938 15712 6944
rect 15856 5234 15884 6956
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15672 4554 15700 5102
rect 15856 4554 15884 5170
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15856 4146 15884 4490
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15856 3074 15884 4082
rect 15948 3534 15976 8463
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16132 7886 16160 8366
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16040 7002 16068 7686
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15856 3046 15976 3074
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15580 2746 15700 2774
rect 15672 1902 15700 2746
rect 15660 1896 15712 1902
rect 15660 1838 15712 1844
rect 15856 800 15884 2926
rect 15948 2514 15976 3046
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 16040 2310 16068 6938
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16132 2650 16160 6190
rect 16224 4162 16252 8622
rect 16592 7478 16620 12158
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16960 11898 16988 14758
rect 17052 11898 17080 18566
rect 17420 18170 17448 19450
rect 17512 18222 17540 20334
rect 17604 19242 17632 22066
rect 17592 19236 17644 19242
rect 17592 19178 17644 19184
rect 17604 18970 17632 19178
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17328 18142 17448 18170
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17130 17912 17186 17921
rect 17130 17847 17186 17856
rect 17144 17270 17172 17847
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17236 16250 17264 16458
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17222 16144 17278 16153
rect 17222 16079 17224 16088
rect 17276 16079 17278 16088
rect 17224 16050 17276 16056
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 15337 17172 15846
rect 17130 15328 17186 15337
rect 17130 15263 17186 15272
rect 17236 15162 17264 16050
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17328 14074 17356 18142
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17314 13560 17370 13569
rect 17314 13495 17316 13504
rect 17368 13495 17370 13504
rect 17316 13466 17368 13472
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11286 16712 11630
rect 16672 11280 16724 11286
rect 16672 11222 16724 11228
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16684 7342 16712 11222
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16776 10810 16804 11086
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16854 10704 16910 10713
rect 16854 10639 16910 10648
rect 16868 9994 16896 10639
rect 16960 10441 16988 11154
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16946 10432 17002 10441
rect 16946 10367 17002 10376
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 6254 16344 6734
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16408 4729 16436 7210
rect 16500 6934 16528 7210
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16500 6118 16528 6666
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16488 5636 16540 5642
rect 16592 5624 16620 6802
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16684 5642 16712 6258
rect 16540 5596 16620 5624
rect 16488 5578 16540 5584
rect 16592 4758 16620 5596
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16684 5234 16712 5578
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16684 5030 16712 5170
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16580 4752 16632 4758
rect 16394 4720 16450 4729
rect 16580 4694 16632 4700
rect 16394 4655 16450 4664
rect 16224 4134 16344 4162
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16224 800 16252 4014
rect 16316 3126 16344 4134
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16408 2310 16436 4082
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16592 800 16620 2858
rect 16776 2446 16804 9862
rect 16960 9518 16988 10367
rect 17052 10198 17080 10610
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7478 16896 7686
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16960 6798 16988 9454
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16960 5778 16988 6734
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 17144 3058 17172 13126
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17236 11121 17264 12786
rect 17328 12646 17356 13262
rect 17420 12986 17448 17478
rect 17512 16998 17540 17682
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 13870 17540 16934
rect 17604 16574 17632 18770
rect 17696 17610 17724 24142
rect 17788 19310 17816 25350
rect 17972 25140 18000 25434
rect 18432 25294 18460 28018
rect 18512 27872 18564 27878
rect 18510 27840 18512 27849
rect 18564 27840 18566 27849
rect 18510 27775 18566 27784
rect 18616 26042 18644 28698
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 18616 25498 18644 25978
rect 18708 25838 18736 29786
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18892 28762 18920 29582
rect 19076 29238 19104 35498
rect 19536 34082 19564 43726
rect 19536 34066 19748 34082
rect 19536 34060 19760 34066
rect 19536 34054 19708 34060
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19248 33856 19300 33862
rect 19248 33798 19300 33804
rect 19260 33318 19288 33798
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 19260 32570 19288 33254
rect 19444 32910 19472 33934
rect 19536 33522 19564 34054
rect 19708 34002 19760 34008
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19248 32564 19300 32570
rect 19248 32506 19300 32512
rect 19260 32026 19288 32506
rect 19444 32230 19472 32846
rect 19616 32496 19668 32502
rect 19668 32456 19748 32484
rect 19616 32438 19668 32444
rect 19720 32230 19748 32456
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19708 32224 19760 32230
rect 19708 32166 19760 32172
rect 19248 32020 19300 32026
rect 19248 31962 19300 31968
rect 19260 31754 19288 31962
rect 19444 31822 19472 32166
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19248 31748 19300 31754
rect 19248 31690 19300 31696
rect 19260 31414 19288 31690
rect 19248 31408 19300 31414
rect 19248 31350 19300 31356
rect 19260 30938 19288 31350
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19260 30666 19288 30874
rect 19444 30802 19472 31758
rect 19720 31482 19748 31826
rect 19708 31476 19760 31482
rect 19708 31418 19760 31424
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19248 30660 19300 30666
rect 19248 30602 19300 30608
rect 19260 30394 19288 30602
rect 19248 30388 19300 30394
rect 19248 30330 19300 30336
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19168 29306 19196 29446
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19064 29232 19116 29238
rect 19064 29174 19116 29180
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18800 27062 18828 28154
rect 18788 27056 18840 27062
rect 18788 26998 18840 27004
rect 18800 26518 18828 26998
rect 18984 26790 19012 28562
rect 19260 27282 19288 29990
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19352 28558 19380 29650
rect 19616 29504 19668 29510
rect 19616 29446 19668 29452
rect 19524 29028 19576 29034
rect 19444 28988 19524 29016
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19168 27254 19288 27282
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 18788 26512 18840 26518
rect 18788 26454 18840 26460
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18604 25492 18656 25498
rect 18604 25434 18656 25440
rect 18420 25288 18472 25294
rect 18418 25256 18420 25265
rect 18472 25256 18474 25265
rect 18616 25226 18644 25434
rect 18418 25191 18474 25200
rect 18604 25220 18656 25226
rect 17880 25112 18000 25140
rect 17880 24954 17908 25112
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 18328 24880 18380 24886
rect 18328 24822 18380 24828
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17880 19922 17908 24550
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23746 18368 24822
rect 18432 24818 18460 25191
rect 18604 25162 18656 25168
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18524 24206 18552 25094
rect 18616 24970 18644 25162
rect 18616 24942 18736 24970
rect 18708 24818 18736 24942
rect 18696 24812 18748 24818
rect 18748 24772 18828 24800
rect 18696 24754 18748 24760
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18248 23718 18368 23746
rect 18248 23118 18276 23718
rect 18328 23248 18380 23254
rect 18328 23190 18380 23196
rect 18420 23248 18472 23254
rect 18420 23190 18472 23196
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17788 18766 17816 19246
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17788 17678 17816 18702
rect 18340 18630 18368 23190
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17866 17912 17922 17921
rect 17922 17882 18000 17898
rect 17922 17876 18012 17882
rect 17922 17870 17960 17876
rect 17866 17847 17922 17856
rect 17960 17818 18012 17824
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17880 17610 17908 17750
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17696 16640 17724 17546
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18432 17270 18460 23190
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16726 17908 17070
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18432 16794 18460 16934
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17696 16612 17816 16640
rect 17604 16546 17724 16574
rect 17696 15366 17724 16546
rect 17788 16522 17816 16612
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17788 16046 17816 16458
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 12238 17356 12378
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17222 11112 17278 11121
rect 17222 11047 17278 11056
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17236 7546 17264 7754
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17236 4826 17264 6258
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17328 3534 17356 10406
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17420 6497 17448 7482
rect 17406 6488 17462 6497
rect 17406 6423 17462 6432
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17420 5370 17448 6190
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17512 4706 17540 13262
rect 17604 10742 17632 14486
rect 17696 11830 17724 15302
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17684 11824 17736 11830
rect 17788 11801 17816 12922
rect 17684 11766 17736 11772
rect 17774 11792 17830 11801
rect 17774 11727 17830 11736
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17788 11218 17816 11630
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17788 10130 17816 11154
rect 17880 11014 17908 15846
rect 18432 15366 18460 16730
rect 18524 16114 18552 24006
rect 18616 22098 18644 24686
rect 18800 23202 18828 24772
rect 18984 24274 19012 26726
rect 19064 24676 19116 24682
rect 19064 24618 19116 24624
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18880 24132 18932 24138
rect 18880 24074 18932 24080
rect 18892 23866 18920 24074
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18892 23497 18920 23802
rect 18878 23488 18934 23497
rect 18878 23423 18934 23432
rect 18696 23180 18748 23186
rect 18800 23174 19012 23202
rect 18696 23122 18748 23128
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18708 21434 18736 23122
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18800 22778 18828 23054
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18800 22658 18828 22714
rect 18800 22630 18920 22658
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18800 21622 18828 22510
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18616 21406 18736 21434
rect 18616 20398 18644 21406
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18708 21146 18736 21286
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 20534 18828 20742
rect 18892 20534 18920 22630
rect 18984 22574 19012 23174
rect 19076 22982 19104 24618
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19076 22778 19104 22918
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18972 22568 19024 22574
rect 18972 22510 19024 22516
rect 19076 21690 19104 22578
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18880 20528 18932 20534
rect 18880 20470 18932 20476
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18800 19718 18828 20470
rect 19168 20466 19196 27254
rect 19352 27146 19380 28494
rect 19444 27606 19472 28988
rect 19524 28970 19576 28976
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19444 27334 19472 27542
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 19260 27130 19472 27146
rect 19248 27124 19472 27130
rect 19300 27118 19472 27124
rect 19248 27066 19300 27072
rect 19444 26450 19472 27118
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19444 24818 19472 26386
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19260 20874 19288 23734
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19352 20346 19380 24550
rect 19444 24274 19472 24754
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19444 20602 19472 24210
rect 19536 22094 19564 28358
rect 19628 25974 19656 29446
rect 19708 28416 19760 28422
rect 19708 28358 19760 28364
rect 19720 28218 19748 28358
rect 19708 28212 19760 28218
rect 19708 28154 19760 28160
rect 19616 25968 19668 25974
rect 19616 25910 19668 25916
rect 19812 25294 19840 49846
rect 19996 38554 20024 53382
rect 21180 46368 21232 46374
rect 21180 46310 21232 46316
rect 21088 43716 21140 43722
rect 21088 43658 21140 43664
rect 19984 38548 20036 38554
rect 19984 38490 20036 38496
rect 20628 35556 20680 35562
rect 20628 35498 20680 35504
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 19996 33318 20024 33866
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 20536 33312 20588 33318
rect 20536 33254 20588 33260
rect 19892 33040 19944 33046
rect 19892 32982 19944 32988
rect 19904 32842 19932 32982
rect 19892 32836 19944 32842
rect 19892 32778 19944 32784
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 19904 27402 19932 31078
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 20088 30394 20116 30534
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 20548 30190 20576 33254
rect 20640 30326 20668 35498
rect 21100 34746 21128 43658
rect 21192 35834 21220 46310
rect 21364 43648 21416 43654
rect 21364 43590 21416 43596
rect 21272 42764 21324 42770
rect 21272 42706 21324 42712
rect 21180 35828 21232 35834
rect 21180 35770 21232 35776
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 21100 33930 21128 34682
rect 21088 33924 21140 33930
rect 21088 33866 21140 33872
rect 21100 33590 21128 33866
rect 21192 33862 21220 35566
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 21088 33584 21140 33590
rect 21088 33526 21140 33532
rect 21100 32502 21128 33526
rect 21088 32496 21140 32502
rect 21088 32438 21140 32444
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20812 31952 20864 31958
rect 20812 31894 20864 31900
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20536 30184 20588 30190
rect 20536 30126 20588 30132
rect 20352 30048 20404 30054
rect 20352 29990 20404 29996
rect 19984 27668 20036 27674
rect 19984 27610 20036 27616
rect 19892 27396 19944 27402
rect 19892 27338 19944 27344
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19892 25152 19944 25158
rect 19892 25094 19944 25100
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19720 23798 19748 24074
rect 19800 23860 19852 23866
rect 19800 23802 19852 23808
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19628 22778 19656 23666
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19720 23186 19748 23598
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19720 22642 19748 23122
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19536 22066 19748 22094
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19156 20324 19208 20330
rect 19352 20318 19472 20346
rect 19156 20266 19208 20272
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18708 19514 18736 19654
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18616 18086 18644 18770
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18432 14006 18460 15302
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18524 13841 18552 15846
rect 18616 15570 18644 18022
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18708 16998 18736 17818
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18510 13832 18566 13841
rect 18510 13767 18566 13776
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 17972 13326 18000 13466
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17880 10198 17908 10950
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10606 18368 12786
rect 18432 12481 18460 13466
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18418 12472 18474 12481
rect 18418 12407 18474 12416
rect 18524 12345 18552 12854
rect 18510 12336 18566 12345
rect 18510 12271 18566 12280
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11898 18460 12038
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 18326 10160 18382 10169
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17960 10124 18012 10130
rect 18326 10095 18328 10104
rect 17960 10066 18012 10072
rect 18380 10095 18382 10104
rect 18328 10066 18380 10072
rect 17972 9908 18000 10066
rect 17880 9880 18000 9908
rect 18236 9920 18288 9926
rect 17880 9722 17908 9880
rect 18288 9880 18368 9908
rect 18236 9862 18288 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 9042 18276 9454
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17604 8430 17632 8502
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17604 5794 17632 8230
rect 17696 7993 17724 8910
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18248 8401 18276 8434
rect 18234 8392 18290 8401
rect 18234 8327 18290 8336
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17682 7984 17738 7993
rect 17682 7919 17738 7928
rect 17880 7546 17908 8026
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17696 6730 17724 7278
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17696 5914 17724 6666
rect 17788 5914 17816 7142
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17880 6440 17908 6666
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17880 6412 18000 6440
rect 17972 6322 18000 6412
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17774 5808 17830 5817
rect 17604 5766 17724 5794
rect 17512 4678 17632 4706
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17316 3120 17368 3126
rect 17236 3080 17316 3108
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17236 2774 17264 3080
rect 17316 3062 17368 3068
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 16960 2746 17264 2774
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16960 800 16988 2746
rect 17328 2514 17356 2790
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17420 2122 17448 4014
rect 17512 3194 17540 4558
rect 17604 4146 17632 4678
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17696 2938 17724 5766
rect 17774 5743 17830 5752
rect 17788 5234 17816 5743
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17880 4486 17908 6190
rect 18340 5778 18368 9880
rect 18432 7274 18460 10406
rect 18510 10296 18566 10305
rect 18510 10231 18566 10240
rect 18524 9722 18552 10231
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18420 7268 18472 7274
rect 18420 7210 18472 7216
rect 18524 7206 18552 8366
rect 18616 7886 18644 14962
rect 18708 13190 18736 15642
rect 18800 15094 18828 19110
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18892 18086 18920 18294
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18892 17882 18920 18022
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18892 13870 18920 17070
rect 18984 14890 19012 18634
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18892 12782 18920 13806
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18696 12640 18748 12646
rect 18748 12588 18828 12594
rect 18696 12582 18828 12588
rect 18708 12566 18828 12582
rect 18800 12442 18828 12566
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18786 12336 18842 12345
rect 18786 12271 18842 12280
rect 18800 12238 18828 12271
rect 18788 12232 18840 12238
rect 18694 12200 18750 12209
rect 18788 12174 18840 12180
rect 18694 12135 18696 12144
rect 18748 12135 18750 12144
rect 18696 12106 18748 12112
rect 18800 10538 18828 12174
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18892 10441 18920 12038
rect 18878 10432 18934 10441
rect 18878 10367 18934 10376
rect 18694 10160 18750 10169
rect 18694 10095 18750 10104
rect 18788 10124 18840 10130
rect 18708 9926 18736 10095
rect 18788 10066 18840 10072
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18694 9752 18750 9761
rect 18694 9687 18750 9696
rect 18708 9382 18736 9687
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 8566 18736 9318
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18602 7168 18658 7177
rect 18524 5817 18552 7142
rect 18602 7103 18658 7112
rect 18510 5808 18566 5817
rect 18328 5772 18380 5778
rect 18510 5743 18566 5752
rect 18328 5714 18380 5720
rect 18418 5672 18474 5681
rect 18418 5607 18474 5616
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17788 2961 17816 3946
rect 18340 3482 18368 5510
rect 18248 3454 18368 3482
rect 18248 3398 18276 3454
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17328 2094 17448 2122
rect 17604 2910 17724 2938
rect 17774 2952 17830 2961
rect 17604 2106 17632 2910
rect 17774 2887 17830 2896
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17592 2100 17644 2106
rect 17328 800 17356 2094
rect 17592 2042 17644 2048
rect 17696 800 17724 2790
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 3334
rect 18432 3058 18460 5607
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18524 2122 18552 4082
rect 18616 3670 18644 7103
rect 18708 4010 18736 8366
rect 18800 7206 18828 10066
rect 18892 10062 18920 10367
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18984 9908 19012 13670
rect 19076 10713 19104 20198
rect 19168 19378 19196 20266
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19168 12306 19196 12786
rect 19260 12374 19288 17546
rect 19352 14550 19380 20198
rect 19444 17746 19472 20318
rect 19536 19514 19564 21286
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 16114 19472 16390
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19444 13326 19472 16050
rect 19628 15434 19656 20946
rect 19720 19854 19748 22066
rect 19812 20942 19840 23802
rect 19904 23633 19932 25094
rect 19996 23730 20024 27610
rect 20076 27328 20128 27334
rect 20076 27270 20128 27276
rect 20088 26790 20116 27270
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19890 23624 19946 23633
rect 19890 23559 19946 23568
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19904 23118 19932 23462
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19996 21486 20024 22510
rect 20088 21894 20116 25162
rect 20260 23520 20312 23526
rect 20260 23462 20312 23468
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20088 21690 20116 21830
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20180 21622 20208 21830
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 19984 21480 20036 21486
rect 19904 21428 19984 21434
rect 19904 21422 20036 21428
rect 19904 21406 20024 21422
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19904 19786 19932 21406
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19812 17746 19840 19722
rect 19904 19378 19932 19722
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19522 15192 19578 15201
rect 19522 15127 19578 15136
rect 19536 14006 19564 15127
rect 19720 14550 19748 17614
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19812 16182 19840 17546
rect 19800 16176 19852 16182
rect 19800 16118 19852 16124
rect 19708 14544 19760 14550
rect 19708 14486 19760 14492
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19628 13938 19656 14214
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19720 12714 19748 13942
rect 19708 12708 19760 12714
rect 19708 12650 19760 12656
rect 19812 12434 19840 14214
rect 19720 12406 19840 12434
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19260 12186 19288 12310
rect 19168 12158 19288 12186
rect 19432 12164 19484 12170
rect 19168 11150 19196 12158
rect 19432 12106 19484 12112
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19444 12050 19472 12106
rect 19156 11144 19208 11150
rect 19260 11121 19288 12038
rect 19444 12022 19656 12050
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19156 11086 19208 11092
rect 19246 11112 19302 11121
rect 19246 11047 19302 11056
rect 19062 10704 19118 10713
rect 19062 10639 19118 10648
rect 19352 10606 19380 11494
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19444 10169 19472 11154
rect 19536 10985 19564 11222
rect 19522 10976 19578 10985
rect 19522 10911 19578 10920
rect 19522 10840 19578 10849
rect 19522 10775 19578 10784
rect 19536 10742 19564 10775
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19430 10160 19486 10169
rect 19536 10130 19564 10406
rect 19430 10095 19486 10104
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19156 9920 19208 9926
rect 18984 9880 19104 9908
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18892 9353 18920 9454
rect 18878 9344 18934 9353
rect 18878 9279 18934 9288
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18800 5352 18828 6734
rect 18892 5778 18920 7278
rect 18984 7177 19012 9658
rect 19076 9382 19104 9880
rect 19156 9862 19208 9868
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 9178 19104 9318
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19168 8090 19196 9862
rect 19352 9674 19380 9862
rect 19524 9716 19576 9722
rect 19248 9648 19300 9654
rect 19352 9646 19472 9674
rect 19524 9658 19576 9664
rect 19248 9590 19300 9596
rect 19260 9489 19288 9590
rect 19246 9480 19302 9489
rect 19444 9466 19472 9646
rect 19246 9415 19302 9424
rect 19352 9438 19472 9466
rect 19248 9376 19300 9382
rect 19246 9344 19248 9353
rect 19300 9344 19302 9353
rect 19246 9279 19302 9288
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19260 7342 19288 8978
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 18970 7168 19026 7177
rect 18970 7103 19026 7112
rect 18970 7032 19026 7041
rect 19352 6984 19380 9438
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9110 19472 9318
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19536 8974 19564 9658
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 18970 6967 19026 6976
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18880 5364 18932 5370
rect 18800 5324 18880 5352
rect 18880 5306 18932 5312
rect 18892 5030 18920 5306
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18892 4826 18920 4966
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18708 2650 18736 3538
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18432 2094 18552 2122
rect 18432 800 18460 2094
rect 18892 1714 18920 3606
rect 18984 3058 19012 6967
rect 19076 6956 19380 6984
rect 19076 4146 19104 6956
rect 19444 6882 19472 8842
rect 19522 8256 19578 8265
rect 19522 8191 19578 8200
rect 19536 7886 19564 8191
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19628 7698 19656 12022
rect 19720 8498 19748 12406
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11694 19840 12038
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 19536 7670 19656 7698
rect 19536 6934 19564 7670
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19352 6854 19472 6882
rect 19524 6928 19576 6934
rect 19524 6870 19576 6876
rect 19352 6662 19380 6854
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19352 6458 19380 6598
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 19076 3602 19104 3878
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18800 1686 18920 1714
rect 18800 800 18828 1686
rect 19168 800 19196 5714
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19260 2378 19288 5578
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 5098 19380 5510
rect 19444 5302 19472 6598
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19628 5234 19656 7482
rect 19616 5228 19668 5234
rect 19536 5188 19616 5216
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19430 4720 19486 4729
rect 19536 4690 19564 5188
rect 19616 5170 19668 5176
rect 19616 5092 19668 5098
rect 19616 5034 19668 5040
rect 19628 4729 19656 5034
rect 19614 4720 19670 4729
rect 19430 4655 19486 4664
rect 19524 4684 19576 4690
rect 19444 3534 19472 4655
rect 19614 4655 19670 4664
rect 19524 4626 19576 4632
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19536 3534 19564 4490
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19248 2372 19300 2378
rect 19248 2314 19300 2320
rect 19444 2106 19472 2382
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19536 800 19564 3334
rect 19720 2774 19748 7754
rect 19812 7154 19840 11494
rect 19904 9994 19932 18566
rect 19996 18290 20024 19246
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19996 16794 20024 17138
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20088 15162 20116 21014
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20180 16590 20208 19858
rect 20272 17610 20300 23462
rect 20364 20466 20392 29990
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20548 29306 20576 29446
rect 20536 29300 20588 29306
rect 20536 29242 20588 29248
rect 20548 29034 20576 29242
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20640 28150 20668 28494
rect 20824 28490 20852 31894
rect 20916 29102 20944 32166
rect 21100 31822 21128 32438
rect 21192 32366 21220 33798
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 30666 21036 31622
rect 20996 30660 21048 30666
rect 20996 30602 21048 30608
rect 20904 29096 20956 29102
rect 20904 29038 20956 29044
rect 20916 28490 20944 29038
rect 21008 28626 21036 30602
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 20904 28484 20956 28490
rect 20904 28426 20956 28432
rect 20628 28144 20680 28150
rect 20628 28086 20680 28092
rect 20536 27940 20588 27946
rect 20536 27882 20588 27888
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20456 24410 20484 24686
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20456 23186 20484 24346
rect 20548 24070 20576 27882
rect 20996 27872 21048 27878
rect 20996 27814 21048 27820
rect 21008 26586 21036 27814
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 20996 26444 21048 26450
rect 20996 26386 21048 26392
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20824 23186 20852 23666
rect 21008 23662 21036 26386
rect 21100 26314 21128 26726
rect 21088 26308 21140 26314
rect 21088 26250 21140 26256
rect 21100 25498 21128 26250
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 21100 24818 21128 25434
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 21100 24138 21128 24754
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20364 17338 20392 19314
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20180 16182 20208 16526
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20180 15570 20208 16118
rect 20548 16046 20576 22102
rect 20732 19514 20760 22374
rect 20996 21412 21048 21418
rect 20996 21354 21048 21360
rect 21008 20942 21036 21354
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21192 20534 21220 23530
rect 21180 20528 21232 20534
rect 21180 20470 21232 20476
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21008 16794 21036 16934
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21008 16522 21036 16730
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19996 11830 20024 14962
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20180 12442 20208 14554
rect 20258 14512 20314 14521
rect 20258 14447 20314 14456
rect 20272 14414 20300 14447
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20088 11830 20116 12378
rect 20180 12238 20208 12378
rect 20272 12306 20300 13194
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19996 11150 20024 11630
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20180 11354 20208 11562
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19892 9988 19944 9994
rect 19892 9930 19944 9936
rect 19996 9926 20024 10950
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 19984 9920 20036 9926
rect 20088 9908 20116 10678
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20180 10033 20208 10542
rect 20166 10024 20222 10033
rect 20166 9959 20222 9968
rect 20168 9920 20220 9926
rect 20088 9880 20168 9908
rect 19984 9862 20036 9868
rect 20168 9862 20220 9868
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 7410 19932 9318
rect 19996 8362 20024 9862
rect 20180 9722 20208 9862
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19812 7126 20024 7154
rect 19892 6928 19944 6934
rect 19892 6870 19944 6876
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19812 5846 19840 6598
rect 19800 5840 19852 5846
rect 19800 5782 19852 5788
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19628 2746 19748 2774
rect 19628 2446 19656 2746
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19812 2292 19840 4762
rect 19904 3058 19932 6870
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19904 2514 19932 2790
rect 19996 2650 20024 7126
rect 20088 3738 20116 9522
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 20180 4214 20208 9386
rect 20272 9042 20300 12242
rect 20364 12102 20392 15302
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20364 11082 20392 11562
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20456 10266 20484 14486
rect 20548 12782 20576 15982
rect 20640 15366 20668 16458
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15706 20760 15846
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20640 14958 20668 15302
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20732 12434 20760 13330
rect 20824 12714 20852 16050
rect 21008 15434 21036 16458
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 21100 13841 21128 18022
rect 21086 13832 21142 13841
rect 21086 13767 21142 13776
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20732 12406 20852 12434
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20364 9042 20392 10134
rect 20456 9926 20484 10202
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20272 7546 20300 8978
rect 20444 7880 20496 7886
rect 20442 7848 20444 7857
rect 20496 7848 20498 7857
rect 20442 7783 20498 7792
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20364 6866 20392 7346
rect 20456 7002 20484 7346
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20272 5914 20300 6394
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 20364 4010 20392 6258
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20260 4004 20312 4010
rect 20260 3946 20312 3952
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20272 3738 20300 3946
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 20456 2292 20484 5782
rect 20548 4026 20576 11698
rect 20640 11558 20668 11766
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20640 11150 20668 11290
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20732 10606 20760 12106
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20718 10160 20774 10169
rect 20718 10095 20774 10104
rect 20732 9994 20760 10095
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20732 9518 20760 9930
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 6769 20668 7822
rect 20732 7342 20760 8026
rect 20720 7336 20772 7342
rect 20718 7304 20720 7313
rect 20772 7304 20774 7313
rect 20718 7239 20774 7248
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20626 6760 20682 6769
rect 20626 6695 20682 6704
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20640 5642 20668 6190
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 20732 4078 20760 7142
rect 20824 6798 20852 12406
rect 20916 11694 20944 12854
rect 21008 12850 21036 13126
rect 21100 12986 21128 13466
rect 21192 12986 21220 19178
rect 21284 13258 21312 42706
rect 21376 33114 21404 43590
rect 21468 41614 21496 53450
rect 22296 53038 22324 53518
rect 23308 53242 23336 53586
rect 23400 53582 23428 56063
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 23400 53242 23428 53518
rect 23940 53440 23992 53446
rect 23940 53382 23992 53388
rect 23296 53236 23348 53242
rect 23296 53178 23348 53184
rect 23388 53236 23440 53242
rect 23388 53178 23440 53184
rect 22284 53032 22336 53038
rect 22284 52974 22336 52980
rect 23664 52896 23716 52902
rect 23664 52838 23716 52844
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 23388 50176 23440 50182
rect 23388 50118 23440 50124
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 23400 48142 23428 50118
rect 23388 48136 23440 48142
rect 23388 48078 23440 48084
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 21732 42016 21784 42022
rect 21732 41958 21784 41964
rect 21456 41608 21508 41614
rect 21456 41550 21508 41556
rect 21364 33108 21416 33114
rect 21364 33050 21416 33056
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21652 26450 21680 27270
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21548 25696 21600 25702
rect 21548 25638 21600 25644
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21456 22704 21508 22710
rect 21456 22646 21508 22652
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21376 16250 21404 21898
rect 21468 20806 21496 22646
rect 21560 22642 21588 25638
rect 21652 23118 21680 25638
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21468 20602 21496 20742
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21468 15552 21496 19178
rect 21376 15524 21496 15552
rect 21376 13938 21404 15524
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21468 15026 21496 15370
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14362 21496 14758
rect 21560 14482 21588 20266
rect 21640 19984 21692 19990
rect 21640 19926 21692 19932
rect 21652 19310 21680 19926
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21652 15502 21680 18838
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21468 14334 21588 14362
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 6390 20944 6734
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 21008 5710 21036 11154
rect 21284 11082 21312 12922
rect 21376 12753 21404 13262
rect 21468 12986 21496 13398
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21560 12866 21588 14334
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21468 12838 21588 12866
rect 21362 12744 21418 12753
rect 21362 12679 21418 12688
rect 21362 11928 21418 11937
rect 21362 11863 21364 11872
rect 21416 11863 21418 11872
rect 21364 11834 21416 11840
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21468 11014 21496 12838
rect 21652 12434 21680 13806
rect 21744 12442 21772 41958
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23296 40180 23348 40186
rect 23296 40122 23348 40128
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 22020 34950 22048 35634
rect 22008 34944 22060 34950
rect 22008 34886 22060 34892
rect 21916 33584 21968 33590
rect 21916 33526 21968 33532
rect 21928 33114 21956 33526
rect 21916 33108 21968 33114
rect 21916 33050 21968 33056
rect 21824 33040 21876 33046
rect 21824 32982 21876 32988
rect 21836 32434 21864 32982
rect 21928 32842 21956 33050
rect 21916 32836 21968 32842
rect 21916 32778 21968 32784
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21836 32230 21864 32370
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21836 29034 21864 32166
rect 22020 31686 22048 34886
rect 22112 31686 22140 35702
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 22192 34944 22244 34950
rect 22192 34886 22244 34892
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 21916 31340 21968 31346
rect 21916 31282 21968 31288
rect 21928 31142 21956 31282
rect 22020 31210 22048 31622
rect 22008 31204 22060 31210
rect 22008 31146 22060 31152
rect 22204 31142 22232 34886
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22296 33590 22324 34002
rect 22376 33924 22428 33930
rect 22376 33866 22428 33872
rect 22388 33590 22416 33866
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 22296 32978 22324 33526
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22388 33114 22416 33390
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22296 32502 22324 32914
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22296 31346 22324 32438
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22376 31272 22428 31278
rect 22376 31214 22428 31220
rect 22284 31204 22336 31210
rect 22284 31146 22336 31152
rect 21916 31136 21968 31142
rect 22192 31136 22244 31142
rect 21968 31084 22048 31090
rect 21916 31078 22048 31084
rect 22192 31078 22244 31084
rect 21928 31062 22048 31078
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21836 28082 21864 28970
rect 21916 28688 21968 28694
rect 21916 28630 21968 28636
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21928 23866 21956 28630
rect 22020 26518 22048 31062
rect 22296 28422 22324 31146
rect 22388 30666 22416 31214
rect 22376 30660 22428 30666
rect 22376 30602 22428 30608
rect 22480 30326 22508 34886
rect 22572 33658 22600 35566
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22560 33652 22612 33658
rect 22560 33594 22612 33600
rect 22756 33114 22784 35090
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 23020 34196 23072 34202
rect 23020 34138 23072 34144
rect 23032 33454 23060 34138
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 23216 33658 23244 33798
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 23020 33448 23072 33454
rect 22848 33396 23020 33402
rect 22848 33390 23072 33396
rect 22848 33374 23060 33390
rect 22744 33108 22796 33114
rect 22744 33050 22796 33056
rect 22744 31952 22796 31958
rect 22744 31894 22796 31900
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 26586 22140 26862
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22008 26512 22060 26518
rect 22008 26454 22060 26460
rect 22020 25838 22048 26454
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 22112 23066 22140 25638
rect 22204 24818 22232 26386
rect 22296 26246 22324 28358
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 22388 27402 22416 27814
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 22284 26240 22336 26246
rect 22284 26182 22336 26188
rect 22296 26042 22324 26182
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22296 24274 22324 24890
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22204 23730 22232 24210
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22020 23038 22140 23066
rect 22020 22522 22048 23038
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 22642 22140 22918
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22020 22494 22140 22522
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21836 16998 21864 19110
rect 21928 18986 21956 21286
rect 22020 21010 22048 21490
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22112 19530 22140 22494
rect 22204 22098 22232 23666
rect 22296 23526 22324 24006
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 22296 21962 22324 23462
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 21418 22324 21898
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 20058 22232 20402
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22112 19502 22324 19530
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 21928 18958 22048 18986
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21928 16114 21956 16390
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15978 21956 16050
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 22020 15450 22048 18958
rect 22204 18766 22232 19382
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22112 18290 22140 18566
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22296 17921 22324 19502
rect 22388 18358 22416 26726
rect 22480 26042 22508 29446
rect 22572 28150 22600 31622
rect 22652 31408 22704 31414
rect 22652 31350 22704 31356
rect 22664 30938 22692 31350
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22572 26926 22600 27950
rect 22664 26994 22692 30602
rect 22756 27130 22784 31894
rect 22848 30190 22876 33374
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23308 31890 23336 40122
rect 23676 39982 23704 52838
rect 23848 52624 23900 52630
rect 23848 52566 23900 52572
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23860 35894 23888 52566
rect 23492 35866 23888 35894
rect 23492 32774 23520 35866
rect 23572 33652 23624 33658
rect 23572 33594 23624 33600
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 23296 31884 23348 31890
rect 23296 31826 23348 31832
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23032 31414 23060 31758
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 23480 31136 23532 31142
rect 23480 31078 23532 31084
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 23492 30326 23520 31078
rect 23480 30320 23532 30326
rect 23480 30262 23532 30268
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22848 27554 22876 29786
rect 23308 29186 23336 30126
rect 23308 29158 23428 29186
rect 23400 29102 23428 29158
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23204 28688 23256 28694
rect 23204 28630 23256 28636
rect 23216 28422 23244 28630
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23400 28150 23428 29038
rect 23492 28370 23520 30262
rect 23584 28558 23612 33594
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23860 32842 23888 33254
rect 23848 32836 23900 32842
rect 23848 32778 23900 32784
rect 23860 31754 23888 32778
rect 23768 31726 23888 31754
rect 23768 30138 23796 31726
rect 23952 30190 23980 53382
rect 24504 52698 24532 56200
rect 25318 55448 25374 55457
rect 25318 55383 25374 55392
rect 24766 54632 24822 54641
rect 24766 54567 24822 54576
rect 24676 53984 24728 53990
rect 24676 53926 24728 53932
rect 24688 53582 24716 53926
rect 24676 53576 24728 53582
rect 24676 53518 24728 53524
rect 24584 53440 24636 53446
rect 24584 53382 24636 53388
rect 24492 52692 24544 52698
rect 24492 52634 24544 52640
rect 24504 52494 24532 52634
rect 24492 52488 24544 52494
rect 24492 52430 24544 52436
rect 24596 52018 24624 53382
rect 24780 53242 24808 54567
rect 24858 53816 24914 53825
rect 24858 53751 24914 53760
rect 24768 53236 24820 53242
rect 24768 53178 24820 53184
rect 24872 53038 24900 53751
rect 25332 53242 25360 55383
rect 25884 54194 25912 56200
rect 25872 54188 25924 54194
rect 25872 54130 25924 54136
rect 25320 53236 25372 53242
rect 25320 53178 25372 53184
rect 24860 53032 24912 53038
rect 24860 52974 24912 52980
rect 25502 53000 25558 53009
rect 25502 52935 25504 52944
rect 25556 52935 25558 52944
rect 25504 52906 25556 52912
rect 24676 52896 24728 52902
rect 24676 52838 24728 52844
rect 24584 52012 24636 52018
rect 24584 51954 24636 51960
rect 24584 51808 24636 51814
rect 24584 51750 24636 51756
rect 24596 50318 24624 51750
rect 24584 50312 24636 50318
rect 24584 50254 24636 50260
rect 24216 49836 24268 49842
rect 24216 49778 24268 49784
rect 24228 49434 24256 49778
rect 24216 49428 24268 49434
rect 24216 49370 24268 49376
rect 24032 48000 24084 48006
rect 24032 47942 24084 47948
rect 24044 43858 24072 47942
rect 24688 45554 24716 52838
rect 24952 52420 25004 52426
rect 24952 52362 25004 52368
rect 24964 52193 24992 52362
rect 24950 52184 25006 52193
rect 24950 52119 24952 52128
rect 25004 52119 25006 52128
rect 24952 52090 25004 52096
rect 25516 52018 25544 52906
rect 25964 52488 26016 52494
rect 25964 52430 26016 52436
rect 25504 52012 25556 52018
rect 25504 51954 25556 51960
rect 25228 51808 25280 51814
rect 25228 51750 25280 51756
rect 24950 51368 25006 51377
rect 24950 51303 24952 51312
rect 25004 51303 25006 51312
rect 24952 51274 25004 51280
rect 25044 50924 25096 50930
rect 25044 50866 25096 50872
rect 24952 50720 25004 50726
rect 24952 50662 25004 50668
rect 24766 49736 24822 49745
rect 24766 49671 24822 49680
rect 24780 49434 24808 49671
rect 24768 49428 24820 49434
rect 24768 49370 24820 49376
rect 24860 49224 24912 49230
rect 24860 49166 24912 49172
rect 24872 48929 24900 49166
rect 24858 48920 24914 48929
rect 24858 48855 24860 48864
rect 24912 48855 24914 48864
rect 24860 48826 24912 48832
rect 24860 48136 24912 48142
rect 24858 48104 24860 48113
rect 24912 48104 24914 48113
rect 24858 48039 24914 48048
rect 24872 47802 24900 48039
rect 24860 47796 24912 47802
rect 24860 47738 24912 47744
rect 24504 45526 24716 45554
rect 24032 43852 24084 43858
rect 24032 43794 24084 43800
rect 24504 42090 24532 45526
rect 24964 45014 24992 50662
rect 25056 50561 25084 50866
rect 25042 50552 25098 50561
rect 25042 50487 25098 50496
rect 25136 49088 25188 49094
rect 25136 49030 25188 49036
rect 25148 48822 25176 49030
rect 25136 48816 25188 48822
rect 25136 48758 25188 48764
rect 25136 48000 25188 48006
rect 25136 47942 25188 47948
rect 25148 47734 25176 47942
rect 25136 47728 25188 47734
rect 25136 47670 25188 47676
rect 25240 47598 25268 51750
rect 25780 51332 25832 51338
rect 25780 51274 25832 51280
rect 25228 47592 25280 47598
rect 25228 47534 25280 47540
rect 25688 47524 25740 47530
rect 25688 47466 25740 47472
rect 25318 47288 25374 47297
rect 25318 47223 25374 47232
rect 25332 47054 25360 47223
rect 25320 47048 25372 47054
rect 25320 46990 25372 46996
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25332 46481 25360 46514
rect 25318 46472 25374 46481
rect 25318 46407 25374 46416
rect 25320 45960 25372 45966
rect 25320 45902 25372 45908
rect 25044 45824 25096 45830
rect 25044 45766 25096 45772
rect 24952 45008 25004 45014
rect 24952 44950 25004 44956
rect 24676 44396 24728 44402
rect 24676 44338 24728 44344
rect 24688 44033 24716 44338
rect 24674 44024 24730 44033
rect 24674 43959 24730 43968
rect 24860 43648 24912 43654
rect 24860 43590 24912 43596
rect 24872 42838 24900 43590
rect 24952 43308 25004 43314
rect 24952 43250 25004 43256
rect 24964 43217 24992 43250
rect 24950 43208 25006 43217
rect 24950 43143 25006 43152
rect 24860 42832 24912 42838
rect 24860 42774 24912 42780
rect 24860 42696 24912 42702
rect 24860 42638 24912 42644
rect 24872 42401 24900 42638
rect 24858 42392 24914 42401
rect 24858 42327 24860 42336
rect 24912 42327 24914 42336
rect 24860 42298 24912 42304
rect 24492 42084 24544 42090
rect 24492 42026 24544 42032
rect 24860 41608 24912 41614
rect 24858 41576 24860 41585
rect 24912 41576 24914 41585
rect 24780 41534 24858 41562
rect 24780 41274 24808 41534
rect 24858 41511 24914 41520
rect 24768 41268 24820 41274
rect 24768 41210 24820 41216
rect 24860 40928 24912 40934
rect 24860 40870 24912 40876
rect 24124 39296 24176 39302
rect 24124 39238 24176 39244
rect 24032 32496 24084 32502
rect 24032 32438 24084 32444
rect 24044 32026 24072 32438
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 24044 31414 24072 31962
rect 24136 31958 24164 39238
rect 24872 38865 24900 40870
rect 25056 40746 25084 45766
rect 25332 45665 25360 45902
rect 25318 45656 25374 45665
rect 25318 45591 25374 45600
rect 25412 45484 25464 45490
rect 25412 45426 25464 45432
rect 25228 45280 25280 45286
rect 25228 45222 25280 45228
rect 25136 42560 25188 42566
rect 25136 42502 25188 42508
rect 25148 42294 25176 42502
rect 25136 42288 25188 42294
rect 25136 42230 25188 42236
rect 25056 40718 25176 40746
rect 24858 38856 24914 38865
rect 24858 38791 24914 38800
rect 24768 38752 24820 38758
rect 24768 38694 24820 38700
rect 25044 38752 25096 38758
rect 25044 38694 25096 38700
rect 24780 38321 24808 38694
rect 24766 38312 24822 38321
rect 24766 38247 24822 38256
rect 24860 37868 24912 37874
rect 24860 37810 24912 37816
rect 24872 37505 24900 37810
rect 24858 37496 24914 37505
rect 24858 37431 24914 37440
rect 24952 36780 25004 36786
rect 24952 36722 25004 36728
rect 24964 36689 24992 36722
rect 24950 36680 25006 36689
rect 24950 36615 25006 36624
rect 24768 36168 24820 36174
rect 24768 36110 24820 36116
rect 24676 36032 24728 36038
rect 24676 35974 24728 35980
rect 24688 35698 24716 35974
rect 24780 35873 24808 36110
rect 24766 35864 24822 35873
rect 24766 35799 24822 35808
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24216 33856 24268 33862
rect 24216 33798 24268 33804
rect 24124 31952 24176 31958
rect 24124 31894 24176 31900
rect 24032 31408 24084 31414
rect 24032 31350 24084 31356
rect 24044 30598 24072 31350
rect 24032 30592 24084 30598
rect 24032 30534 24084 30540
rect 24044 30326 24072 30534
rect 24032 30320 24084 30326
rect 24032 30262 24084 30268
rect 23940 30184 23992 30190
rect 23768 30110 23888 30138
rect 23940 30126 23992 30132
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23768 29782 23796 29990
rect 23756 29776 23808 29782
rect 23756 29718 23808 29724
rect 23860 29306 23888 30110
rect 24044 29594 24072 30262
rect 23952 29566 24072 29594
rect 23848 29300 23900 29306
rect 23848 29242 23900 29248
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23768 28762 23796 29038
rect 23756 28756 23808 28762
rect 23756 28698 23808 28704
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23492 28342 23612 28370
rect 23388 28144 23440 28150
rect 23388 28086 23440 28092
rect 23480 28144 23532 28150
rect 23480 28086 23532 28092
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22848 27526 22968 27554
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22560 26920 22612 26926
rect 22940 26874 22968 27526
rect 22560 26862 22612 26868
rect 22848 26846 22968 26874
rect 22560 26512 22612 26518
rect 22560 26454 22612 26460
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22468 24880 22520 24886
rect 22468 24822 22520 24828
rect 22480 21554 22508 24822
rect 22572 21690 22600 26454
rect 22848 26314 22876 26846
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 26042 23060 26182
rect 23020 26036 23072 26042
rect 23020 25978 23072 25984
rect 22744 25832 22796 25838
rect 22744 25774 22796 25780
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22664 24410 22692 24550
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22664 23730 22692 24210
rect 22756 23798 22784 25774
rect 22848 25498 22876 25774
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 23308 24750 23336 27814
rect 23400 27538 23428 28086
rect 23492 27606 23520 28086
rect 23480 27600 23532 27606
rect 23480 27542 23532 27548
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23400 26926 23428 27474
rect 23584 27062 23612 28342
rect 23676 27674 23704 28562
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 23664 27396 23716 27402
rect 23664 27338 23716 27344
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 23400 24682 23428 26862
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23492 25498 23520 25842
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 23676 24834 23704 27338
rect 23492 24818 23704 24834
rect 23480 24812 23704 24818
rect 23532 24806 23704 24812
rect 23480 24754 23532 24760
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 23388 24676 23440 24682
rect 23388 24618 23440 24624
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22848 23662 22876 24618
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23204 23792 23256 23798
rect 23256 23740 23336 23746
rect 23204 23734 23336 23740
rect 23216 23718 23336 23734
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22466 21448 22522 21457
rect 22466 21383 22468 21392
rect 22520 21383 22522 21392
rect 22468 21354 22520 21360
rect 22480 20262 22508 21354
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19786 22508 20198
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22282 17912 22338 17921
rect 22282 17847 22338 17856
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 21836 15422 22048 15450
rect 21836 14414 21864 15422
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21560 12406 21680 12434
rect 21732 12436 21784 12442
rect 21456 11008 21508 11014
rect 21178 10976 21234 10985
rect 21456 10950 21508 10956
rect 21178 10911 21234 10920
rect 21192 10742 21220 10911
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 21180 10736 21232 10742
rect 21180 10678 21232 10684
rect 21100 9722 21128 10678
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21284 10266 21312 10542
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 21192 9178 21220 9454
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21088 7268 21140 7274
rect 21088 7210 21140 7216
rect 21100 6662 21128 7210
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20904 5092 20956 5098
rect 20824 5052 20904 5080
rect 20720 4072 20772 4078
rect 20548 3998 20668 4026
rect 20720 4014 20772 4020
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20640 3890 20668 3998
rect 20548 2446 20576 3878
rect 20640 3862 20760 3890
rect 20732 3534 20760 3862
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 19812 2264 19932 2292
rect 20456 2264 20668 2292
rect 19904 800 19932 2264
rect 20260 1284 20312 1290
rect 20260 1226 20312 1232
rect 20272 800 20300 1226
rect 20640 800 20668 2264
rect 20824 1290 20852 5052
rect 20904 5034 20956 5040
rect 21100 4486 21128 6598
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20916 3194 20944 4082
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21192 2774 21220 8774
rect 21272 7948 21324 7954
rect 21376 7936 21404 10474
rect 21560 9110 21588 12406
rect 21732 12378 21784 12384
rect 21744 11830 21772 12378
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21836 11286 21864 14214
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 21928 11218 21956 15302
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 12986 22048 14962
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 22112 12918 22140 14418
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22020 12730 22048 12786
rect 22020 12702 22140 12730
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22020 11898 22048 12242
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11286 22048 11494
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22020 10418 22048 10746
rect 22112 10418 22140 12702
rect 22020 10390 22140 10418
rect 21824 10192 21876 10198
rect 21824 10134 21876 10140
rect 21836 9926 21864 10134
rect 21824 9920 21876 9926
rect 21638 9888 21694 9897
rect 22100 9920 22152 9926
rect 21824 9862 21876 9868
rect 22020 9880 22100 9908
rect 21638 9823 21694 9832
rect 21652 9382 21680 9823
rect 22020 9722 22048 9880
rect 22100 9862 22152 9868
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 22008 9716 22060 9722
rect 22204 9704 22232 17546
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22296 15570 22324 16118
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22284 13796 22336 13802
rect 22284 13738 22336 13744
rect 22296 11626 22324 13738
rect 22388 13190 22416 16934
rect 22572 16726 22600 20334
rect 22756 19310 22784 21626
rect 22848 20602 22876 23054
rect 23308 22658 23336 23718
rect 23400 22778 23428 24278
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23662 23612 24006
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23308 22630 23428 22658
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23020 22092 23072 22098
rect 23020 22034 23072 22040
rect 23032 21554 23060 22034
rect 23124 21690 23152 22170
rect 23204 22024 23256 22030
rect 23308 22001 23336 22510
rect 23400 22234 23428 22630
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23204 21966 23256 21972
rect 23294 21992 23350 22001
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23216 21622 23244 21966
rect 23294 21927 23350 21936
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22756 17338 22784 18022
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22848 17218 22876 17478
rect 22756 17190 22876 17218
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22284 11620 22336 11626
rect 22284 11562 22336 11568
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22296 11082 22324 11222
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22388 10130 22416 12582
rect 22480 11529 22508 14486
rect 22572 13870 22600 16526
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22664 15570 22692 15846
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22664 14006 22692 15370
rect 22652 14000 22704 14006
rect 22652 13942 22704 13948
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22664 12782 22692 13806
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22466 11520 22522 11529
rect 22466 11455 22522 11464
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22282 10024 22338 10033
rect 22282 9959 22338 9968
rect 22296 9722 22324 9959
rect 22008 9658 22060 9664
rect 22112 9676 22232 9704
rect 22284 9716 22336 9722
rect 21836 9602 21864 9658
rect 22112 9602 22140 9676
rect 22284 9658 22336 9664
rect 21836 9574 21956 9602
rect 21928 9518 21956 9574
rect 22020 9574 22140 9602
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21324 7908 21404 7936
rect 21272 7890 21324 7896
rect 21284 6934 21312 7890
rect 21456 7812 21508 7818
rect 21456 7754 21508 7760
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21376 7342 21404 7686
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 21284 5710 21312 6326
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21376 5370 21404 7142
rect 21468 7002 21496 7754
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21284 4826 21312 5102
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21284 4078 21312 4762
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 21376 3398 21404 5102
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21468 2774 21496 6054
rect 21560 5370 21588 9046
rect 21652 8906 21680 9318
rect 21640 8900 21692 8906
rect 21640 8842 21692 8848
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21744 6390 21772 8774
rect 21732 6384 21784 6390
rect 21732 6326 21784 6332
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21638 5808 21694 5817
rect 21638 5743 21694 5752
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21560 4282 21588 4490
rect 21652 4282 21680 5743
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21548 3120 21600 3126
rect 21548 3062 21600 3068
rect 21560 2854 21588 3062
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21008 2746 21220 2774
rect 21376 2746 21496 2774
rect 20812 1284 20864 1290
rect 20812 1226 20864 1232
rect 21008 800 21036 2746
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21284 1970 21312 2246
rect 21272 1964 21324 1970
rect 21272 1906 21324 1912
rect 21376 800 21404 2746
rect 21744 800 21772 6190
rect 21836 4049 21864 9454
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21928 7546 21956 7890
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21928 6322 21956 7482
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 21916 5568 21968 5574
rect 21914 5536 21916 5545
rect 21968 5536 21970 5545
rect 21914 5471 21970 5480
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21928 4486 21956 5306
rect 22020 4622 22048 9574
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22112 7954 22140 9454
rect 22296 9194 22324 9658
rect 22296 9166 22416 9194
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 22112 4282 22140 4966
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 21916 4208 21968 4214
rect 21916 4150 21968 4156
rect 22020 4162 22048 4218
rect 21822 4040 21878 4049
rect 21822 3975 21878 3984
rect 21928 3890 21956 4150
rect 22020 4134 22140 4162
rect 21928 3862 22048 3890
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21928 3058 21956 3674
rect 22020 3058 22048 3862
rect 22112 3398 22140 4134
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22204 3126 22232 5170
rect 22296 3126 22324 8434
rect 22388 7818 22416 9166
rect 22480 8906 22508 11290
rect 22572 10742 22600 12650
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 22664 10674 22692 12718
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22572 9994 22600 10134
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22572 9897 22600 9930
rect 22558 9888 22614 9897
rect 22558 9823 22614 9832
rect 22664 9518 22692 10610
rect 22756 10606 22784 17190
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22848 15162 22876 17070
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 22940 16182 22968 16730
rect 23308 16674 23336 21830
rect 23386 19544 23442 19553
rect 23492 19514 23520 22918
rect 23584 21350 23612 23598
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23386 19479 23442 19488
rect 23480 19508 23532 19514
rect 23400 18834 23428 19479
rect 23480 19450 23532 19456
rect 23584 19446 23612 20334
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23676 19446 23704 19994
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23584 17626 23612 19382
rect 23492 17598 23612 17626
rect 23492 17202 23520 17598
rect 23768 17270 23796 28698
rect 23860 27538 23888 29242
rect 23952 28422 23980 29566
rect 24124 28960 24176 28966
rect 24124 28902 24176 28908
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 23952 28150 23980 28358
rect 23940 28144 23992 28150
rect 23940 28086 23992 28092
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23952 27470 23980 28086
rect 24030 27704 24086 27713
rect 24030 27639 24086 27648
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23952 27062 23980 27406
rect 23940 27056 23992 27062
rect 23940 26998 23992 27004
rect 23848 25220 23900 25226
rect 23848 25162 23900 25168
rect 23860 24449 23888 25162
rect 23952 24886 23980 26998
rect 24044 26382 24072 27639
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 23940 24880 23992 24886
rect 23940 24822 23992 24828
rect 23952 24614 23980 24822
rect 23940 24608 23992 24614
rect 23940 24550 23992 24556
rect 23846 24440 23902 24449
rect 23846 24375 23902 24384
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23860 22642 23888 23802
rect 23952 23798 23980 24550
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23952 23526 23980 23734
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 24044 21457 24072 21558
rect 24030 21448 24086 21457
rect 24030 21383 24086 21392
rect 24044 21350 24072 21383
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24044 20602 24072 21286
rect 24032 20596 24084 20602
rect 24032 20538 24084 20544
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 23952 18290 23980 20198
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24136 18086 24164 28902
rect 24228 28218 24256 33798
rect 24596 31754 24624 35430
rect 24860 35080 24912 35086
rect 24858 35048 24860 35057
rect 24912 35048 24914 35057
rect 24858 34983 24914 34992
rect 24768 33312 24820 33318
rect 24768 33254 24820 33260
rect 24780 32609 24808 33254
rect 24860 32768 24912 32774
rect 24860 32710 24912 32716
rect 24766 32600 24822 32609
rect 24872 32586 24900 32710
rect 24872 32558 24992 32586
rect 24766 32535 24822 32544
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24504 31726 24624 31754
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24216 28212 24268 28218
rect 24216 28154 24268 28160
rect 24216 20936 24268 20942
rect 24216 20878 24268 20884
rect 24228 20058 24256 20878
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24228 19446 24256 19654
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24412 18698 24440 28358
rect 24504 18698 24532 31726
rect 24872 29714 24900 31962
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 24596 29510 24624 29582
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24596 28529 24624 29446
rect 24872 29345 24900 29514
rect 24858 29336 24914 29345
rect 24858 29271 24914 29280
rect 24964 29186 24992 32558
rect 25056 32042 25084 38694
rect 25148 35834 25176 40718
rect 25136 35828 25188 35834
rect 25136 35770 25188 35776
rect 25240 35018 25268 45222
rect 25424 44849 25452 45426
rect 25410 44840 25466 44849
rect 25320 44804 25372 44810
rect 25410 44775 25466 44784
rect 25320 44746 25372 44752
rect 25332 44538 25360 44746
rect 25504 44736 25556 44742
rect 25504 44678 25556 44684
rect 25320 44532 25372 44538
rect 25320 44474 25372 44480
rect 25320 43716 25372 43722
rect 25320 43658 25372 43664
rect 25332 43450 25360 43658
rect 25320 43444 25372 43450
rect 25320 43386 25372 43392
rect 25320 41472 25372 41478
rect 25320 41414 25372 41420
rect 25332 41206 25360 41414
rect 25320 41200 25372 41206
rect 25320 41142 25372 41148
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25332 40526 25360 40695
rect 25320 40520 25372 40526
rect 25320 40462 25372 40468
rect 25412 40384 25464 40390
rect 25412 40326 25464 40332
rect 25320 40044 25372 40050
rect 25320 39986 25372 39992
rect 25332 39953 25360 39986
rect 25318 39944 25374 39953
rect 25318 39879 25374 39888
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 25332 39137 25360 39374
rect 25318 39128 25374 39137
rect 25318 39063 25374 39072
rect 25320 38276 25372 38282
rect 25320 38218 25372 38224
rect 25332 38010 25360 38218
rect 25320 38004 25372 38010
rect 25320 37946 25372 37952
rect 25320 37188 25372 37194
rect 25320 37130 25372 37136
rect 25332 36922 25360 37130
rect 25320 36916 25372 36922
rect 25320 36858 25372 36864
rect 25320 35692 25372 35698
rect 25320 35634 25372 35640
rect 25332 35290 25360 35634
rect 25320 35284 25372 35290
rect 25320 35226 25372 35232
rect 25228 35012 25280 35018
rect 25228 34954 25280 34960
rect 25228 34740 25280 34746
rect 25228 34682 25280 34688
rect 25240 33130 25268 34682
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25318 34167 25374 34176
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25332 33425 25360 33934
rect 25318 33416 25374 33425
rect 25318 33351 25374 33360
rect 25240 33102 25360 33130
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 25228 32972 25280 32978
rect 25228 32914 25280 32920
rect 25148 32570 25176 32914
rect 25136 32564 25188 32570
rect 25136 32506 25188 32512
rect 25240 32366 25268 32914
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25056 32014 25176 32042
rect 25044 31952 25096 31958
rect 25044 31894 25096 31900
rect 24872 29158 24992 29186
rect 24872 28626 24900 29158
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24964 28558 24992 29038
rect 24952 28552 25004 28558
rect 24582 28520 24638 28529
rect 24952 28494 25004 28500
rect 24582 28455 24638 28464
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24780 27130 24808 27542
rect 25056 27538 25084 31894
rect 25148 31482 25176 32014
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 25056 26586 25084 27270
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 24860 26512 24912 26518
rect 24860 26454 24912 26460
rect 24872 23202 24900 26454
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 24952 26036 25004 26042
rect 24952 25978 25004 25984
rect 24964 23746 24992 25978
rect 25056 24750 25084 26386
rect 25148 26314 25176 31078
rect 25240 30190 25268 32302
rect 25332 32026 25360 33102
rect 25424 32910 25452 40326
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25412 32564 25464 32570
rect 25412 32506 25464 32512
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25228 30184 25280 30190
rect 25228 30126 25280 30132
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 29306 25360 29582
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25424 28626 25452 32506
rect 25516 31482 25544 44678
rect 25596 37324 25648 37330
rect 25596 37266 25648 37272
rect 25504 31476 25556 31482
rect 25504 31418 25556 31424
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25516 30977 25544 31282
rect 25502 30968 25558 30977
rect 25502 30903 25504 30912
rect 25556 30903 25558 30912
rect 25504 30874 25556 30880
rect 25412 28620 25464 28626
rect 25412 28562 25464 28568
rect 25228 27872 25280 27878
rect 25228 27814 25280 27820
rect 25240 27334 25268 27814
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25410 26888 25466 26897
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25265 25176 25774
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25240 24750 25268 26862
rect 25410 26823 25466 26832
rect 25318 26072 25374 26081
rect 25318 26007 25374 26016
rect 25332 25294 25360 26007
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25056 23866 25084 24686
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 24964 23718 25084 23746
rect 24872 23174 24992 23202
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24872 22817 24900 22986
rect 24858 22808 24914 22817
rect 24858 22743 24914 22752
rect 24964 22658 24992 23174
rect 24872 22630 24992 22658
rect 24872 22098 24900 22630
rect 24860 22092 24912 22098
rect 25056 22094 25084 23718
rect 25134 23624 25190 23633
rect 25134 23559 25190 23568
rect 25148 22710 25176 23559
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 25240 22234 25268 24686
rect 25332 23866 25360 25230
rect 25424 24206 25452 26823
rect 25504 26376 25556 26382
rect 25504 26318 25556 26324
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25332 23050 25360 23462
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25228 22228 25280 22234
rect 25228 22170 25280 22176
rect 24860 22034 24912 22040
rect 24964 22066 25084 22094
rect 24858 21176 24914 21185
rect 24768 21140 24820 21146
rect 24858 21111 24914 21120
rect 24768 21082 24820 21088
rect 24674 20360 24730 20369
rect 24674 20295 24730 20304
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24596 18766 24624 19654
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24400 18692 24452 18698
rect 24400 18634 24452 18640
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 24688 18222 24716 20295
rect 24780 19854 24808 21082
rect 24872 21010 24900 21111
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24964 20874 24992 22066
rect 25424 21486 25452 23122
rect 25412 21480 25464 21486
rect 25412 21422 25464 21428
rect 25044 21072 25096 21078
rect 25044 21014 25096 21020
rect 24952 20868 25004 20874
rect 24952 20810 25004 20816
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24858 18728 24914 18737
rect 24858 18663 24914 18672
rect 24952 18692 25004 18698
rect 24872 18358 24900 18663
rect 24952 18634 25004 18640
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 24858 17912 24914 17921
rect 24858 17847 24914 17856
rect 24872 17746 24900 17847
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23216 16646 23336 16674
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 23216 16130 23244 16646
rect 23492 16266 23520 17138
rect 23846 17096 23902 17105
rect 23846 17031 23902 17040
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23308 16250 23520 16266
rect 23296 16244 23520 16250
rect 23348 16238 23520 16244
rect 23296 16186 23348 16192
rect 23216 16102 23336 16130
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23308 15586 23336 16102
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23216 15558 23336 15586
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 23216 15094 23244 15558
rect 23294 15464 23350 15473
rect 23294 15399 23350 15408
rect 23308 15094 23336 15399
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22848 12986 22876 13942
rect 23204 13864 23256 13870
rect 23256 13824 23336 13852
rect 23204 13806 23256 13812
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22848 12374 22876 12922
rect 23308 12918 23336 13824
rect 23400 13258 23428 14010
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22848 11354 22876 12174
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22834 11248 22890 11257
rect 23308 11234 23336 12242
rect 22834 11183 22890 11192
rect 23216 11206 23336 11234
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22558 9072 22614 9081
rect 22558 9007 22614 9016
rect 22572 8974 22600 9007
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22388 5545 22416 6802
rect 22374 5536 22430 5545
rect 22374 5471 22430 5480
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22020 2446 22048 2586
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22098 2408 22154 2417
rect 22098 2343 22154 2352
rect 22112 1834 22140 2343
rect 22100 1828 22152 1834
rect 22100 1770 22152 1776
rect 22204 1601 22232 2518
rect 22296 2446 22324 2926
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22190 1592 22246 1601
rect 22190 1527 22246 1536
rect 22112 870 22232 898
rect 22112 800 22140 870
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22204 762 22232 870
rect 22388 762 22416 3402
rect 22480 800 22508 8366
rect 22756 7313 22784 9998
rect 22848 9178 22876 11183
rect 23216 10810 23244 11206
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23308 9330 23336 11086
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23400 10577 23428 11018
rect 23386 10568 23442 10577
rect 23386 10503 23442 10512
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23400 10130 23428 10406
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23400 9518 23428 10066
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23308 9302 23428 9330
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22848 7970 22876 8502
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22848 7942 22968 7970
rect 22940 7546 22968 7942
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 22742 7304 22798 7313
rect 22742 7239 22798 7248
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22742 7032 22798 7041
rect 22950 7035 23258 7044
rect 22560 6996 22612 7002
rect 22742 6967 22798 6976
rect 22560 6938 22612 6944
rect 22204 734 22416 762
rect 22466 0 22522 800
rect 22572 762 22600 6938
rect 22652 6928 22704 6934
rect 22652 6870 22704 6876
rect 22664 3058 22692 6870
rect 22756 4282 22784 6967
rect 23308 6882 23336 9114
rect 23400 8090 23428 9302
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23216 6854 23336 6882
rect 23018 6352 23074 6361
rect 23018 6287 23074 6296
rect 23032 6254 23060 6287
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 23216 6202 23244 6854
rect 23400 6474 23428 7482
rect 23492 7410 23520 15914
rect 23584 15366 23612 16662
rect 23860 16590 23888 17031
rect 24228 16794 24256 17206
rect 24596 16794 24624 17614
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23584 13734 23612 15302
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23846 13832 23902 13841
rect 23846 13767 23902 13776
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23860 13326 23888 13767
rect 23952 13530 23980 14350
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 24136 12442 24164 14962
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 23860 10198 23888 10678
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 23952 9178 23980 11698
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23756 7744 23808 7750
rect 23676 7692 23756 7698
rect 23676 7686 23808 7692
rect 23676 7670 23796 7686
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23676 6934 23704 7670
rect 23664 6928 23716 6934
rect 23664 6870 23716 6876
rect 23400 6446 23612 6474
rect 23676 6458 23704 6870
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23768 6458 23796 6598
rect 23216 6174 23336 6202
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23110 5672 23166 5681
rect 23110 5607 23166 5616
rect 23124 5574 23152 5607
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 23308 4214 23336 6174
rect 23478 5808 23534 5817
rect 23478 5743 23534 5752
rect 23492 5642 23520 5743
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 23400 4865 23428 5578
rect 23584 5522 23612 6446
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23492 5494 23612 5522
rect 23386 4856 23442 4865
rect 23386 4791 23442 4800
rect 23492 4706 23520 5494
rect 23400 4678 23520 4706
rect 23662 4720 23718 4729
rect 23296 4208 23348 4214
rect 23296 4150 23348 4156
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23204 3664 23256 3670
rect 23204 3606 23256 3612
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 3126 22876 3334
rect 23216 3233 23244 3606
rect 23202 3224 23258 3233
rect 23202 3159 23258 3168
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 23400 2774 23428 4678
rect 23662 4655 23718 4664
rect 23676 4554 23704 4655
rect 23754 4584 23810 4593
rect 23664 4548 23716 4554
rect 23754 4519 23810 4528
rect 23664 4490 23716 4496
rect 23768 4486 23796 4519
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23492 3738 23520 4082
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23860 3194 23888 8298
rect 23940 8016 23992 8022
rect 23940 7958 23992 7964
rect 23952 7449 23980 7958
rect 23938 7440 23994 7449
rect 23938 7375 23940 7384
rect 23992 7375 23994 7384
rect 23940 7346 23992 7352
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 23952 5681 23980 6734
rect 23938 5672 23994 5681
rect 23938 5607 23994 5616
rect 24044 4146 24072 10950
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24136 9518 24164 10134
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24136 7886 24164 9454
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24136 7750 24164 7822
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 6390 24164 7686
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24136 5914 24164 6326
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 24044 4026 24072 4082
rect 24044 3998 24164 4026
rect 24032 3936 24084 3942
rect 24030 3904 24032 3913
rect 24084 3904 24086 3913
rect 24030 3839 24086 3848
rect 23938 3496 23994 3505
rect 23938 3431 23994 3440
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23570 2952 23626 2961
rect 23570 2887 23626 2896
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23308 2746 23428 2774
rect 23308 2564 23336 2746
rect 23216 2536 23336 2564
rect 22756 870 22876 898
rect 22756 762 22784 870
rect 22848 800 22876 870
rect 23216 800 23244 2536
rect 23584 800 23612 2887
rect 23952 800 23980 3431
rect 24136 3194 24164 3998
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24228 3058 24256 11630
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24320 6390 24348 10202
rect 24412 9586 24440 15642
rect 24596 10266 24624 15982
rect 24688 15570 24716 17478
rect 24766 16280 24822 16289
rect 24766 16215 24822 16224
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24780 14958 24808 16215
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24688 10062 24716 14826
rect 24858 14648 24914 14657
rect 24858 14583 24914 14592
rect 24872 14482 24900 14583
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 10849 24808 12174
rect 24872 11914 24900 14214
rect 24964 12434 24992 18634
rect 25056 17746 25084 21014
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 19514 25176 20334
rect 25332 20058 25360 20810
rect 25424 20602 25452 21422
rect 25516 20942 25544 26318
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25148 17746 25176 19450
rect 25228 18148 25280 18154
rect 25228 18090 25280 18096
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 25056 14414 25084 17546
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25240 13938 25268 18090
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 13394 25084 13670
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 25134 13016 25190 13025
rect 25134 12951 25190 12960
rect 24964 12406 25084 12434
rect 24950 12200 25006 12209
rect 24950 12135 24952 12144
rect 25004 12135 25006 12144
rect 24952 12106 25004 12112
rect 24872 11886 24992 11914
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24872 11393 24900 11766
rect 24964 11762 24992 11886
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24766 10840 24822 10849
rect 24766 10775 24822 10784
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24398 7848 24454 7857
rect 24398 7783 24454 7792
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24320 5914 24348 6326
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 24412 4826 24440 7783
rect 24492 6656 24544 6662
rect 24492 6598 24544 6604
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24308 4548 24360 4554
rect 24308 4490 24360 4496
rect 24320 4146 24348 4490
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 24320 800 24348 4082
rect 24504 2106 24532 6598
rect 24596 5710 24624 8366
rect 24688 6662 24716 9862
rect 24766 9752 24822 9761
rect 24766 9687 24822 9696
rect 24780 8430 24808 9687
rect 24950 8936 25006 8945
rect 24950 8871 24952 8880
rect 25004 8871 25006 8880
rect 24952 8842 25004 8848
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24950 7984 25006 7993
rect 24950 7919 25006 7928
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24872 7313 24900 7414
rect 24858 7304 24914 7313
rect 24768 7268 24820 7274
rect 24858 7239 24914 7248
rect 24768 7210 24820 7216
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 24596 3534 24624 3878
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 2446 24624 3334
rect 24688 3194 24716 6258
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24780 2774 24808 7210
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 24872 6497 24900 6666
rect 24858 6488 24914 6497
rect 24858 6423 24914 6432
rect 24964 5846 24992 7919
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 25056 5234 25084 12406
rect 25148 11830 25176 12951
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25608 11286 25636 37266
rect 25700 29866 25728 47466
rect 25792 30054 25820 51274
rect 25872 38208 25924 38214
rect 25872 38150 25924 38156
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 25700 29838 25820 29866
rect 25688 29776 25740 29782
rect 25688 29718 25740 29724
rect 25700 23118 25728 29718
rect 25792 23322 25820 29838
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25884 22094 25912 38150
rect 25976 32230 26004 52430
rect 26148 48612 26200 48618
rect 26148 48554 26200 48560
rect 26056 35488 26108 35494
rect 26056 35430 26108 35436
rect 25964 32224 26016 32230
rect 25964 32166 26016 32172
rect 25964 27872 26016 27878
rect 25964 27814 26016 27820
rect 25976 26314 26004 27814
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 25976 23526 26004 26250
rect 25964 23520 26016 23526
rect 25964 23462 26016 23468
rect 25792 22066 25912 22094
rect 25792 11558 25820 22066
rect 26068 17882 26096 35430
rect 26160 31754 26188 48554
rect 26516 47184 26568 47190
rect 26516 47126 26568 47132
rect 26160 31726 26280 31754
rect 26148 31476 26200 31482
rect 26148 31418 26200 31424
rect 26160 18426 26188 31418
rect 26252 25974 26280 31726
rect 26528 29170 26556 47126
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26240 25968 26292 25974
rect 26240 25910 26292 25916
rect 26148 18420 26200 18426
rect 26148 18362 26200 18368
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 25596 11280 25648 11286
rect 25596 11222 25648 11228
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 24780 2746 24900 2774
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24492 2100 24544 2106
rect 24492 2042 24544 2048
rect 22572 734 22784 762
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24872 785 24900 2746
rect 24858 776 24914 785
rect 24858 711 24914 720
rect 25042 0 25098 800
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3422 8744 3478 8800
rect 4066 6432 4122 6488
rect 3790 4120 3846 4176
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3974 1844 3976 1864
rect 3976 1844 4028 1864
rect 4028 1844 4030 1864
rect 3974 1808 4030 1844
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 23386 56072 23442 56128
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 8850 12280 8906 12336
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 10046 9016 10102 9072
rect 9954 7384 10010 7440
rect 11518 10512 11574 10568
rect 10874 6196 10876 6216
rect 10876 6196 10928 6216
rect 10928 6196 10930 6216
rect 10874 6160 10930 6196
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 13450 25764 13506 25800
rect 13450 25744 13452 25764
rect 13452 25744 13504 25764
rect 13504 25744 13506 25764
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 13542 25336 13598 25392
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 15566 27276 15568 27296
rect 15568 27276 15620 27296
rect 15620 27276 15622 27296
rect 15566 27240 15622 27276
rect 15290 24792 15346 24848
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 11978 11056 12034 11112
rect 11426 9424 11482 9480
rect 12346 11620 12402 11656
rect 12346 11600 12348 11620
rect 12348 11600 12400 11620
rect 12400 11600 12402 11620
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13358 11736 13414 11792
rect 12254 4528 12310 4584
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13542 12280 13598 12336
rect 13542 11892 13598 11928
rect 13542 11872 13544 11892
rect 13544 11872 13596 11892
rect 13596 11872 13598 11892
rect 13542 11228 13544 11248
rect 13544 11228 13596 11248
rect 13596 11228 13598 11248
rect 13542 11192 13598 11228
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12714 6432 12770 6488
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 13450 6704 13506 6760
rect 13450 6296 13506 6352
rect 12990 6196 12992 6216
rect 12992 6196 13044 6216
rect 13044 6196 13046 6216
rect 12990 6160 13046 6196
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 14738 12416 14794 12472
rect 13818 8336 13874 8392
rect 13082 5228 13138 5264
rect 13082 5208 13084 5228
rect 13084 5208 13136 5228
rect 13136 5208 13138 5228
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14554 10512 14610 10568
rect 16302 25200 16358 25256
rect 15106 11600 15162 11656
rect 14370 6860 14426 6896
rect 14370 6840 14372 6860
rect 14372 6840 14424 6860
rect 14424 6840 14426 6860
rect 14186 5908 14242 5944
rect 14186 5888 14188 5908
rect 14188 5888 14240 5908
rect 14240 5888 14242 5908
rect 14738 5244 14740 5264
rect 14740 5244 14792 5264
rect 14792 5244 14794 5264
rect 14738 5208 14794 5244
rect 15290 10240 15346 10296
rect 15198 7248 15254 7304
rect 15382 6316 15438 6352
rect 15382 6296 15384 6316
rect 15384 6296 15436 6316
rect 15436 6296 15438 6316
rect 15198 6160 15254 6216
rect 15474 5752 15530 5808
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 16026 12144 16082 12200
rect 16026 11872 16082 11928
rect 16026 11192 16082 11248
rect 16854 18264 16910 18320
rect 17130 25744 17186 25800
rect 17406 25644 17408 25664
rect 17408 25644 17460 25664
rect 17460 25644 17462 25664
rect 17406 25608 17462 25644
rect 17222 22752 17278 22808
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17590 25336 17646 25392
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 16118 9988 16174 10024
rect 16118 9968 16120 9988
rect 16120 9968 16172 9988
rect 16172 9968 16174 9988
rect 15934 8472 15990 8528
rect 17130 17856 17186 17912
rect 17222 16108 17278 16144
rect 17222 16088 17224 16108
rect 17224 16088 17276 16108
rect 17276 16088 17278 16108
rect 17130 15272 17186 15328
rect 17314 13524 17370 13560
rect 17314 13504 17316 13524
rect 17316 13504 17368 13524
rect 17368 13504 17370 13524
rect 16854 10648 16910 10704
rect 16946 10376 17002 10432
rect 16394 4664 16450 4720
rect 18510 27820 18512 27840
rect 18512 27820 18564 27840
rect 18564 27820 18566 27840
rect 18510 27784 18566 27820
rect 18418 25236 18420 25256
rect 18420 25236 18472 25256
rect 18472 25236 18474 25256
rect 18418 25200 18474 25236
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17866 17856 17922 17912
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17222 11056 17278 11112
rect 17406 6432 17462 6488
rect 17774 11736 17830 11792
rect 18878 23432 18934 23488
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18510 13776 18566 13832
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18418 12416 18474 12472
rect 18510 12280 18566 12336
rect 18326 10124 18382 10160
rect 18326 10104 18328 10124
rect 18328 10104 18380 10124
rect 18380 10104 18382 10124
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18234 8336 18290 8392
rect 17682 7928 17738 7984
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17774 5752 17830 5808
rect 18510 10240 18566 10296
rect 18786 12280 18842 12336
rect 18694 12164 18750 12200
rect 18694 12144 18696 12164
rect 18696 12144 18748 12164
rect 18748 12144 18750 12164
rect 18878 10376 18934 10432
rect 18694 10104 18750 10160
rect 18694 9696 18750 9752
rect 18602 7112 18658 7168
rect 18510 5752 18566 5808
rect 18418 5616 18474 5672
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17774 2896 17830 2952
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 19890 23568 19946 23624
rect 19522 15136 19578 15192
rect 19246 11056 19302 11112
rect 19062 10648 19118 10704
rect 19522 10920 19578 10976
rect 19522 10784 19578 10840
rect 19430 10104 19486 10160
rect 18878 9288 18934 9344
rect 19246 9424 19302 9480
rect 19246 9324 19248 9344
rect 19248 9324 19300 9344
rect 19300 9324 19302 9344
rect 19246 9288 19302 9324
rect 18970 7112 19026 7168
rect 18970 6976 19026 7032
rect 19522 8200 19578 8256
rect 19430 4664 19486 4720
rect 19614 4664 19670 4720
rect 20258 14456 20314 14512
rect 20166 9968 20222 10024
rect 21086 13776 21142 13832
rect 20442 7828 20444 7848
rect 20444 7828 20496 7848
rect 20496 7828 20498 7848
rect 20442 7792 20498 7828
rect 20718 10104 20774 10160
rect 20718 7284 20720 7304
rect 20720 7284 20772 7304
rect 20772 7284 20774 7304
rect 20718 7248 20774 7284
rect 20626 6704 20682 6760
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 21362 12688 21418 12744
rect 21362 11892 21418 11928
rect 21362 11872 21364 11892
rect 21364 11872 21416 11892
rect 21416 11872 21418 11892
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 25318 55392 25374 55448
rect 24766 54576 24822 54632
rect 24858 53760 24914 53816
rect 25502 52964 25558 53000
rect 25502 52944 25504 52964
rect 25504 52944 25556 52964
rect 25556 52944 25558 52964
rect 24950 52148 25006 52184
rect 24950 52128 24952 52148
rect 24952 52128 25004 52148
rect 25004 52128 25006 52148
rect 24950 51332 25006 51368
rect 24950 51312 24952 51332
rect 24952 51312 25004 51332
rect 25004 51312 25006 51332
rect 24766 49680 24822 49736
rect 24858 48884 24914 48920
rect 24858 48864 24860 48884
rect 24860 48864 24912 48884
rect 24912 48864 24914 48884
rect 24858 48084 24860 48104
rect 24860 48084 24912 48104
rect 24912 48084 24914 48104
rect 24858 48048 24914 48084
rect 25042 50496 25098 50552
rect 25318 47232 25374 47288
rect 25318 46416 25374 46472
rect 24674 43968 24730 44024
rect 24950 43152 25006 43208
rect 24858 42356 24914 42392
rect 24858 42336 24860 42356
rect 24860 42336 24912 42356
rect 24912 42336 24914 42356
rect 24858 41556 24860 41576
rect 24860 41556 24912 41576
rect 24912 41556 24914 41576
rect 24858 41520 24914 41556
rect 25318 45600 25374 45656
rect 24858 38800 24914 38856
rect 24766 38256 24822 38312
rect 24858 37440 24914 37496
rect 24950 36624 25006 36680
rect 24766 35808 24822 35864
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22466 21412 22522 21448
rect 22466 21392 22468 21412
rect 22468 21392 22520 21412
rect 22520 21392 22522 21412
rect 22282 17856 22338 17912
rect 21178 10920 21234 10976
rect 21638 9832 21694 9888
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23294 21936 23350 21992
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22466 11464 22522 11520
rect 22282 9968 22338 10024
rect 21638 5752 21694 5808
rect 21914 5516 21916 5536
rect 21916 5516 21968 5536
rect 21968 5516 21970 5536
rect 21914 5480 21970 5516
rect 21822 3984 21878 4040
rect 22558 9832 22614 9888
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23386 19488 23442 19544
rect 24030 27648 24086 27704
rect 23846 24384 23902 24440
rect 24030 21392 24086 21448
rect 24858 35028 24860 35048
rect 24860 35028 24912 35048
rect 24912 35028 24914 35048
rect 24858 34992 24914 35028
rect 24766 32544 24822 32600
rect 24858 29280 24914 29336
rect 25410 44784 25466 44840
rect 25318 40704 25374 40760
rect 25318 39888 25374 39944
rect 25318 39072 25374 39128
rect 25318 34176 25374 34232
rect 25318 33360 25374 33416
rect 24582 28464 24638 28520
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30096 25374 30152
rect 25502 30932 25558 30968
rect 25502 30912 25504 30932
rect 25504 30912 25556 30932
rect 25556 30912 25558 30932
rect 25134 25200 25190 25256
rect 25410 26832 25466 26888
rect 25318 26016 25374 26072
rect 24858 22752 24914 22808
rect 25134 23568 25190 23624
rect 24858 21120 24914 21176
rect 24674 20304 24730 20360
rect 24858 18672 24914 18728
rect 24858 17856 24914 17912
rect 23846 17040 23902 17096
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 23294 15408 23350 15464
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22834 11192 22890 11248
rect 22558 9016 22614 9072
rect 22374 5480 22430 5536
rect 22098 2352 22154 2408
rect 22190 1536 22246 1592
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23386 10512 23442 10568
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22742 7248 22798 7304
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22742 6976 22798 7032
rect 23018 6296 23074 6352
rect 23846 13776 23902 13832
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 23110 5616 23166 5672
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 23478 5752 23534 5808
rect 23386 4800 23442 4856
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23202 3168 23258 3224
rect 23662 4664 23718 4720
rect 23754 4528 23810 4584
rect 23938 7404 23994 7440
rect 23938 7384 23940 7404
rect 23940 7384 23992 7404
rect 23992 7384 23994 7404
rect 23938 5616 23994 5672
rect 24030 3884 24032 3904
rect 24032 3884 24084 3904
rect 24084 3884 24086 3904
rect 24030 3848 24086 3884
rect 23938 3440 23994 3496
rect 23570 2896 23626 2952
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24766 16224 24822 16280
rect 24858 14592 24914 14648
rect 25134 12960 25190 13016
rect 24950 12164 25006 12200
rect 24950 12144 24952 12164
rect 24952 12144 25004 12164
rect 25004 12144 25006 12164
rect 24858 11328 24914 11384
rect 24766 10784 24822 10840
rect 24398 7792 24454 7848
rect 24766 9696 24822 9752
rect 24950 8900 25006 8936
rect 24950 8880 24952 8900
rect 24952 8880 25004 8900
rect 25004 8880 25006 8900
rect 24950 7928 25006 7984
rect 24858 7248 24914 7304
rect 24858 6432 24914 6488
rect 25134 8064 25190 8120
rect 24858 720 24914 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23430 56133 23490 56206
rect 26200 56176 27000 56206
rect 23381 56128 23490 56133
rect 23381 56072 23386 56128
rect 23442 56072 23490 56128
rect 23381 56070 23490 56072
rect 23381 56067 23447 56070
rect 25313 55450 25379 55453
rect 26200 55450 27000 55480
rect 25313 55448 27000 55450
rect 25313 55392 25318 55448
rect 25374 55392 27000 55448
rect 25313 55390 27000 55392
rect 25313 55387 25379 55390
rect 26200 55360 27000 55390
rect 24761 54634 24827 54637
rect 26200 54634 27000 54664
rect 24761 54632 27000 54634
rect 24761 54576 24766 54632
rect 24822 54576 27000 54632
rect 24761 54574 27000 54576
rect 24761 54571 24827 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 24853 53818 24919 53821
rect 26200 53818 27000 53848
rect 24853 53816 27000 53818
rect 24853 53760 24858 53816
rect 24914 53760 27000 53816
rect 24853 53758 27000 53760
rect 24853 53755 24919 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 25497 53002 25563 53005
rect 26200 53002 27000 53032
rect 25497 53000 27000 53002
rect 25497 52944 25502 53000
rect 25558 52944 27000 53000
rect 25497 52942 27000 52944
rect 25497 52939 25563 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24945 52186 25011 52189
rect 26200 52186 27000 52216
rect 24945 52184 27000 52186
rect 24945 52128 24950 52184
rect 25006 52128 27000 52184
rect 24945 52126 27000 52128
rect 24945 52123 25011 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 24945 51370 25011 51373
rect 26200 51370 27000 51400
rect 24945 51368 27000 51370
rect 24945 51312 24950 51368
rect 25006 51312 27000 51368
rect 24945 51310 27000 51312
rect 24945 51307 25011 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 25037 50554 25103 50557
rect 26200 50554 27000 50584
rect 25037 50552 27000 50554
rect 25037 50496 25042 50552
rect 25098 50496 27000 50552
rect 25037 50494 27000 50496
rect 25037 50491 25103 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 24761 49738 24827 49741
rect 26200 49738 27000 49768
rect 24761 49736 27000 49738
rect 24761 49680 24766 49736
rect 24822 49680 27000 49736
rect 24761 49678 27000 49680
rect 24761 49675 24827 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 24853 48922 24919 48925
rect 26200 48922 27000 48952
rect 24853 48920 27000 48922
rect 24853 48864 24858 48920
rect 24914 48864 27000 48920
rect 24853 48862 27000 48864
rect 24853 48859 24919 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 24853 48106 24919 48109
rect 26200 48106 27000 48136
rect 24853 48104 27000 48106
rect 24853 48048 24858 48104
rect 24914 48048 27000 48104
rect 24853 48046 27000 48048
rect 24853 48043 24919 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25313 46474 25379 46477
rect 26200 46474 27000 46504
rect 25313 46472 27000 46474
rect 25313 46416 25318 46472
rect 25374 46416 27000 46472
rect 25313 46414 27000 46416
rect 25313 46411 25379 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 25313 45658 25379 45661
rect 26200 45658 27000 45688
rect 25313 45656 27000 45658
rect 25313 45600 25318 45656
rect 25374 45600 27000 45656
rect 25313 45598 27000 45600
rect 25313 45595 25379 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25405 44842 25471 44845
rect 26200 44842 27000 44872
rect 25405 44840 27000 44842
rect 25405 44784 25410 44840
rect 25466 44784 27000 44840
rect 25405 44782 27000 44784
rect 25405 44779 25471 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24669 44026 24735 44029
rect 26200 44026 27000 44056
rect 24669 44024 27000 44026
rect 24669 43968 24674 44024
rect 24730 43968 27000 44024
rect 24669 43966 27000 43968
rect 24669 43963 24735 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 24945 43210 25011 43213
rect 26200 43210 27000 43240
rect 24945 43208 27000 43210
rect 24945 43152 24950 43208
rect 25006 43152 27000 43208
rect 24945 43150 27000 43152
rect 24945 43147 25011 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 24853 42394 24919 42397
rect 26200 42394 27000 42424
rect 24853 42392 27000 42394
rect 24853 42336 24858 42392
rect 24914 42336 27000 42392
rect 24853 42334 27000 42336
rect 24853 42331 24919 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 24853 41578 24919 41581
rect 26200 41578 27000 41608
rect 24853 41576 27000 41578
rect 24853 41520 24858 41576
rect 24914 41520 27000 41576
rect 24853 41518 27000 41520
rect 24853 41515 24919 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 25313 39946 25379 39949
rect 26200 39946 27000 39976
rect 25313 39944 27000 39946
rect 25313 39888 25318 39944
rect 25374 39888 27000 39944
rect 25313 39886 27000 39888
rect 25313 39883 25379 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25313 39130 25379 39133
rect 26200 39130 27000 39160
rect 25313 39128 27000 39130
rect 25313 39072 25318 39128
rect 25374 39072 27000 39128
rect 25313 39070 27000 39072
rect 25313 39067 25379 39070
rect 26200 39040 27000 39070
rect 21398 38796 21404 38860
rect 21468 38858 21474 38860
rect 24853 38858 24919 38861
rect 21468 38856 24919 38858
rect 21468 38800 24858 38856
rect 24914 38800 24919 38856
rect 21468 38798 24919 38800
rect 21468 38796 21474 38798
rect 24853 38795 24919 38798
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 24761 38314 24827 38317
rect 26200 38314 27000 38344
rect 24761 38312 27000 38314
rect 24761 38256 24766 38312
rect 24822 38256 27000 38312
rect 24761 38254 27000 38256
rect 24761 38251 24827 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 24853 37498 24919 37501
rect 26200 37498 27000 37528
rect 24853 37496 27000 37498
rect 24853 37440 24858 37496
rect 24914 37440 27000 37496
rect 24853 37438 27000 37440
rect 24853 37435 24919 37438
rect 26200 37408 27000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 24945 36682 25011 36685
rect 26200 36682 27000 36712
rect 24945 36680 27000 36682
rect 24945 36624 24950 36680
rect 25006 36624 27000 36680
rect 24945 36622 27000 36624
rect 24945 36619 25011 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 24761 35866 24827 35869
rect 26200 35866 27000 35896
rect 24761 35864 27000 35866
rect 24761 35808 24766 35864
rect 24822 35808 27000 35864
rect 24761 35806 27000 35808
rect 24761 35803 24827 35806
rect 26200 35776 27000 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 24853 35050 24919 35053
rect 26200 35050 27000 35080
rect 24853 35048 27000 35050
rect 24853 34992 24858 35048
rect 24914 34992 27000 35048
rect 24853 34990 27000 34992
rect 24853 34987 24919 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 25313 33418 25379 33421
rect 26200 33418 27000 33448
rect 25313 33416 27000 33418
rect 25313 33360 25318 33416
rect 25374 33360 27000 33416
rect 25313 33358 27000 33360
rect 25313 33355 25379 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 24761 32602 24827 32605
rect 26200 32602 27000 32632
rect 24761 32600 27000 32602
rect 24761 32544 24766 32600
rect 24822 32544 27000 32600
rect 24761 32542 27000 32544
rect 24761 32539 24827 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 25497 30970 25563 30973
rect 26200 30970 27000 31000
rect 25497 30968 27000 30970
rect 25497 30912 25502 30968
rect 25558 30912 27000 30968
rect 25497 30910 27000 30912
rect 25497 30907 25563 30910
rect 26200 30880 27000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 24853 29338 24919 29341
rect 26200 29338 27000 29368
rect 24853 29336 27000 29338
rect 24853 29280 24858 29336
rect 24914 29280 27000 29336
rect 24853 29278 27000 29280
rect 24853 29275 24919 29278
rect 26200 29248 27000 29278
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 24577 28522 24643 28525
rect 26200 28522 27000 28552
rect 24577 28520 27000 28522
rect 24577 28464 24582 28520
rect 24638 28464 27000 28520
rect 24577 28462 27000 28464
rect 24577 28459 24643 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 18505 27844 18571 27845
rect 18454 27780 18460 27844
rect 18524 27842 18571 27844
rect 18524 27840 18616 27842
rect 18566 27784 18616 27840
rect 18524 27782 18616 27784
rect 18524 27780 18571 27782
rect 18505 27779 18571 27780
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24025 27706 24091 27709
rect 26200 27706 27000 27736
rect 24025 27704 27000 27706
rect 24025 27648 24030 27704
rect 24086 27648 27000 27704
rect 24025 27646 27000 27648
rect 24025 27643 24091 27646
rect 26200 27616 27000 27646
rect 15561 27298 15627 27301
rect 15694 27298 15700 27300
rect 15561 27296 15700 27298
rect 15561 27240 15566 27296
rect 15622 27240 15700 27296
rect 15561 27238 15700 27240
rect 15561 27235 15627 27238
rect 15694 27236 15700 27238
rect 15764 27236 15770 27300
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25405 26890 25471 26893
rect 26200 26890 27000 26920
rect 25405 26888 27000 26890
rect 25405 26832 25410 26888
rect 25466 26832 27000 26888
rect 25405 26830 27000 26832
rect 25405 26827 25471 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 25313 26074 25379 26077
rect 26200 26074 27000 26104
rect 25313 26072 27000 26074
rect 25313 26016 25318 26072
rect 25374 26016 27000 26072
rect 25313 26014 27000 26016
rect 25313 26011 25379 26014
rect 26200 25984 27000 26014
rect 13445 25802 13511 25805
rect 17125 25802 17191 25805
rect 13445 25800 17191 25802
rect 13445 25744 13450 25800
rect 13506 25744 17130 25800
rect 17186 25744 17191 25800
rect 13445 25742 17191 25744
rect 13445 25739 13511 25742
rect 17125 25739 17191 25742
rect 17401 25666 17467 25669
rect 17718 25666 17724 25668
rect 17401 25664 17724 25666
rect 17401 25608 17406 25664
rect 17462 25608 17724 25664
rect 17401 25606 17724 25608
rect 17401 25603 17467 25606
rect 17718 25604 17724 25606
rect 17788 25604 17794 25668
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 13537 25394 13603 25397
rect 17585 25394 17651 25397
rect 13537 25392 17651 25394
rect 13537 25336 13542 25392
rect 13598 25336 17590 25392
rect 17646 25336 17651 25392
rect 13537 25334 17651 25336
rect 13537 25331 13603 25334
rect 17585 25331 17651 25334
rect 16297 25258 16363 25261
rect 18413 25258 18479 25261
rect 16297 25256 18479 25258
rect 16297 25200 16302 25256
rect 16358 25200 18418 25256
rect 18474 25200 18479 25256
rect 16297 25198 18479 25200
rect 16297 25195 16363 25198
rect 18413 25195 18479 25198
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 15285 24850 15351 24853
rect 16430 24850 16436 24852
rect 15285 24848 16436 24850
rect 15285 24792 15290 24848
rect 15346 24792 16436 24848
rect 15285 24790 16436 24792
rect 15285 24787 15351 24790
rect 16430 24788 16436 24790
rect 16500 24788 16506 24852
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 23841 24442 23907 24445
rect 26200 24442 27000 24472
rect 23841 24440 27000 24442
rect 23841 24384 23846 24440
rect 23902 24384 27000 24440
rect 23841 24382 27000 24384
rect 23841 24379 23907 24382
rect 26200 24352 27000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 14222 23564 14228 23628
rect 14292 23626 14298 23628
rect 19885 23626 19951 23629
rect 14292 23624 19951 23626
rect 14292 23568 19890 23624
rect 19946 23568 19951 23624
rect 14292 23566 19951 23568
rect 14292 23564 14298 23566
rect 19885 23563 19951 23566
rect 25129 23626 25195 23629
rect 26200 23626 27000 23656
rect 25129 23624 27000 23626
rect 25129 23568 25134 23624
rect 25190 23568 27000 23624
rect 25129 23566 27000 23568
rect 25129 23563 25195 23566
rect 26200 23536 27000 23566
rect 18873 23490 18939 23493
rect 19006 23490 19012 23492
rect 18873 23488 19012 23490
rect 18873 23432 18878 23488
rect 18934 23432 19012 23488
rect 18873 23430 19012 23432
rect 18873 23427 18939 23430
rect 19006 23428 19012 23430
rect 19076 23428 19082 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 17217 22812 17283 22813
rect 17166 22810 17172 22812
rect 17126 22750 17172 22810
rect 17236 22808 17283 22812
rect 17278 22752 17283 22808
rect 17166 22748 17172 22750
rect 17236 22748 17283 22752
rect 17217 22747 17283 22748
rect 24853 22810 24919 22813
rect 26200 22810 27000 22840
rect 24853 22808 27000 22810
rect 24853 22752 24858 22808
rect 24914 22752 27000 22808
rect 24853 22750 27000 22752
rect 24853 22747 24919 22750
rect 26200 22720 27000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 23289 21994 23355 21997
rect 26200 21994 27000 22024
rect 23289 21992 27000 21994
rect 23289 21936 23294 21992
rect 23350 21936 27000 21992
rect 23289 21934 27000 21936
rect 23289 21931 23355 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 22461 21450 22527 21453
rect 24025 21450 24091 21453
rect 22461 21448 24091 21450
rect 22461 21392 22466 21448
rect 22522 21392 24030 21448
rect 24086 21392 24091 21448
rect 22461 21390 24091 21392
rect 22461 21387 22527 21390
rect 24025 21387 24091 21390
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 24853 21178 24919 21181
rect 26200 21178 27000 21208
rect 24853 21176 27000 21178
rect 24853 21120 24858 21176
rect 24914 21120 27000 21176
rect 24853 21118 27000 21120
rect 24853 21115 24919 21118
rect 26200 21088 27000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 24669 20362 24735 20365
rect 26200 20362 27000 20392
rect 24669 20360 27000 20362
rect 24669 20304 24674 20360
rect 24730 20304 27000 20360
rect 24669 20302 27000 20304
rect 24669 20299 24735 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 23381 19546 23447 19549
rect 26200 19546 27000 19576
rect 23381 19544 27000 19546
rect 23381 19488 23386 19544
rect 23442 19488 27000 19544
rect 23381 19486 27000 19488
rect 23381 19483 23447 19486
rect 26200 19456 27000 19486
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 24853 18730 24919 18733
rect 26200 18730 27000 18760
rect 24853 18728 27000 18730
rect 24853 18672 24858 18728
rect 24914 18672 27000 18728
rect 24853 18670 27000 18672
rect 24853 18667 24919 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 16849 18324 16915 18325
rect 16798 18322 16804 18324
rect 16758 18262 16804 18322
rect 16868 18320 16915 18324
rect 16910 18264 16915 18320
rect 16798 18260 16804 18262
rect 16868 18260 16915 18264
rect 16849 18259 16915 18260
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 17125 17914 17191 17917
rect 17718 17914 17724 17916
rect 17125 17912 17724 17914
rect 17125 17856 17130 17912
rect 17186 17856 17724 17912
rect 17125 17854 17724 17856
rect 17125 17851 17191 17854
rect 17718 17852 17724 17854
rect 17788 17914 17794 17916
rect 17861 17914 17927 17917
rect 17788 17912 17927 17914
rect 17788 17856 17866 17912
rect 17922 17856 17927 17912
rect 17788 17854 17927 17856
rect 17788 17852 17794 17854
rect 17861 17851 17927 17854
rect 20662 17852 20668 17916
rect 20732 17914 20738 17916
rect 22277 17914 22343 17917
rect 20732 17912 22343 17914
rect 20732 17856 22282 17912
rect 22338 17856 22343 17912
rect 20732 17854 22343 17856
rect 20732 17852 20738 17854
rect 22277 17851 22343 17854
rect 24853 17914 24919 17917
rect 26200 17914 27000 17944
rect 24853 17912 27000 17914
rect 24853 17856 24858 17912
rect 24914 17856 27000 17912
rect 24853 17854 27000 17856
rect 24853 17851 24919 17854
rect 26200 17824 27000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 23841 17098 23907 17101
rect 26200 17098 27000 17128
rect 23841 17096 27000 17098
rect 23841 17040 23846 17096
rect 23902 17040 27000 17096
rect 23841 17038 27000 17040
rect 23841 17035 23907 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 24761 16282 24827 16285
rect 26200 16282 27000 16312
rect 24761 16280 27000 16282
rect 24761 16224 24766 16280
rect 24822 16224 27000 16280
rect 24761 16222 27000 16224
rect 24761 16219 24827 16222
rect 26200 16192 27000 16222
rect 17217 16148 17283 16149
rect 17166 16084 17172 16148
rect 17236 16146 17283 16148
rect 17236 16144 17328 16146
rect 17278 16088 17328 16144
rect 17236 16086 17328 16088
rect 17236 16084 17283 16086
rect 17217 16083 17283 16084
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 23289 15466 23355 15469
rect 26200 15466 27000 15496
rect 23289 15464 27000 15466
rect 23289 15408 23294 15464
rect 23350 15408 27000 15464
rect 23289 15406 27000 15408
rect 23289 15403 23355 15406
rect 26200 15376 27000 15406
rect 16982 15268 16988 15332
rect 17052 15330 17058 15332
rect 17125 15330 17191 15333
rect 17052 15328 17191 15330
rect 17052 15272 17130 15328
rect 17186 15272 17191 15328
rect 17052 15270 17191 15272
rect 17052 15268 17058 15270
rect 17125 15267 17191 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 19517 15194 19583 15197
rect 20662 15194 20668 15196
rect 19517 15192 20668 15194
rect 19517 15136 19522 15192
rect 19578 15136 20668 15192
rect 19517 15134 20668 15136
rect 19517 15131 19583 15134
rect 20662 15132 20668 15134
rect 20732 15132 20738 15196
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 24853 14650 24919 14653
rect 26200 14650 27000 14680
rect 24853 14648 27000 14650
rect 24853 14592 24858 14648
rect 24914 14592 27000 14648
rect 24853 14590 27000 14592
rect 24853 14587 24919 14590
rect 26200 14560 27000 14590
rect 20253 14514 20319 14517
rect 21398 14514 21404 14516
rect 20253 14512 21404 14514
rect 20253 14456 20258 14512
rect 20314 14456 21404 14512
rect 20253 14454 21404 14456
rect 20253 14451 20319 14454
rect 21398 14452 21404 14454
rect 21468 14452 21474 14516
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 18505 13834 18571 13837
rect 18638 13834 18644 13836
rect 18505 13832 18644 13834
rect 18505 13776 18510 13832
rect 18566 13776 18644 13832
rect 18505 13774 18644 13776
rect 18505 13771 18571 13774
rect 18638 13772 18644 13774
rect 18708 13772 18714 13836
rect 20662 13772 20668 13836
rect 20732 13834 20738 13836
rect 21081 13834 21147 13837
rect 20732 13832 21147 13834
rect 20732 13776 21086 13832
rect 21142 13776 21147 13832
rect 20732 13774 21147 13776
rect 20732 13772 20738 13774
rect 21081 13771 21147 13774
rect 23841 13834 23907 13837
rect 26200 13834 27000 13864
rect 23841 13832 27000 13834
rect 23841 13776 23846 13832
rect 23902 13776 27000 13832
rect 23841 13774 27000 13776
rect 23841 13771 23907 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 16798 13500 16804 13564
rect 16868 13562 16874 13564
rect 17309 13562 17375 13565
rect 16868 13560 17375 13562
rect 16868 13504 17314 13560
rect 17370 13504 17375 13560
rect 16868 13502 17375 13504
rect 16868 13500 16874 13502
rect 17309 13499 17375 13502
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 25129 13018 25195 13021
rect 26200 13018 27000 13048
rect 25129 13016 27000 13018
rect 25129 12960 25134 13016
rect 25190 12960 27000 13016
rect 25129 12958 27000 12960
rect 25129 12955 25195 12958
rect 26200 12928 27000 12958
rect 21357 12746 21423 12749
rect 24158 12746 24164 12748
rect 21357 12744 24164 12746
rect 21357 12688 21362 12744
rect 21418 12688 24164 12744
rect 21357 12686 24164 12688
rect 21357 12683 21423 12686
rect 24158 12684 24164 12686
rect 24228 12684 24234 12748
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 14733 12474 14799 12477
rect 18413 12474 18479 12477
rect 14733 12472 18479 12474
rect 14733 12416 14738 12472
rect 14794 12416 18418 12472
rect 18474 12416 18479 12472
rect 14733 12414 18479 12416
rect 14733 12411 14799 12414
rect 18413 12411 18479 12414
rect 8845 12338 8911 12341
rect 13537 12338 13603 12341
rect 8845 12336 13603 12338
rect 8845 12280 8850 12336
rect 8906 12280 13542 12336
rect 13598 12280 13603 12336
rect 8845 12278 13603 12280
rect 8845 12275 8911 12278
rect 13537 12275 13603 12278
rect 18505 12338 18571 12341
rect 18781 12338 18847 12341
rect 18505 12336 18847 12338
rect 18505 12280 18510 12336
rect 18566 12280 18786 12336
rect 18842 12280 18847 12336
rect 18505 12278 18847 12280
rect 18505 12275 18571 12278
rect 18781 12275 18847 12278
rect 16021 12202 16087 12205
rect 18689 12202 18755 12205
rect 16021 12200 18755 12202
rect 16021 12144 16026 12200
rect 16082 12144 18694 12200
rect 18750 12144 18755 12200
rect 16021 12142 18755 12144
rect 16021 12139 16087 12142
rect 18689 12139 18755 12142
rect 24945 12202 25011 12205
rect 26200 12202 27000 12232
rect 24945 12200 27000 12202
rect 24945 12144 24950 12200
rect 25006 12144 27000 12200
rect 24945 12142 27000 12144
rect 24945 12139 25011 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 13537 11930 13603 11933
rect 16021 11930 16087 11933
rect 21357 11932 21423 11933
rect 21357 11930 21404 11932
rect 13537 11928 16087 11930
rect 13537 11872 13542 11928
rect 13598 11872 16026 11928
rect 16082 11872 16087 11928
rect 13537 11870 16087 11872
rect 21312 11928 21404 11930
rect 21312 11872 21362 11928
rect 21312 11870 21404 11872
rect 13537 11867 13603 11870
rect 16021 11867 16087 11870
rect 21357 11868 21404 11870
rect 21468 11868 21474 11932
rect 21357 11867 21423 11868
rect 13353 11794 13419 11797
rect 17769 11794 17835 11797
rect 13353 11792 17835 11794
rect 13353 11736 13358 11792
rect 13414 11736 17774 11792
rect 17830 11736 17835 11792
rect 13353 11734 17835 11736
rect 13353 11731 13419 11734
rect 17769 11731 17835 11734
rect 12341 11658 12407 11661
rect 14406 11658 14412 11660
rect 12341 11656 14412 11658
rect 12341 11600 12346 11656
rect 12402 11600 14412 11656
rect 12341 11598 14412 11600
rect 12341 11595 12407 11598
rect 14406 11596 14412 11598
rect 14476 11658 14482 11660
rect 15101 11658 15167 11661
rect 14476 11656 15167 11658
rect 14476 11600 15106 11656
rect 15162 11600 15167 11656
rect 14476 11598 15167 11600
rect 14476 11596 14482 11598
rect 15101 11595 15167 11598
rect 22461 11522 22527 11525
rect 22461 11520 22754 11522
rect 22461 11464 22466 11520
rect 22522 11464 22754 11520
rect 22461 11462 22754 11464
rect 22461 11459 22527 11462
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 13537 11252 13603 11253
rect 13486 11250 13492 11252
rect 13410 11190 13492 11250
rect 13556 11250 13603 11252
rect 15694 11250 15700 11252
rect 13556 11248 15700 11250
rect 13598 11192 15700 11248
rect 13486 11188 13492 11190
rect 13556 11190 15700 11192
rect 13556 11188 13603 11190
rect 15694 11188 15700 11190
rect 15764 11250 15770 11252
rect 16021 11250 16087 11253
rect 15764 11248 16087 11250
rect 15764 11192 16026 11248
rect 16082 11192 16087 11248
rect 15764 11190 16087 11192
rect 22694 11250 22754 11462
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 22829 11250 22895 11253
rect 22694 11248 22895 11250
rect 22694 11192 22834 11248
rect 22890 11192 22895 11248
rect 22694 11190 22895 11192
rect 15764 11188 15770 11190
rect 13537 11187 13603 11188
rect 16021 11187 16087 11190
rect 22829 11187 22895 11190
rect 11973 11114 12039 11117
rect 17217 11114 17283 11117
rect 19241 11116 19307 11117
rect 19190 11114 19196 11116
rect 11973 11112 17283 11114
rect 11973 11056 11978 11112
rect 12034 11056 17222 11112
rect 17278 11056 17283 11112
rect 11973 11054 17283 11056
rect 19150 11054 19196 11114
rect 19260 11112 19307 11116
rect 19302 11056 19307 11112
rect 11973 11051 12039 11054
rect 17217 11051 17283 11054
rect 19190 11052 19196 11054
rect 19260 11052 19307 11056
rect 19241 11051 19307 11052
rect 19517 10978 19583 10981
rect 21173 10978 21239 10981
rect 19517 10976 21239 10978
rect 19517 10920 19522 10976
rect 19578 10920 21178 10976
rect 21234 10920 21239 10976
rect 19517 10918 21239 10920
rect 19517 10915 19583 10918
rect 21173 10915 21239 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 19517 10842 19583 10845
rect 24761 10842 24827 10845
rect 19517 10840 24827 10842
rect 19517 10784 19522 10840
rect 19578 10784 24766 10840
rect 24822 10784 24827 10840
rect 19517 10782 24827 10784
rect 19517 10779 19583 10782
rect 24761 10779 24827 10782
rect 16849 10706 16915 10709
rect 19057 10706 19123 10709
rect 16849 10704 19123 10706
rect 16849 10648 16854 10704
rect 16910 10648 19062 10704
rect 19118 10648 19123 10704
rect 16849 10646 19123 10648
rect 16849 10643 16915 10646
rect 19057 10643 19123 10646
rect 11513 10570 11579 10573
rect 14549 10570 14615 10573
rect 11513 10568 14615 10570
rect 11513 10512 11518 10568
rect 11574 10512 14554 10568
rect 14610 10512 14615 10568
rect 11513 10510 14615 10512
rect 11513 10507 11579 10510
rect 14549 10507 14615 10510
rect 23381 10570 23447 10573
rect 26200 10570 27000 10600
rect 23381 10568 27000 10570
rect 23381 10512 23386 10568
rect 23442 10512 27000 10568
rect 23381 10510 27000 10512
rect 23381 10507 23447 10510
rect 26200 10480 27000 10510
rect 16941 10434 17007 10437
rect 18873 10434 18939 10437
rect 16941 10432 18939 10434
rect 16941 10376 16946 10432
rect 17002 10376 18878 10432
rect 18934 10376 18939 10432
rect 16941 10374 18939 10376
rect 16941 10371 17007 10374
rect 18873 10371 18939 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 15285 10298 15351 10301
rect 18505 10298 18571 10301
rect 15285 10296 18571 10298
rect 15285 10240 15290 10296
rect 15346 10240 18510 10296
rect 18566 10240 18571 10296
rect 15285 10238 18571 10240
rect 15285 10235 15351 10238
rect 18505 10235 18571 10238
rect 18321 10162 18387 10165
rect 18454 10162 18460 10164
rect 18321 10160 18460 10162
rect 18321 10104 18326 10160
rect 18382 10104 18460 10160
rect 18321 10102 18460 10104
rect 18321 10099 18387 10102
rect 18454 10100 18460 10102
rect 18524 10162 18530 10164
rect 18689 10162 18755 10165
rect 18524 10160 18755 10162
rect 18524 10104 18694 10160
rect 18750 10104 18755 10160
rect 18524 10102 18755 10104
rect 18524 10100 18530 10102
rect 18689 10099 18755 10102
rect 19425 10162 19491 10165
rect 20713 10162 20779 10165
rect 19425 10160 20779 10162
rect 19425 10104 19430 10160
rect 19486 10104 20718 10160
rect 20774 10104 20779 10160
rect 19425 10102 20779 10104
rect 19425 10099 19491 10102
rect 20713 10099 20779 10102
rect 16113 10026 16179 10029
rect 20161 10026 20227 10029
rect 22277 10026 22343 10029
rect 16113 10024 19442 10026
rect 16113 9968 16118 10024
rect 16174 9968 19442 10024
rect 16113 9966 19442 9968
rect 16113 9963 16179 9966
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 18689 9756 18755 9757
rect 18638 9692 18644 9756
rect 18708 9754 18755 9756
rect 18708 9752 18800 9754
rect 18750 9696 18800 9752
rect 18708 9694 18800 9696
rect 18708 9692 18755 9694
rect 18689 9691 18755 9692
rect 19382 9618 19442 9966
rect 20161 10024 22343 10026
rect 20161 9968 20166 10024
rect 20222 9968 22282 10024
rect 22338 9968 22343 10024
rect 20161 9966 22343 9968
rect 20161 9963 20227 9966
rect 22277 9963 22343 9966
rect 21633 9890 21699 9893
rect 22553 9890 22619 9893
rect 21633 9888 22619 9890
rect 21633 9832 21638 9888
rect 21694 9832 22558 9888
rect 22614 9832 22619 9888
rect 21633 9830 22619 9832
rect 21633 9827 21699 9830
rect 22553 9827 22619 9830
rect 24761 9754 24827 9757
rect 26200 9754 27000 9784
rect 24761 9752 27000 9754
rect 24761 9696 24766 9752
rect 24822 9696 27000 9752
rect 24761 9694 27000 9696
rect 24761 9691 24827 9694
rect 26200 9664 27000 9694
rect 23422 9618 23428 9620
rect 19382 9558 23428 9618
rect 23422 9556 23428 9558
rect 23492 9556 23498 9620
rect 11421 9482 11487 9485
rect 19241 9482 19307 9485
rect 11421 9480 19307 9482
rect 11421 9424 11426 9480
rect 11482 9424 19246 9480
rect 19302 9424 19307 9480
rect 11421 9422 19307 9424
rect 11421 9419 11487 9422
rect 19241 9419 19307 9422
rect 18873 9346 18939 9349
rect 19241 9346 19307 9349
rect 18873 9344 19307 9346
rect 18873 9288 18878 9344
rect 18934 9288 19246 9344
rect 19302 9288 19307 9344
rect 18873 9286 19307 9288
rect 18873 9283 18939 9286
rect 19241 9283 19307 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 10041 9074 10107 9077
rect 22553 9074 22619 9077
rect 10041 9072 22619 9074
rect 10041 9016 10046 9072
rect 10102 9016 22558 9072
rect 22614 9016 22619 9072
rect 10041 9014 22619 9016
rect 10041 9011 10107 9014
rect 22553 9011 22619 9014
rect 24945 8938 25011 8941
rect 26200 8938 27000 8968
rect 24945 8936 27000 8938
rect 24945 8880 24950 8936
rect 25006 8880 27000 8936
rect 24945 8878 27000 8880
rect 24945 8875 25011 8878
rect 26200 8848 27000 8878
rect 0 8802 800 8832
rect 3417 8802 3483 8805
rect 0 8800 3483 8802
rect 0 8744 3422 8800
rect 3478 8744 3483 8800
rect 0 8742 3483 8744
rect 0 8712 800 8742
rect 3417 8739 3483 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 15929 8530 15995 8533
rect 16982 8530 16988 8532
rect 15929 8528 16988 8530
rect 15929 8472 15934 8528
rect 15990 8472 16988 8528
rect 15929 8470 16988 8472
rect 15929 8467 15995 8470
rect 16982 8468 16988 8470
rect 17052 8468 17058 8532
rect 13813 8394 13879 8397
rect 18229 8394 18295 8397
rect 13813 8392 18295 8394
rect 13813 8336 13818 8392
rect 13874 8336 18234 8392
rect 18290 8336 18295 8392
rect 13813 8334 18295 8336
rect 13813 8331 13879 8334
rect 18229 8331 18295 8334
rect 19517 8258 19583 8261
rect 20662 8258 20668 8260
rect 19517 8256 20668 8258
rect 19517 8200 19522 8256
rect 19578 8200 20668 8256
rect 19517 8198 20668 8200
rect 19517 8195 19583 8198
rect 20662 8196 20668 8198
rect 20732 8196 20738 8260
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 17677 7986 17743 7989
rect 24945 7986 25011 7989
rect 17677 7984 25011 7986
rect 17677 7928 17682 7984
rect 17738 7928 24950 7984
rect 25006 7928 25011 7984
rect 17677 7926 25011 7928
rect 17677 7923 17743 7926
rect 24945 7923 25011 7926
rect 20437 7850 20503 7853
rect 24393 7850 24459 7853
rect 20437 7848 24459 7850
rect 20437 7792 20442 7848
rect 20498 7792 24398 7848
rect 24454 7792 24459 7848
rect 20437 7790 24459 7792
rect 20437 7787 20503 7790
rect 24393 7787 24459 7790
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 9949 7442 10015 7445
rect 23933 7442 23999 7445
rect 9949 7440 23999 7442
rect 9949 7384 9954 7440
rect 10010 7384 23938 7440
rect 23994 7384 23999 7440
rect 9949 7382 23999 7384
rect 9949 7379 10015 7382
rect 23933 7379 23999 7382
rect 15193 7306 15259 7309
rect 16430 7306 16436 7308
rect 15193 7304 16436 7306
rect 15193 7248 15198 7304
rect 15254 7248 16436 7304
rect 15193 7246 16436 7248
rect 15193 7243 15259 7246
rect 16430 7244 16436 7246
rect 16500 7306 16506 7308
rect 20713 7306 20779 7309
rect 22737 7306 22803 7309
rect 16500 7304 20779 7306
rect 16500 7248 20718 7304
rect 20774 7248 20779 7304
rect 16500 7246 20779 7248
rect 16500 7244 16506 7246
rect 20713 7243 20779 7246
rect 22694 7304 22803 7306
rect 22694 7248 22742 7304
rect 22798 7248 22803 7304
rect 22694 7243 22803 7248
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 18597 7170 18663 7173
rect 18965 7170 19031 7173
rect 18597 7168 19031 7170
rect 18597 7112 18602 7168
rect 18658 7112 18970 7168
rect 19026 7112 19031 7168
rect 18597 7110 19031 7112
rect 18597 7107 18663 7110
rect 18965 7107 19031 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22694 7037 22754 7243
rect 26200 7216 27000 7246
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 18965 7034 19031 7037
rect 19190 7034 19196 7036
rect 18965 7032 19196 7034
rect 18965 6976 18970 7032
rect 19026 6976 19196 7032
rect 18965 6974 19196 6976
rect 18965 6971 19031 6974
rect 19190 6972 19196 6974
rect 19260 6972 19266 7036
rect 22694 7032 22803 7037
rect 22694 6976 22742 7032
rect 22798 6976 22803 7032
rect 22694 6974 22803 6976
rect 22737 6971 22803 6974
rect 14365 6900 14431 6901
rect 14365 6898 14412 6900
rect 14320 6896 14412 6898
rect 14320 6840 14370 6896
rect 14320 6838 14412 6840
rect 14365 6836 14412 6838
rect 14476 6836 14482 6900
rect 14365 6835 14431 6836
rect 13445 6762 13511 6765
rect 20621 6762 20687 6765
rect 13445 6760 20687 6762
rect 13445 6704 13450 6760
rect 13506 6704 20626 6760
rect 20682 6704 20687 6760
rect 13445 6702 20687 6704
rect 13445 6699 13511 6702
rect 20621 6699 20687 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 4061 6490 4127 6493
rect 0 6488 4127 6490
rect 0 6432 4066 6488
rect 4122 6432 4127 6488
rect 0 6430 4127 6432
rect 0 6400 800 6430
rect 4061 6427 4127 6430
rect 12709 6490 12775 6493
rect 17401 6490 17467 6493
rect 12709 6488 17467 6490
rect 12709 6432 12714 6488
rect 12770 6432 17406 6488
rect 17462 6432 17467 6488
rect 12709 6430 17467 6432
rect 12709 6427 12775 6430
rect 17401 6427 17467 6430
rect 24853 6490 24919 6493
rect 26200 6490 27000 6520
rect 24853 6488 27000 6490
rect 24853 6432 24858 6488
rect 24914 6432 27000 6488
rect 24853 6430 27000 6432
rect 24853 6427 24919 6430
rect 26200 6400 27000 6430
rect 13445 6356 13511 6357
rect 13445 6354 13492 6356
rect 13400 6352 13492 6354
rect 13400 6296 13450 6352
rect 13400 6294 13492 6296
rect 13445 6292 13492 6294
rect 13556 6292 13562 6356
rect 15377 6354 15443 6357
rect 23013 6354 23079 6357
rect 15377 6352 23079 6354
rect 15377 6296 15382 6352
rect 15438 6296 23018 6352
rect 23074 6296 23079 6352
rect 15377 6294 23079 6296
rect 13445 6291 13511 6292
rect 15377 6291 15443 6294
rect 23013 6291 23079 6294
rect 10869 6218 10935 6221
rect 12985 6218 13051 6221
rect 15193 6218 15259 6221
rect 10869 6216 15259 6218
rect 10869 6160 10874 6216
rect 10930 6160 12990 6216
rect 13046 6160 15198 6216
rect 15254 6160 15259 6216
rect 10869 6158 15259 6160
rect 10869 6155 10935 6158
rect 12985 6155 13051 6158
rect 15193 6155 15259 6158
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 14181 5948 14247 5949
rect 14181 5946 14228 5948
rect 14136 5944 14228 5946
rect 14136 5888 14186 5944
rect 14136 5886 14228 5888
rect 14181 5884 14228 5886
rect 14292 5884 14298 5948
rect 14181 5883 14247 5884
rect 15469 5810 15535 5813
rect 17769 5810 17835 5813
rect 15469 5808 17835 5810
rect 15469 5752 15474 5808
rect 15530 5752 17774 5808
rect 17830 5752 17835 5808
rect 15469 5750 17835 5752
rect 15469 5747 15535 5750
rect 17769 5747 17835 5750
rect 18505 5810 18571 5813
rect 21633 5810 21699 5813
rect 23473 5812 23539 5813
rect 18505 5808 21699 5810
rect 18505 5752 18510 5808
rect 18566 5752 21638 5808
rect 21694 5752 21699 5808
rect 18505 5750 21699 5752
rect 18505 5747 18571 5750
rect 21633 5747 21699 5750
rect 23422 5748 23428 5812
rect 23492 5810 23539 5812
rect 23492 5808 23584 5810
rect 23534 5752 23584 5808
rect 23492 5750 23584 5752
rect 23492 5748 23539 5750
rect 23473 5747 23539 5748
rect 18413 5674 18479 5677
rect 23105 5674 23171 5677
rect 18413 5672 23171 5674
rect 18413 5616 18418 5672
rect 18474 5616 23110 5672
rect 23166 5616 23171 5672
rect 18413 5614 23171 5616
rect 18413 5611 18479 5614
rect 23105 5611 23171 5614
rect 23933 5674 23999 5677
rect 26200 5674 27000 5704
rect 23933 5672 27000 5674
rect 23933 5616 23938 5672
rect 23994 5616 27000 5672
rect 23933 5614 27000 5616
rect 23933 5611 23999 5614
rect 26200 5584 27000 5614
rect 21909 5538 21975 5541
rect 22369 5538 22435 5541
rect 21909 5536 22435 5538
rect 21909 5480 21914 5536
rect 21970 5480 22374 5536
rect 22430 5480 22435 5536
rect 21909 5478 22435 5480
rect 21909 5475 21975 5478
rect 22369 5475 22435 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 13077 5266 13143 5269
rect 14733 5266 14799 5269
rect 13077 5264 14799 5266
rect 13077 5208 13082 5264
rect 13138 5208 14738 5264
rect 14794 5208 14799 5264
rect 13077 5206 14799 5208
rect 13077 5203 13143 5206
rect 14733 5203 14799 5206
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23381 4858 23447 4861
rect 26200 4858 27000 4888
rect 23381 4856 27000 4858
rect 23381 4800 23386 4856
rect 23442 4800 27000 4856
rect 23381 4798 27000 4800
rect 23381 4795 23447 4798
rect 26200 4768 27000 4798
rect 16389 4722 16455 4725
rect 19425 4722 19491 4725
rect 16389 4720 19491 4722
rect 16389 4664 16394 4720
rect 16450 4664 19430 4720
rect 19486 4664 19491 4720
rect 16389 4662 19491 4664
rect 16389 4659 16455 4662
rect 19425 4659 19491 4662
rect 19609 4722 19675 4725
rect 23657 4722 23723 4725
rect 19609 4720 23723 4722
rect 19609 4664 19614 4720
rect 19670 4664 23662 4720
rect 23718 4664 23723 4720
rect 19609 4662 23723 4664
rect 19609 4659 19675 4662
rect 23657 4659 23723 4662
rect 12249 4586 12315 4589
rect 23749 4586 23815 4589
rect 12249 4584 23815 4586
rect 12249 4528 12254 4584
rect 12310 4528 23754 4584
rect 23810 4528 23815 4584
rect 12249 4526 23815 4528
rect 12249 4523 12315 4526
rect 23749 4523 23815 4526
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 0 4178 800 4208
rect 3785 4178 3851 4181
rect 0 4176 3851 4178
rect 0 4120 3790 4176
rect 3846 4120 3851 4176
rect 0 4118 3851 4120
rect 0 4088 800 4118
rect 3785 4115 3851 4118
rect 21817 4042 21883 4045
rect 26200 4042 27000 4072
rect 21817 4040 27000 4042
rect 21817 3984 21822 4040
rect 21878 3984 27000 4040
rect 21817 3982 27000 3984
rect 21817 3979 21883 3982
rect 26200 3952 27000 3982
rect 24025 3906 24091 3909
rect 24158 3906 24164 3908
rect 24025 3904 24164 3906
rect 24025 3848 24030 3904
rect 24086 3848 24164 3904
rect 24025 3846 24164 3848
rect 24025 3843 24091 3846
rect 24158 3844 24164 3846
rect 24228 3844 24234 3908
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 19006 3436 19012 3500
rect 19076 3498 19082 3500
rect 23933 3498 23999 3501
rect 19076 3496 23999 3498
rect 19076 3440 23938 3496
rect 23994 3440 23999 3496
rect 19076 3438 23999 3440
rect 19076 3436 19082 3438
rect 23933 3435 23999 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 23197 3226 23263 3229
rect 26200 3226 27000 3256
rect 23197 3224 27000 3226
rect 23197 3168 23202 3224
rect 23258 3168 27000 3224
rect 23197 3166 27000 3168
rect 23197 3163 23263 3166
rect 26200 3136 27000 3166
rect 17769 2954 17835 2957
rect 23565 2954 23631 2957
rect 17769 2952 23631 2954
rect 17769 2896 17774 2952
rect 17830 2896 23570 2952
rect 23626 2896 23631 2952
rect 17769 2894 23631 2896
rect 17769 2891 17835 2894
rect 23565 2891 23631 2894
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 22093 2410 22159 2413
rect 26200 2410 27000 2440
rect 22093 2408 27000 2410
rect 22093 2352 22098 2408
rect 22154 2352 27000 2408
rect 22093 2350 27000 2352
rect 22093 2347 22159 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 3969 1866 4035 1869
rect 0 1864 4035 1866
rect 0 1808 3974 1864
rect 4030 1808 4035 1864
rect 0 1806 4035 1808
rect 0 1776 800 1806
rect 3969 1803 4035 1806
rect 22185 1594 22251 1597
rect 26200 1594 27000 1624
rect 22185 1592 27000 1594
rect 22185 1536 22190 1592
rect 22246 1536 27000 1592
rect 22185 1534 27000 1536
rect 22185 1531 22251 1534
rect 26200 1504 27000 1534
rect 24853 778 24919 781
rect 26200 778 27000 808
rect 24853 776 27000 778
rect 24853 720 24858 776
rect 24914 720 27000 776
rect 24853 718 27000 720
rect 24853 715 24919 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 21404 38796 21468 38860
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 18460 27840 18524 27844
rect 18460 27784 18510 27840
rect 18510 27784 18524 27840
rect 18460 27780 18524 27784
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 15700 27236 15764 27300
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 17724 25604 17788 25668
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 16436 24788 16500 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 14228 23564 14292 23628
rect 19012 23428 19076 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 17172 22808 17236 22812
rect 17172 22752 17222 22808
rect 17222 22752 17236 22808
rect 17172 22748 17236 22752
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 16804 18320 16868 18324
rect 16804 18264 16854 18320
rect 16854 18264 16868 18320
rect 16804 18260 16868 18264
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 17724 17852 17788 17916
rect 20668 17852 20732 17916
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 17172 16144 17236 16148
rect 17172 16088 17222 16144
rect 17222 16088 17236 16144
rect 17172 16084 17236 16088
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 16988 15268 17052 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 20668 15132 20732 15196
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 21404 14452 21468 14516
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18644 13772 18708 13836
rect 20668 13772 20732 13836
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 16804 13500 16868 13564
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 24164 12684 24228 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 21404 11928 21468 11932
rect 21404 11872 21418 11928
rect 21418 11872 21468 11928
rect 21404 11868 21468 11872
rect 14412 11596 14476 11660
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 13492 11248 13556 11252
rect 13492 11192 13542 11248
rect 13542 11192 13556 11248
rect 13492 11188 13556 11192
rect 15700 11188 15764 11252
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 19196 11112 19260 11116
rect 19196 11056 19246 11112
rect 19246 11056 19260 11112
rect 19196 11052 19260 11056
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 18460 10100 18524 10164
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18644 9752 18708 9756
rect 18644 9696 18694 9752
rect 18694 9696 18708 9752
rect 18644 9692 18708 9696
rect 23428 9556 23492 9620
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 16988 8468 17052 8532
rect 20668 8196 20732 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 16436 7244 16500 7308
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 19196 6972 19260 7036
rect 14412 6896 14476 6900
rect 14412 6840 14426 6896
rect 14426 6840 14476 6896
rect 14412 6836 14476 6840
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 13492 6352 13556 6356
rect 13492 6296 13506 6352
rect 13506 6296 13556 6352
rect 13492 6292 13556 6296
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 14228 5944 14292 5948
rect 14228 5888 14242 5944
rect 14242 5888 14292 5944
rect 14228 5884 14292 5888
rect 23428 5808 23492 5812
rect 23428 5752 23478 5808
rect 23478 5752 23492 5808
rect 23428 5748 23492 5752
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 24164 3844 24228 3908
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 19012 3436 19076 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 21403 38860 21469 38861
rect 21403 38796 21404 38860
rect 21468 38796 21469 38860
rect 21403 38795 21469 38796
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 15699 27300 15765 27301
rect 15699 27236 15700 27300
rect 15764 27236 15765 27300
rect 15699 27235 15765 27236
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 14227 23628 14293 23629
rect 14227 23564 14228 23628
rect 14292 23564 14293 23628
rect 14227 23563 14293 23564
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 13491 11252 13557 11253
rect 13491 11188 13492 11252
rect 13556 11188 13557 11252
rect 13491 11187 13557 11188
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 13494 6357 13554 11187
rect 13491 6356 13557 6357
rect 13491 6292 13492 6356
rect 13556 6292 13557 6356
rect 13491 6291 13557 6292
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 14230 5949 14290 23563
rect 14411 11660 14477 11661
rect 14411 11596 14412 11660
rect 14476 11596 14477 11660
rect 14411 11595 14477 11596
rect 14414 6901 14474 11595
rect 15702 11253 15762 27235
rect 17944 27232 18264 28256
rect 18459 27844 18525 27845
rect 18459 27780 18460 27844
rect 18524 27780 18525 27844
rect 18459 27779 18525 27780
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17723 25668 17789 25669
rect 17723 25604 17724 25668
rect 17788 25604 17789 25668
rect 17723 25603 17789 25604
rect 16435 24852 16501 24853
rect 16435 24788 16436 24852
rect 16500 24788 16501 24852
rect 16435 24787 16501 24788
rect 15699 11252 15765 11253
rect 15699 11188 15700 11252
rect 15764 11188 15765 11252
rect 15699 11187 15765 11188
rect 16438 7309 16498 24787
rect 17171 22812 17237 22813
rect 17171 22748 17172 22812
rect 17236 22748 17237 22812
rect 17171 22747 17237 22748
rect 16803 18324 16869 18325
rect 16803 18260 16804 18324
rect 16868 18260 16869 18324
rect 16803 18259 16869 18260
rect 16806 13565 16866 18259
rect 17174 16149 17234 22747
rect 17726 17917 17786 25603
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17723 17916 17789 17917
rect 17723 17852 17724 17916
rect 17788 17852 17789 17916
rect 17723 17851 17789 17852
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17171 16148 17237 16149
rect 17171 16084 17172 16148
rect 17236 16084 17237 16148
rect 17171 16083 17237 16084
rect 16987 15332 17053 15333
rect 16987 15268 16988 15332
rect 17052 15268 17053 15332
rect 16987 15267 17053 15268
rect 16803 13564 16869 13565
rect 16803 13500 16804 13564
rect 16868 13500 16869 13564
rect 16803 13499 16869 13500
rect 16990 8533 17050 15267
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 18462 10165 18522 27779
rect 19011 23492 19077 23493
rect 19011 23428 19012 23492
rect 19076 23428 19077 23492
rect 19011 23427 19077 23428
rect 18643 13836 18709 13837
rect 18643 13772 18644 13836
rect 18708 13772 18709 13836
rect 18643 13771 18709 13772
rect 18459 10164 18525 10165
rect 18459 10100 18460 10164
rect 18524 10100 18525 10164
rect 18459 10099 18525 10100
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 18646 9757 18706 13771
rect 18643 9756 18709 9757
rect 18643 9692 18644 9756
rect 18708 9692 18709 9756
rect 18643 9691 18709 9692
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 16987 8532 17053 8533
rect 16987 8468 16988 8532
rect 17052 8468 17053 8532
rect 16987 8467 17053 8468
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 16435 7308 16501 7309
rect 16435 7244 16436 7308
rect 16500 7244 16501 7308
rect 16435 7243 16501 7244
rect 14411 6900 14477 6901
rect 14411 6836 14412 6900
rect 14476 6836 14477 6900
rect 14411 6835 14477 6836
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 14227 5948 14293 5949
rect 14227 5884 14228 5948
rect 14292 5884 14293 5948
rect 14227 5883 14293 5884
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 19014 3501 19074 23427
rect 20667 17916 20733 17917
rect 20667 17852 20668 17916
rect 20732 17852 20733 17916
rect 20667 17851 20733 17852
rect 20670 15197 20730 17851
rect 20667 15196 20733 15197
rect 20667 15132 20668 15196
rect 20732 15132 20733 15196
rect 20667 15131 20733 15132
rect 21406 14517 21466 38795
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 21403 14516 21469 14517
rect 21403 14452 21404 14516
rect 21468 14452 21469 14516
rect 21403 14451 21469 14452
rect 20667 13836 20733 13837
rect 20667 13772 20668 13836
rect 20732 13772 20733 13836
rect 20667 13771 20733 13772
rect 19195 11116 19261 11117
rect 19195 11052 19196 11116
rect 19260 11052 19261 11116
rect 19195 11051 19261 11052
rect 19198 7037 19258 11051
rect 20670 8261 20730 13771
rect 21406 11933 21466 14451
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 24163 12748 24229 12749
rect 24163 12684 24164 12748
rect 24228 12684 24229 12748
rect 24163 12683 24229 12684
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 21403 11932 21469 11933
rect 21403 11868 21404 11932
rect 21468 11868 21469 11932
rect 21403 11867 21469 11868
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 23427 9620 23493 9621
rect 23427 9556 23428 9620
rect 23492 9556 23493 9620
rect 23427 9555 23493 9556
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 20667 8260 20733 8261
rect 20667 8196 20668 8260
rect 20732 8196 20733 8260
rect 20667 8195 20733 8196
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 19195 7036 19261 7037
rect 19195 6972 19196 7036
rect 19260 6972 19261 7036
rect 19195 6971 19261 6972
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 23430 5813 23490 9555
rect 23427 5812 23493 5813
rect 23427 5748 23428 5812
rect 23492 5748 23493 5812
rect 23427 5747 23493 5748
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 24166 3909 24226 12683
rect 24163 3908 24229 3909
rect 24163 3844 24164 3908
rect 24228 3844 24229 3908
rect 24163 3843 24229 3844
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 19011 3500 19077 3501
rect 19011 3436 19012 3500
rect 19076 3436 19077 3500
rect 19011 3435 19077 3436
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15456 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_
timestamp 1679235063
transform 1 0 11040 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 1679235063
transform 1 0 18032 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _108_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1679235063
transform 1 0 21344 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _110_
timestamp 1679235063
transform 1 0 10304 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_
timestamp 1679235063
transform 1 0 24472 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_
timestamp 1679235063
transform 1 0 9660 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 1679235063
transform 1 0 9752 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1679235063
transform 1 0 25024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1679235063
transform 1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1679235063
transform 1 0 25024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1679235063
transform 1 0 21988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1679235063
transform 1 0 20792 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1679235063
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1679235063
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1679235063
transform 1 0 22172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1679235063
transform 1 0 20792 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1679235063
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1679235063
transform 1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1679235063
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 21804 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 24196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1679235063
transform 1 0 23368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1679235063
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1679235063
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1679235063
transform 1 0 5152 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 6532 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1679235063
transform 1 0 7544 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1679235063
transform 1 0 9200 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1679235063
transform 1 0 8280 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1679235063
transform 1 0 9384 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1679235063
transform 1 0 10396 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1679235063
transform 1 0 11408 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1679235063
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1679235063
transform 1 0 20424 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1679235063
transform 1 0 18400 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1679235063
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1679235063
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1679235063
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1679235063
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 22908 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 25300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1679235063
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1679235063
transform 1 0 24196 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform 1 0 25024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1679235063
transform 1 0 24012 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1679235063
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 11132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 9200 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 15272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 14168 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16284 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 15456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 15272 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 14168 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__S
timestamp 1679235063
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 15732 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__S
timestamp 1679235063
transform 1 0 14352 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15272 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__S
timestamp 1679235063
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 17296 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__S
timestamp 1679235063
transform 1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11684 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 11040 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11684 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 10120 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11316 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11132 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 8280 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 8832 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8648 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 16744 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 15732 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 15548 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 15824 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 16928 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 19320 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 19504 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1679235063
transform 1 0 25300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold11_A
timestamp 1679235063
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1679235063
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold13_A
timestamp 1679235063
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold14_A
timestamp 1679235063
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold15_A
timestamp 1679235063
transform 1 0 9476 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold16_A
timestamp 1679235063
transform 1 0 15916 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold17_A
timestamp 1679235063
transform 1 0 9108 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold18_A
timestamp 1679235063
transform 1 0 13800 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold19_A
timestamp 1679235063
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold20_A
timestamp 1679235063
transform 1 0 18124 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold21_A
timestamp 1679235063
transform 1 0 10764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold22_A
timestamp 1679235063
transform 1 0 24288 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold23_A
timestamp 1679235063
transform 1 0 24288 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold24_A
timestamp 1679235063
transform 1 0 24656 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold25_A
timestamp 1679235063
transform 1 0 24288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold26_A
timestamp 1679235063
transform 1 0 24656 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold27_A
timestamp 1679235063
transform 1 0 24288 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold28_A
timestamp 1679235063
transform 1 0 24656 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold29_A
timestamp 1679235063
transform 1 0 24656 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold30_A
timestamp 1679235063
transform 1 0 24104 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold31_A
timestamp 1679235063
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold32_A
timestamp 1679235063
transform 1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold33_A
timestamp 1679235063
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold34_A
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold37_A
timestamp 1679235063
transform 1 0 23000 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 24748 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 24748 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 24748 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 24748 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 24748 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 24748 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 24748 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 24748 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 24748 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 24748 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 22080 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 22816 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 24748 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 24748 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 5244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 7636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 8280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 8004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 3864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 24472 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 24472 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 24012 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 22632 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 25024 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 25208 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 23368 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1679235063
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1679235063
transform 1 0 22540 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform 1 0 23184 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform 1 0 24380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1679235063
transform 1 0 25300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1679235063
transform 1 0 25024 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19504 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22448 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20240 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22816 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23184 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19504 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19964 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18768 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18768 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19688 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22080 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23092 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24012 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21896 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19136 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18676 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20424 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19964 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 15456 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15640 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 11316 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13156 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15824 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15272 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15456 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16928 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18124 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17020 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19688 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19872 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22264 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22448 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22724 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19320 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19964 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19688 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_45.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22356 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_47.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_49.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 25208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16928 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16744 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 16560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16744 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 13340 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 7268 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16008 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16192 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16192 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 9016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16192 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 10304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 18676 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18492 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16192 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15088 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15272 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18032 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19044 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14720 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18492 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17848 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18032 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21160 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20976 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22448 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 25208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5060 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8188 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6532 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6532 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7636 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9292 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 7268 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6440 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7728 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9936 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 7728 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6900 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7728 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9752 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8004 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 9108 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 14996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12604 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11592 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9016 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15824 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17020 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 15088 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195
timestamp 1679235063
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15916 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13800 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 11868 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 13340 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12420 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10212 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196
timestamp 1679235063
transform 1 0 15640 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14720 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12696 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 13800 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12144 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11592 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10028 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197
timestamp 1679235063
transform 1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14812 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 9476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8648 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16376 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13248 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10580 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10212 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 15548 0 1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 12512 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 10304 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 9568 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 14628 0 -1 46784
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 11592 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 9384 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 8924 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9108 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 13432 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 10304 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 7544 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 7912 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6624 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15916 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10212 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 12604 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 10212 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 12420 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 17296 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 17204 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 19228 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 14076 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 14352 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 14628 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 15364 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 20332 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 22172 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 19872 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 22080 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp 1679235063
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1679235063
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1679235063
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1679235063
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1679235063
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1679235063
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1679235063
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1679235063
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1679235063
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1679235063
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1679235063
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1679235063
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1679235063
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263
timestamp 1679235063
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1679235063
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1679235063
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35
timestamp 1679235063
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1679235063
transform 1 0 4968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1679235063
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_72
timestamp 1679235063
transform 1 0 7728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1679235063
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1679235063
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1679235063
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1679235063
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1679235063
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1679235063
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1679235063
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1679235063
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1679235063
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1679235063
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_247
timestamp 1679235063
transform 1 0 23828 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_253
timestamp 1679235063
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1679235063
transform 1 0 24840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1679235063
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_5
timestamp 1679235063
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1679235063
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_24
timestamp 1679235063
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1679235063
transform 1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1679235063
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1679235063
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1679235063
transform 1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1679235063
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_72
timestamp 1679235063
transform 1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1679235063
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1679235063
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1679235063
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1679235063
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1679235063
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1679235063
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_183
timestamp 1679235063
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1679235063
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_235
timestamp 1679235063
transform 1 0 22724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_239
timestamp 1679235063
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1679235063
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1679235063
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1679235063
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_28
timestamp 1679235063
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1679235063
transform 1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1679235063
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1679235063
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1679235063
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1679235063
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1679235063
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1679235063
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_83
timestamp 1679235063
transform 1 0 8740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1679235063
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_104
timestamp 1679235063
transform 1 0 10672 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1679235063
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1679235063
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1679235063
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1679235063
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1679235063
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1679235063
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_231
timestamp 1679235063
transform 1 0 22356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1679235063
transform 1 0 23000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1679235063
transform 1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_252
timestamp 1679235063
transform 1 0 24288 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1679235063
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_16
timestamp 1679235063
transform 1 0 2576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1679235063
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1679235063
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_66
timestamp 1679235063
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1679235063
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1679235063
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_107
timestamp 1679235063
transform 1 0 10948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1679235063
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1679235063
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1679235063
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1679235063
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1679235063
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_192
timestamp 1679235063
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1679235063
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1679235063
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_248
timestamp 1679235063
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_259
timestamp 1679235063
transform 1 0 24932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1679235063
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 1679235063
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_68
timestamp 1679235063
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_80
timestamp 1679235063
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_92
timestamp 1679235063
transform 1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1679235063
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_120
timestamp 1679235063
transform 1 0 12144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_127
timestamp 1679235063
transform 1 0 12788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_151
timestamp 1679235063
transform 1 0 14996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1679235063
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1679235063
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1679235063
transform 1 0 17204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1679235063
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1679235063
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1679235063
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_263
timestamp 1679235063
transform 1 0 25300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1679235063
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1679235063
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1679235063
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1679235063
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_143
timestamp 1679235063
transform 1 0 14260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1679235063
transform 1 0 14536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1679235063
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1679235063
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1679235063
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1679235063
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_248
timestamp 1679235063
transform 1 0 23920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_259
timestamp 1679235063
transform 1 0 24932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_124
timestamp 1679235063
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_130
timestamp 1679235063
transform 1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1679235063
transform 1 0 14168 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1679235063
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1679235063
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_180
timestamp 1679235063
transform 1 0 17664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1679235063
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1679235063
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_247
timestamp 1679235063
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_255
timestamp 1679235063
transform 1 0 24564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_263
timestamp 1679235063
transform 1 0 25300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1679235063
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_129
timestamp 1679235063
transform 1 0 12972 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1679235063
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1679235063
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_150
timestamp 1679235063
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1679235063
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1679235063
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1679235063
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1679235063
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1679235063
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1679235063
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1679235063
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1679235063
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1679235063
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1679235063
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_130
timestamp 1679235063
transform 1 0 13064 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1679235063
transform 1 0 13616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1679235063
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1679235063
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_180
timestamp 1679235063
transform 1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_186
timestamp 1679235063
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1679235063
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1679235063
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1679235063
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1679235063
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1679235063
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1679235063
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_158
timestamp 1679235063
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_169
timestamp 1679235063
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_173
timestamp 1679235063
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1679235063
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1679235063
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_203
timestamp 1679235063
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_207
timestamp 1679235063
transform 1 0 20148 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1679235063
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_248
timestamp 1679235063
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_259
timestamp 1679235063
transform 1 0 24932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1679235063
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1679235063
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_118
timestamp 1679235063
transform 1 0 11960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_126
timestamp 1679235063
transform 1 0 12696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1679235063
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1679235063
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1679235063
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_146
timestamp 1679235063
transform 1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1679235063
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_171
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1679235063
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1679235063
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1679235063
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1679235063
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1679235063
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_111
timestamp 1679235063
transform 1 0 11316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1679235063
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1679235063
transform 1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_152
timestamp 1679235063
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_158
timestamp 1679235063
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp 1679235063
transform 1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_176
timestamp 1679235063
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_199
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_221
timestamp 1679235063
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_229
timestamp 1679235063
transform 1 0 22172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_233
timestamp 1679235063
transform 1 0 22540 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_258
timestamp 1679235063
transform 1 0 24840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_262
timestamp 1679235063
transform 1 0 25208 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1679235063
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1679235063
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1679235063
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_109
timestamp 1679235063
transform 1 0 11132 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1679235063
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1679235063
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1679235063
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1679235063
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1679235063
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1679235063
transform 1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1679235063
transform 1 0 19504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1679235063
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1679235063
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1679235063
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_261
timestamp 1679235063
transform 1 0 25116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_265
timestamp 1679235063
transform 1 0 25484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1679235063
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1679235063
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1679235063
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1679235063
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_155
timestamp 1679235063
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1679235063
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1679235063
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_174
timestamp 1679235063
transform 1 0 17112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1679235063
transform 1 0 17848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_192
timestamp 1679235063
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1679235063
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1679235063
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_231
timestamp 1679235063
transform 1 0 22356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_235
timestamp 1679235063
transform 1 0 22724 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_245
timestamp 1679235063
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1679235063
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1679235063
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1679235063
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1679235063
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1679235063
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1679235063
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_109
timestamp 1679235063
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1679235063
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_131
timestamp 1679235063
transform 1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1679235063
transform 1 0 13616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_147
timestamp 1679235063
transform 1 0 14628 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1679235063
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1679235063
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1679235063
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1679235063
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1679235063
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_230
timestamp 1679235063
transform 1 0 22264 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_234
timestamp 1679235063
transform 1 0 22632 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_237
timestamp 1679235063
transform 1 0 22908 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_259
timestamp 1679235063
transform 1 0 24932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_265
timestamp 1679235063
transform 1 0 25484 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1679235063
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1679235063
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1679235063
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1679235063
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1679235063
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1679235063
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1679235063
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_176
timestamp 1679235063
transform 1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_183
timestamp 1679235063
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1679235063
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1679235063
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1679235063
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_231
timestamp 1679235063
transform 1 0 22356 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_259
timestamp 1679235063
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1679235063
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1679235063
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1679235063
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1679235063
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1679235063
transform 1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_104
timestamp 1679235063
transform 1 0 10672 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1679235063
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1679235063
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_152
timestamp 1679235063
transform 1 0 15088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1679235063
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1679235063
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1679235063
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1679235063
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1679235063
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1679235063
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1679235063
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_71
timestamp 1679235063
transform 1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1679235063
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_87
timestamp 1679235063
transform 1 0 9108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1679235063
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1679235063
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1679235063
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_152
timestamp 1679235063
transform 1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1679235063
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_164
timestamp 1679235063
transform 1 0 16192 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1679235063
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1679235063
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1679235063
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1679235063
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1679235063
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1679235063
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1679235063
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1679235063
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_95
timestamp 1679235063
transform 1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1679235063
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1679235063
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1679235063
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1679235063
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1679235063
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1679235063
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1679235063
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_191
timestamp 1679235063
transform 1 0 18676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1679235063
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1679235063
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1679235063
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1679235063
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_234
timestamp 1679235063
transform 1 0 22632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_237
timestamp 1679235063
transform 1 0 22908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_259
timestamp 1679235063
transform 1 0 24932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1679235063
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1679235063
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1679235063
transform 1 0 8372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1679235063
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1679235063
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1679235063
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1679235063
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1679235063
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1679235063
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1679235063
transform 1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1679235063
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1679235063
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1679235063
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1679235063
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1679235063
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_218
timestamp 1679235063
transform 1 0 21160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1679235063
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_258
timestamp 1679235063
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1679235063
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1679235063
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1679235063
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1679235063
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1679235063
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1679235063
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1679235063
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_118
timestamp 1679235063
transform 1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1679235063
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1679235063
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1679235063
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1679235063
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1679235063
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1679235063
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1679235063
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1679235063
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1679235063
transform 1 0 20792 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1679235063
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_230
timestamp 1679235063
transform 1 0 22264 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_234
timestamp 1679235063
transform 1 0 22632 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1679235063
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_263
timestamp 1679235063
transform 1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1679235063
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1679235063
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1679235063
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1679235063
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1679235063
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1679235063
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1679235063
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_152
timestamp 1679235063
transform 1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_156
timestamp 1679235063
transform 1 0 15456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_164
timestamp 1679235063
transform 1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1679235063
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_183
timestamp 1679235063
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1679235063
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_205
timestamp 1679235063
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_211
timestamp 1679235063
transform 1 0 20516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1679235063
transform 1 0 21252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1679235063
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1679235063
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_261
timestamp 1679235063
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1679235063
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1679235063
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1679235063
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1679235063
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1679235063
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1679235063
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1679235063
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_107
timestamp 1679235063
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1679235063
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1679235063
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 1679235063
transform 1 0 14536 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1679235063
transform 1 0 15088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1679235063
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1679235063
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_180
timestamp 1679235063
transform 1 0 17664 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1679235063
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1679235063
transform 1 0 18952 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_200
timestamp 1679235063
transform 1 0 19504 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1679235063
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_217
timestamp 1679235063
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_221
timestamp 1679235063
transform 1 0 21436 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1679235063
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1679235063
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1679235063
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1679235063
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1679235063
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1679235063
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1679235063
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1679235063
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_100
timestamp 1679235063
transform 1 0 10304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1679235063
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1679235063
transform 1 0 12420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_127
timestamp 1679235063
transform 1 0 12788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1679235063
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1679235063
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1679235063
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_150
timestamp 1679235063
transform 1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1679235063
transform 1 0 15272 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1679235063
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1679235063
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1679235063
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_190
timestamp 1679235063
transform 1 0 18584 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1679235063
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1679235063
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_258
timestamp 1679235063
transform 1 0 24840 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1679235063
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1679235063
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1679235063
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1679235063
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1679235063
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1679235063
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1679235063
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1679235063
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1679235063
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1679235063
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1679235063
transform 1 0 11960 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1679235063
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1679235063
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1679235063
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1679235063
transform 1 0 16008 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1679235063
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1679235063
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1679235063
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1679235063
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1679235063
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1679235063
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1679235063
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_247
timestamp 1679235063
transform 1 0 23828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_253
timestamp 1679235063
transform 1 0 24380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1679235063
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1679235063
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1679235063
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1679235063
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp 1679235063
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1679235063
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1679235063
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_108
timestamp 1679235063
transform 1 0 11040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1679235063
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1679235063
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1679235063
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1679235063
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1679235063
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_172
timestamp 1679235063
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_186
timestamp 1679235063
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_190
timestamp 1679235063
transform 1 0 18584 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_199
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1679235063
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1679235063
transform 1 0 20056 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1679235063
transform 1 0 22080 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1679235063
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1679235063
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1679235063
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1679235063
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1679235063
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1679235063
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1679235063
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1679235063
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1679235063
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1679235063
transform 1 0 8464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1679235063
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1679235063
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1679235063
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1679235063
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1679235063
transform 1 0 13616 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1679235063
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1679235063
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_179
timestamp 1679235063
transform 1 0 17572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_186
timestamp 1679235063
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_210
timestamp 1679235063
transform 1 0 20424 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1679235063
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_228
timestamp 1679235063
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1679235063
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1679235063
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1679235063
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1679235063
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1679235063
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1679235063
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1679235063
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1679235063
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1679235063
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1679235063
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_143
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_155
timestamp 1679235063
transform 1 0 15364 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1679235063
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1679235063
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1679235063
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_211
timestamp 1679235063
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1679235063
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1679235063
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1679235063
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1679235063
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1679235063
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1679235063
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1679235063
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1679235063
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1679235063
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1679235063
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_92
timestamp 1679235063
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1679235063
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1679235063
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1679235063
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_134
timestamp 1679235063
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1679235063
transform 1 0 14628 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1679235063
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1679235063
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1679235063
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1679235063
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_195
timestamp 1679235063
transform 1 0 19044 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_206
timestamp 1679235063
transform 1 0 20056 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_214
timestamp 1679235063
transform 1 0 20792 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1679235063
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1679235063
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1679235063
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1679235063
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1679235063
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1679235063
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1679235063
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1679235063
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1679235063
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_95
timestamp 1679235063
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1679235063
transform 1 0 10856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_110
timestamp 1679235063
transform 1 0 11224 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1679235063
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1679235063
transform 1 0 13524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1679235063
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_146
timestamp 1679235063
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_158
timestamp 1679235063
transform 1 0 15640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_170
timestamp 1679235063
transform 1 0 16744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1679235063
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_184
timestamp 1679235063
transform 1 0 18032 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1679235063
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_217
timestamp 1679235063
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_222
timestamp 1679235063
transform 1 0 21528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_226
timestamp 1679235063
transform 1 0 21896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_230
timestamp 1679235063
transform 1 0 22264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_259
timestamp 1679235063
transform 1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1679235063
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1679235063
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1679235063
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1679235063
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1679235063
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1679235063
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1679235063
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1679235063
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_104
timestamp 1679235063
transform 1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1679235063
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_118
timestamp 1679235063
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1679235063
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_148
timestamp 1679235063
transform 1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_154
timestamp 1679235063
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1679235063
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1679235063
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_180
timestamp 1679235063
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_186
timestamp 1679235063
transform 1 0 18216 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_197
timestamp 1679235063
transform 1 0 19228 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1679235063
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1679235063
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1679235063
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1679235063
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1679235063
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1679235063
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1679235063
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1679235063
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1679235063
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1679235063
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1679235063
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1679235063
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1679235063
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1679235063
transform 1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1679235063
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1679235063
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_202
timestamp 1679235063
transform 1 0 19688 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1679235063
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_248
timestamp 1679235063
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1679235063
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_262
timestamp 1679235063
transform 1 0 25208 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1679235063
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1679235063
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1679235063
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1679235063
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 1679235063
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_95
timestamp 1679235063
transform 1 0 9844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1679235063
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1679235063
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1679235063
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1679235063
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1679235063
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1679235063
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1679235063
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1679235063
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_209
timestamp 1679235063
transform 1 0 20332 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_219
timestamp 1679235063
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1679235063
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_230
timestamp 1679235063
transform 1 0 22264 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_234
timestamp 1679235063
transform 1 0 22632 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1679235063
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1679235063
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1679235063
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1679235063
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1679235063
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1679235063
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1679235063
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1679235063
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1679235063
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_90
timestamp 1679235063
transform 1 0 9384 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1679235063
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_103
timestamp 1679235063
transform 1 0 10580 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1679235063
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_128
timestamp 1679235063
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1679235063
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1679235063
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1679235063
transform 1 0 15088 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1679235063
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1679235063
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1679235063
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1679235063
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_208
timestamp 1679235063
transform 1 0 20240 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1679235063
transform 1 0 20608 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_217
timestamp 1679235063
transform 1 0 21068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1679235063
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1679235063
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1679235063
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1679235063
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1679235063
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1679235063
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1679235063
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1679235063
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1679235063
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1679235063
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1679235063
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_118
timestamp 1679235063
transform 1 0 11960 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_150
timestamp 1679235063
transform 1 0 14904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_154
timestamp 1679235063
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1679235063
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1679235063
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1679235063
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 1679235063
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1679235063
transform 1 0 18952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_198
timestamp 1679235063
transform 1 0 19320 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1679235063
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1679235063
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_261
timestamp 1679235063
transform 1 0 25116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1679235063
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1679235063
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1679235063
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1679235063
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1679235063
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1679235063
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1679235063
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_96
timestamp 1679235063
transform 1 0 9936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1679235063
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1679235063
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_117
timestamp 1679235063
transform 1 0 11868 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_127
timestamp 1679235063
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1679235063
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1679235063
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp 1679235063
transform 1 0 16008 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_183
timestamp 1679235063
transform 1 0 17940 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1679235063
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1679235063
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1679235063
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1679235063
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1679235063
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1679235063
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_246
timestamp 1679235063
transform 1 0 23736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1679235063
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1679235063
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1679235063
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1679235063
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1679235063
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_69
timestamp 1679235063
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_75
timestamp 1679235063
transform 1 0 8004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1679235063
transform 1 0 9936 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_100
timestamp 1679235063
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1679235063
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1679235063
transform 1 0 14168 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_148
timestamp 1679235063
transform 1 0 14720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 1679235063
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_174
timestamp 1679235063
transform 1 0 17112 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_186
timestamp 1679235063
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_190
timestamp 1679235063
transform 1 0 18584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_195
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_201
timestamp 1679235063
transform 1 0 19596 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1679235063
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_211
timestamp 1679235063
transform 1 0 20516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1679235063
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1679235063
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1679235063
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1679235063
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1679235063
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1679235063
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1679235063
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1679235063
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1679235063
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_103
timestamp 1679235063
transform 1 0 10580 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_107
timestamp 1679235063
transform 1 0 10948 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_119
timestamp 1679235063
transform 1 0 12052 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1679235063
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_143
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_146
timestamp 1679235063
transform 1 0 14536 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_157
timestamp 1679235063
transform 1 0 15548 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_161
timestamp 1679235063
transform 1 0 15916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_173
timestamp 1679235063
transform 1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_181
timestamp 1679235063
transform 1 0 17756 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_191
timestamp 1679235063
transform 1 0 18676 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1679235063
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1679235063
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_216
timestamp 1679235063
transform 1 0 20976 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1679235063
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_226
timestamp 1679235063
transform 1 0 21896 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1679235063
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1679235063
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1679235063
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1679235063
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1679235063
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_69
timestamp 1679235063
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1679235063
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_99
timestamp 1679235063
transform 1 0 10212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_115
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_127
timestamp 1679235063
transform 1 0 12788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1679235063
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1679235063
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1679235063
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1679235063
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1679235063
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1679235063
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_187
timestamp 1679235063
transform 1 0 18308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_195
timestamp 1679235063
transform 1 0 19044 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1679235063
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1679235063
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1679235063
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_227
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_232
timestamp 1679235063
transform 1 0 22448 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_238
timestamp 1679235063
transform 1 0 23000 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_260
timestamp 1679235063
transform 1 0 25024 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1679235063
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1679235063
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1679235063
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1679235063
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1679235063
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1679235063
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1679235063
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_107
timestamp 1679235063
transform 1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1679235063
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_143
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_155
timestamp 1679235063
transform 1 0 15364 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1679235063
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_219
timestamp 1679235063
transform 1 0 21252 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_223
timestamp 1679235063
transform 1 0 21620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1679235063
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_259
timestamp 1679235063
transform 1 0 24932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1679235063
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1679235063
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1679235063
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1679235063
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1679235063
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1679235063
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1679235063
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1679235063
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1679235063
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_89
timestamp 1679235063
transform 1 0 9292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1679235063
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1679235063
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1679235063
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_128
timestamp 1679235063
transform 1 0 12880 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_149
timestamp 1679235063
transform 1 0 14812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1679235063
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1679235063
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1679235063
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1679235063
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1679235063
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_199
timestamp 1679235063
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1679235063
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1679235063
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_237
timestamp 1679235063
transform 1 0 22908 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_242
timestamp 1679235063
transform 1 0 23368 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1679235063
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1679235063
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1679235063
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1679235063
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1679235063
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1679235063
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1679235063
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1679235063
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1679235063
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1679235063
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1679235063
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp 1679235063
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_105
timestamp 1679235063
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_126
timestamp 1679235063
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1679235063
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1679235063
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1679235063
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_152
timestamp 1679235063
transform 1 0 15088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_156
timestamp 1679235063
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1679235063
transform 1 0 16560 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1679235063
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1679235063
transform 1 0 17848 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_188
timestamp 1679235063
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1679235063
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_199
timestamp 1679235063
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_206
timestamp 1679235063
transform 1 0 20056 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_212
timestamp 1679235063
transform 1 0 20608 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1679235063
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1679235063
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1679235063
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1679235063
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1679235063
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1679235063
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_264
timestamp 1679235063
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1679235063
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1679235063
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1679235063
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1679235063
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1679235063
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1679235063
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1679235063
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1679235063
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_89
timestamp 1679235063
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1679235063
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1679235063
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1679235063
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1679235063
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1679235063
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_129
timestamp 1679235063
transform 1 0 12972 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1679235063
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_148
timestamp 1679235063
transform 1 0 14720 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1679235063
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1679235063
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1679235063
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_174
timestamp 1679235063
transform 1 0 17112 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_178
timestamp 1679235063
transform 1 0 17480 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_190
timestamp 1679235063
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_194
timestamp 1679235063
transform 1 0 18952 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_197
timestamp 1679235063
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_209
timestamp 1679235063
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_221
timestamp 1679235063
transform 1 0 21436 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1679235063
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1679235063
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_240
timestamp 1679235063
transform 1 0 23184 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1679235063
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1679235063
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1679235063
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1679235063
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1679235063
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1679235063
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1679235063
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1679235063
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1679235063
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1679235063
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1679235063
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1679235063
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_107
timestamp 1679235063
transform 1 0 10948 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_113
timestamp 1679235063
transform 1 0 11500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_125
timestamp 1679235063
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1679235063
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1679235063
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_152
timestamp 1679235063
transform 1 0 15088 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_156
timestamp 1679235063
transform 1 0 15456 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_167
timestamp 1679235063
transform 1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1679235063
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_185
timestamp 1679235063
transform 1 0 18124 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_189
timestamp 1679235063
transform 1 0 18492 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_193
timestamp 1679235063
transform 1 0 18860 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1679235063
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_219
timestamp 1679235063
transform 1 0 21252 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1679235063
transform 1 0 21988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_232
timestamp 1679235063
transform 1 0 22448 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1679235063
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1679235063
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1679235063
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_264
timestamp 1679235063
transform 1 0 25392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1679235063
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1679235063
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1679235063
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1679235063
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1679235063
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1679235063
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1679235063
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_85
timestamp 1679235063
transform 1 0 8924 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1679235063
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_115
timestamp 1679235063
transform 1 0 11684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_127
timestamp 1679235063
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1679235063
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1679235063
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1679235063
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1679235063
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1679235063
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_203
timestamp 1679235063
transform 1 0 19780 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_207
timestamp 1679235063
transform 1 0 20148 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_219
timestamp 1679235063
transform 1 0 21252 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_225
timestamp 1679235063
transform 1 0 21804 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_228
timestamp 1679235063
transform 1 0 22080 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1679235063
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1679235063
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1679235063
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1679235063
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1679235063
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1679235063
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1679235063
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1679235063
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_65
timestamp 1679235063
transform 1 0 7084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1679235063
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_89
timestamp 1679235063
transform 1 0 9292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_101
timestamp 1679235063
transform 1 0 10396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_122
timestamp 1679235063
transform 1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_126
timestamp 1679235063
transform 1 0 12696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1679235063
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1679235063
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_162
timestamp 1679235063
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_168
timestamp 1679235063
transform 1 0 16560 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_176
timestamp 1679235063
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1679235063
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1679235063
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_197
timestamp 1679235063
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_202
timestamp 1679235063
transform 1 0 19688 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1679235063
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_248
timestamp 1679235063
transform 1 0 23920 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1679235063
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_264
timestamp 1679235063
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1679235063
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1679235063
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1679235063
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1679235063
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1679235063
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1679235063
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1679235063
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1679235063
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1679235063
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1679235063
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_105
timestamp 1679235063
transform 1 0 10764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1679235063
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1679235063
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_135
timestamp 1679235063
transform 1 0 13524 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_139
timestamp 1679235063
transform 1 0 13892 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1679235063
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_162
timestamp 1679235063
transform 1 0 16008 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1679235063
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1679235063
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_187
timestamp 1679235063
transform 1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_193
timestamp 1679235063
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_196
timestamp 1679235063
transform 1 0 19136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_200
timestamp 1679235063
transform 1 0 19504 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1679235063
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_220
timestamp 1679235063
transform 1 0 21344 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1679235063
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1679235063
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_260
timestamp 1679235063
transform 1 0 25024 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1679235063
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1679235063
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1679235063
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1679235063
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1679235063
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1679235063
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1679235063
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1679235063
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1679235063
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1679235063
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1679235063
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_111
timestamp 1679235063
transform 1 0 11316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_132
timestamp 1679235063
transform 1 0 13248 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1679235063
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1679235063
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_158
timestamp 1679235063
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_166
timestamp 1679235063
transform 1 0 16376 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1679235063
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1679235063
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1679235063
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1679235063
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_245
timestamp 1679235063
transform 1 0 23644 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1679235063
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1679235063
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1679235063
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1679235063
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1679235063
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1679235063
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1679235063
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1679235063
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1679235063
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1679235063
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1679235063
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1679235063
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1679235063
transform 1 0 9292 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1679235063
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1679235063
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_119
timestamp 1679235063
transform 1 0 12052 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_129
timestamp 1679235063
transform 1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_153
timestamp 1679235063
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1679235063
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1679235063
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1679235063
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_186
timestamp 1679235063
transform 1 0 18216 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_201
timestamp 1679235063
transform 1 0 19596 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_207
timestamp 1679235063
transform 1 0 20148 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_212
timestamp 1679235063
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_227
timestamp 1679235063
transform 1 0 21988 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1679235063
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1679235063
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_260
timestamp 1679235063
transform 1 0 25024 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1679235063
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1679235063
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1679235063
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1679235063
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1679235063
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1679235063
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1679235063
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1679235063
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1679235063
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1679235063
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1679235063
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_129
timestamp 1679235063
transform 1 0 12972 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_135
timestamp 1679235063
transform 1 0 13524 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1679235063
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1679235063
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_162
timestamp 1679235063
transform 1 0 16008 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1679235063
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1679235063
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1679235063
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1679235063
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_202
timestamp 1679235063
transform 1 0 19688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_206
timestamp 1679235063
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_216
timestamp 1679235063
transform 1 0 20976 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_228
timestamp 1679235063
transform 1 0 22080 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_238
timestamp 1679235063
transform 1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_243
timestamp 1679235063
transform 1 0 23460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1679235063
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_255
timestamp 1679235063
transform 1 0 24564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1679235063
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1679235063
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1679235063
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1679235063
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1679235063
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1679235063
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1679235063
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1679235063
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1679235063
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1679235063
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_88
timestamp 1679235063
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_100
timestamp 1679235063
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1679235063
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1679235063
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_140
timestamp 1679235063
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_152
timestamp 1679235063
transform 1 0 15088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1679235063
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_173
timestamp 1679235063
transform 1 0 17020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_185
timestamp 1679235063
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_195
timestamp 1679235063
transform 1 0 19044 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_203
timestamp 1679235063
transform 1 0 19780 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_213
timestamp 1679235063
transform 1 0 20700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1679235063
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1679235063
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1679235063
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_240
timestamp 1679235063
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_261
timestamp 1679235063
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_265
timestamp 1679235063
transform 1 0 25484 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1679235063
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1679235063
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1679235063
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1679235063
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1679235063
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1679235063
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1679235063
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1679235063
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1679235063
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1679235063
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_90
timestamp 1679235063
transform 1 0 9384 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_102
timestamp 1679235063
transform 1 0 10488 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_114
timestamp 1679235063
transform 1 0 11592 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_126
timestamp 1679235063
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1679235063
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_141
timestamp 1679235063
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_155
timestamp 1679235063
transform 1 0 15364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_161
timestamp 1679235063
transform 1 0 15916 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_169
timestamp 1679235063
transform 1 0 16652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_190
timestamp 1679235063
transform 1 0 18584 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1679235063
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1679235063
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_201
timestamp 1679235063
transform 1 0 19596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_204
timestamp 1679235063
transform 1 0 19872 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1679235063
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_233
timestamp 1679235063
transform 1 0 22540 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_241
timestamp 1679235063
transform 1 0 23276 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1679235063
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1679235063
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1679235063
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1679235063
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1679235063
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1679235063
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1679235063
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1679235063
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1679235063
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1679235063
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1679235063
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1679235063
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1679235063
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1679235063
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1679235063
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1679235063
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_125
timestamp 1679235063
transform 1 0 12604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_154
timestamp 1679235063
transform 1 0 15272 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_160
timestamp 1679235063
transform 1 0 15824 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_171
timestamp 1679235063
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_197
timestamp 1679235063
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_201
timestamp 1679235063
transform 1 0 19596 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_204
timestamp 1679235063
transform 1 0 19872 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_215
timestamp 1679235063
transform 1 0 20884 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1679235063
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1679235063
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_230
timestamp 1679235063
transform 1 0 22264 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_252
timestamp 1679235063
transform 1 0 24288 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_260
timestamp 1679235063
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1679235063
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1679235063
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1679235063
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1679235063
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1679235063
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1679235063
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1679235063
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1679235063
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1679235063
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1679235063
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1679235063
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1679235063
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1679235063
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1679235063
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1679235063
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1679235063
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1679235063
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1679235063
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_166
timestamp 1679235063
transform 1 0 16376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_190
timestamp 1679235063
transform 1 0 18584 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1679235063
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_219
timestamp 1679235063
transform 1 0 21252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_232
timestamp 1679235063
transform 1 0 22448 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_236
timestamp 1679235063
transform 1 0 22816 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_247
timestamp 1679235063
transform 1 0 23828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1679235063
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1679235063
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1679235063
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1679235063
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1679235063
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1679235063
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1679235063
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1679235063
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1679235063
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1679235063
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1679235063
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1679235063
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1679235063
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1679235063
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1679235063
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1679235063
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1679235063
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1679235063
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1679235063
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1679235063
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1679235063
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1679235063
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_174
timestamp 1679235063
transform 1 0 17112 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_186
timestamp 1679235063
transform 1 0 18216 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_190
timestamp 1679235063
transform 1 0 18584 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_193
timestamp 1679235063
transform 1 0 18860 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_215
timestamp 1679235063
transform 1 0 20884 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_221
timestamp 1679235063
transform 1 0 21436 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1679235063
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1679235063
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_263
timestamp 1679235063
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1679235063
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1679235063
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1679235063
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1679235063
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1679235063
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1679235063
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1679235063
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1679235063
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1679235063
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1679235063
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1679235063
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1679235063
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1679235063
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1679235063
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1679235063
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1679235063
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1679235063
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_166
timestamp 1679235063
transform 1 0 16376 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_174
timestamp 1679235063
transform 1 0 17112 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1679235063
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1679235063
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1679235063
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_202
timestamp 1679235063
transform 1 0 19688 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_215
timestamp 1679235063
transform 1 0 20884 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_223
timestamp 1679235063
transform 1 0 21620 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_228
timestamp 1679235063
transform 1 0 22080 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1679235063
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1679235063
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1679235063
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1679235063
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1679235063
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1679235063
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1679235063
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1679235063
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1679235063
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1679235063
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1679235063
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1679235063
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1679235063
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1679235063
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1679235063
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1679235063
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1679235063
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1679235063
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1679235063
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1679235063
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1679235063
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1679235063
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1679235063
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_193
timestamp 1679235063
transform 1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_198
timestamp 1679235063
transform 1 0 19320 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_220
timestamp 1679235063
transform 1 0 21344 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1679235063
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_247
timestamp 1679235063
transform 1 0 23828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_255
timestamp 1679235063
transform 1 0 24564 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1679235063
transform 1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1679235063
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1679235063
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1679235063
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1679235063
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1679235063
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1679235063
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1679235063
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1679235063
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1679235063
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1679235063
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1679235063
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_90
timestamp 1679235063
transform 1 0 9384 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_102
timestamp 1679235063
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1679235063
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1679235063
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1679235063
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1679235063
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_158
timestamp 1679235063
transform 1 0 15640 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_162
timestamp 1679235063
transform 1 0 16008 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_174
timestamp 1679235063
transform 1 0 17112 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1679235063
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1679235063
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1679235063
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1679235063
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1679235063
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1679235063
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_259
timestamp 1679235063
transform 1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_264
timestamp 1679235063
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1679235063
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1679235063
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1679235063
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1679235063
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1679235063
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1679235063
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1679235063
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1679235063
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1679235063
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1679235063
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1679235063
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1679235063
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1679235063
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1679235063
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1679235063
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1679235063
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1679235063
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1679235063
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1679235063
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1679235063
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1679235063
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1679235063
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_217
timestamp 1679235063
transform 1 0 21068 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1679235063
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1679235063
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1679235063
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1679235063
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_259
timestamp 1679235063
transform 1 0 24932 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1679235063
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1679235063
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1679235063
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1679235063
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1679235063
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1679235063
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1679235063
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1679235063
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1679235063
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1679235063
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1679235063
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1679235063
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1679235063
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1679235063
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1679235063
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1679235063
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1679235063
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1679235063
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1679235063
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1679235063
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1679235063
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1679235063
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1679235063
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1679235063
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1679235063
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1679235063
transform 1 0 21988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1679235063
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_244
timestamp 1679235063
transform 1 0 23552 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_253
timestamp 1679235063
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1679235063
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1679235063
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1679235063
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1679235063
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1679235063
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1679235063
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1679235063
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1679235063
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1679235063
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_81
timestamp 1679235063
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1679235063
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1679235063
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_117
timestamp 1679235063
transform 1 0 11868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_129
timestamp 1679235063
transform 1 0 12972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1679235063
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_153
timestamp 1679235063
transform 1 0 15180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1679235063
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1679235063
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1679235063
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1679235063
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1679235063
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1679235063
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1679235063
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1679235063
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_236
timestamp 1679235063
transform 1 0 22816 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_248
timestamp 1679235063
transform 1 0 23920 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_257
timestamp 1679235063
transform 1 0 24748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_264
timestamp 1679235063
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1679235063
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1679235063
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1679235063
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1679235063
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1679235063
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1679235063
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1679235063
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1679235063
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1679235063
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1679235063
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1679235063
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1679235063
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1679235063
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1679235063
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1679235063
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1679235063
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1679235063
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1679235063
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1679235063
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1679235063
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1679235063
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1679235063
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1679235063
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1679235063
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1679235063
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_245
timestamp 1679235063
transform 1 0 23644 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_249
timestamp 1679235063
transform 1 0 24012 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_253
timestamp 1679235063
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1679235063
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1679235063
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1679235063
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1679235063
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1679235063
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1679235063
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1679235063
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1679235063
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1679235063
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1679235063
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1679235063
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1679235063
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1679235063
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1679235063
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1679235063
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1679235063
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1679235063
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1679235063
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1679235063
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1679235063
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1679235063
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1679235063
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1679235063
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1679235063
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1679235063
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1679235063
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1679235063
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_249
timestamp 1679235063
transform 1 0 24012 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_254
timestamp 1679235063
transform 1 0 24472 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1679235063
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1679235063
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1679235063
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1679235063
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1679235063
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1679235063
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1679235063
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1679235063
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1679235063
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1679235063
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1679235063
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1679235063
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1679235063
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1679235063
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1679235063
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1679235063
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1679235063
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1679235063
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1679235063
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1679235063
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1679235063
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1679235063
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1679235063
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1679235063
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1679235063
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1679235063
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1679235063
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1679235063
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1679235063
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_259
timestamp 1679235063
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_264
timestamp 1679235063
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1679235063
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1679235063
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1679235063
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1679235063
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1679235063
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1679235063
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1679235063
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1679235063
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_81
timestamp 1679235063
transform 1 0 8556 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_85
timestamp 1679235063
transform 1 0 8924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_97
timestamp 1679235063
transform 1 0 10028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_109
timestamp 1679235063
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1679235063
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1679235063
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1679235063
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1679235063
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1679235063
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1679235063
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1679235063
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1679235063
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1679235063
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1679235063
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1679235063
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1679235063
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1679235063
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1679235063
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_249
timestamp 1679235063
transform 1 0 24012 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_254
timestamp 1679235063
transform 1 0 24472 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1679235063
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1679235063
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1679235063
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1679235063
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1679235063
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1679235063
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1679235063
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1679235063
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1679235063
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1679235063
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1679235063
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1679235063
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1679235063
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1679235063
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1679235063
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1679235063
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1679235063
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1679235063
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1679235063
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1679235063
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1679235063
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1679235063
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1679235063
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1679235063
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1679235063
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1679235063
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1679235063
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1679235063
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_253
timestamp 1679235063
transform 1 0 24380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_259
timestamp 1679235063
transform 1 0 24932 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1679235063
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1679235063
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1679235063
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1679235063
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1679235063
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1679235063
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1679235063
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1679235063
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1679235063
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1679235063
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1679235063
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1679235063
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1679235063
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1679235063
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1679235063
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1679235063
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1679235063
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1679235063
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1679235063
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1679235063
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1679235063
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1679235063
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1679235063
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1679235063
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1679235063
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1679235063
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1679235063
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_249
timestamp 1679235063
transform 1 0 24012 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_259
timestamp 1679235063
transform 1 0 24932 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_264
timestamp 1679235063
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1679235063
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1679235063
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1679235063
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1679235063
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1679235063
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1679235063
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1679235063
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1679235063
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1679235063
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1679235063
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1679235063
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1679235063
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1679235063
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1679235063
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1679235063
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1679235063
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1679235063
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1679235063
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1679235063
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1679235063
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1679235063
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1679235063
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1679235063
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1679235063
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1679235063
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1679235063
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1679235063
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1679235063
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_259
timestamp 1679235063
transform 1 0 24932 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1679235063
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1679235063
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1679235063
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1679235063
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1679235063
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1679235063
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1679235063
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1679235063
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1679235063
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1679235063
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1679235063
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1679235063
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1679235063
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1679235063
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1679235063
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1679235063
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1679235063
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1679235063
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1679235063
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1679235063
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1679235063
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1679235063
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1679235063
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1679235063
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1679235063
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1679235063
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1679235063
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_249
timestamp 1679235063
transform 1 0 24012 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_259
timestamp 1679235063
transform 1 0 24932 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1679235063
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1679235063
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1679235063
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1679235063
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1679235063
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1679235063
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1679235063
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1679235063
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1679235063
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1679235063
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1679235063
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1679235063
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1679235063
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1679235063
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1679235063
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1679235063
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1679235063
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1679235063
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1679235063
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1679235063
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1679235063
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1679235063
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1679235063
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1679235063
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1679235063
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1679235063
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1679235063
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1679235063
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_253
timestamp 1679235063
transform 1 0 24380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_259
timestamp 1679235063
transform 1 0 24932 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_264
timestamp 1679235063
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1679235063
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1679235063
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1679235063
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1679235063
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1679235063
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1679235063
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1679235063
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1679235063
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1679235063
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1679235063
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1679235063
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1679235063
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1679235063
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1679235063
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1679235063
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1679235063
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1679235063
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1679235063
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1679235063
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1679235063
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1679235063
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1679235063
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1679235063
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1679235063
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1679235063
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1679235063
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_249
timestamp 1679235063
transform 1 0 24012 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_255
timestamp 1679235063
transform 1 0 24564 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_258
timestamp 1679235063
transform 1 0 24840 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1679235063
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1679235063
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1679235063
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1679235063
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1679235063
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1679235063
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1679235063
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1679235063
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1679235063
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1679235063
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1679235063
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_97
timestamp 1679235063
transform 1 0 10028 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_107
timestamp 1679235063
transform 1 0 10948 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_119
timestamp 1679235063
transform 1 0 12052 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_131
timestamp 1679235063
transform 1 0 13156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1679235063
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1679235063
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1679235063
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1679235063
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1679235063
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1679235063
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1679235063
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1679235063
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1679235063
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1679235063
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1679235063
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1679235063
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1679235063
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_253
timestamp 1679235063
transform 1 0 24380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1679235063
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1679235063
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1679235063
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1679235063
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1679235063
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1679235063
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1679235063
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1679235063
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1679235063
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_81
timestamp 1679235063
transform 1 0 8556 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_89
timestamp 1679235063
transform 1 0 9292 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1679235063
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_117
timestamp 1679235063
transform 1 0 11868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_129
timestamp 1679235063
transform 1 0 12972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_141
timestamp 1679235063
transform 1 0 14076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_153
timestamp 1679235063
transform 1 0 15180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_165
timestamp 1679235063
transform 1 0 16284 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1679235063
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1679235063
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1679235063
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1679235063
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1679235063
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1679235063
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1679235063
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1679235063
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_249
timestamp 1679235063
transform 1 0 24012 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_255
timestamp 1679235063
transform 1 0 24564 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_258
timestamp 1679235063
transform 1 0 24840 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_264
timestamp 1679235063
transform 1 0 25392 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1679235063
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1679235063
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1679235063
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1679235063
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1679235063
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1679235063
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1679235063
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1679235063
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1679235063
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1679235063
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1679235063
transform 1 0 9476 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_100
timestamp 1679235063
transform 1 0 10304 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_112
timestamp 1679235063
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_124
timestamp 1679235063
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1679235063
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1679235063
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1679235063
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1679235063
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1679235063
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1679235063
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1679235063
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1679235063
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1679235063
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1679235063
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1679235063
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1679235063
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1679235063
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1679235063
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1679235063
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1679235063
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1679235063
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1679235063
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1679235063
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1679235063
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1679235063
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1679235063
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1679235063
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1679235063
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1679235063
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1679235063
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1679235063
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1679235063
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1679235063
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1679235063
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1679235063
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1679235063
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1679235063
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1679235063
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1679235063
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1679235063
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1679235063
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1679235063
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1679235063
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1679235063
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1679235063
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_249
timestamp 1679235063
transform 1 0 24012 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_254
timestamp 1679235063
transform 1 0 24472 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1679235063
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1679235063
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1679235063
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1679235063
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1679235063
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1679235063
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1679235063
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1679235063
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1679235063
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1679235063
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1679235063
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1679235063
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1679235063
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1679235063
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1679235063
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1679235063
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1679235063
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1679235063
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1679235063
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1679235063
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1679235063
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1679235063
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_197
timestamp 1679235063
transform 1 0 19228 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_207
timestamp 1679235063
transform 1 0 20148 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_229
timestamp 1679235063
transform 1 0 22172 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_241
timestamp 1679235063
transform 1 0 23276 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_249
timestamp 1679235063
transform 1 0 24012 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_253
timestamp 1679235063
transform 1 0 24380 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_259
timestamp 1679235063
transform 1 0 24932 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_264
timestamp 1679235063
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1679235063
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1679235063
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1679235063
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1679235063
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1679235063
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1679235063
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1679235063
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1679235063
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_81
timestamp 1679235063
transform 1 0 8556 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1679235063
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_101
timestamp 1679235063
transform 1 0 10396 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 1679235063
transform 1 0 11132 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_115
timestamp 1679235063
transform 1 0 11684 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_127
timestamp 1679235063
transform 1 0 12788 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_139
timestamp 1679235063
transform 1 0 13892 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_151
timestamp 1679235063
transform 1 0 14996 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_163
timestamp 1679235063
transform 1 0 16100 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1679235063
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1679235063
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1679235063
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1679235063
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1679235063
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1679235063
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1679235063
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1679235063
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1679235063
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_249
timestamp 1679235063
transform 1 0 24012 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_254
timestamp 1679235063
transform 1 0 24472 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1679235063
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1679235063
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1679235063
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1679235063
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1679235063
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1679235063
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1679235063
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1679235063
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1679235063
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1679235063
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1679235063
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_107
timestamp 1679235063
transform 1 0 10948 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_113
timestamp 1679235063
transform 1 0 11500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_125
timestamp 1679235063
transform 1 0 12604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_137
timestamp 1679235063
transform 1 0 13708 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1679235063
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1679235063
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_165
timestamp 1679235063
transform 1 0 16284 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_179
timestamp 1679235063
transform 1 0 17572 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_191
timestamp 1679235063
transform 1 0 18676 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1679235063
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1679235063
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1679235063
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1679235063
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1679235063
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1679235063
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1679235063
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_253
timestamp 1679235063
transform 1 0 24380 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_259
timestamp 1679235063
transform 1 0 24932 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1679235063
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1679235063
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1679235063
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1679235063
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1679235063
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1679235063
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1679235063
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1679235063
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1679235063
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1679235063
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1679235063
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1679235063
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1679235063
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1679235063
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_125
timestamp 1679235063
transform 1 0 12604 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_133
timestamp 1679235063
transform 1 0 13340 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_147
timestamp 1679235063
transform 1 0 14628 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_159
timestamp 1679235063
transform 1 0 15732 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1679235063
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1679235063
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1679235063
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1679235063
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1679235063
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1679235063
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1679235063
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1679235063
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1679235063
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_249
timestamp 1679235063
transform 1 0 24012 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_259
timestamp 1679235063
transform 1 0 24932 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1679235063
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1679235063
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1679235063
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1679235063
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1679235063
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1679235063
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1679235063
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1679235063
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1679235063
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1679235063
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1679235063
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1679235063
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1679235063
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_121
timestamp 1679235063
transform 1 0 12236 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_129
timestamp 1679235063
transform 1 0 12972 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1679235063
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1679235063
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1679235063
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_153
timestamp 1679235063
transform 1 0 15180 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_170
timestamp 1679235063
transform 1 0 16744 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_182
timestamp 1679235063
transform 1 0 17848 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1679235063
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1679235063
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1679235063
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1679235063
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1679235063
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1679235063
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1679235063
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1679235063
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_259
timestamp 1679235063
transform 1 0 24932 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1679235063
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1679235063
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1679235063
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1679235063
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1679235063
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1679235063
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1679235063
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1679235063
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1679235063
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1679235063
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_93
timestamp 1679235063
transform 1 0 9660 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_99
timestamp 1679235063
transform 1 0 10212 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_106
timestamp 1679235063
transform 1 0 10856 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1679235063
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1679235063
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_121
timestamp 1679235063
transform 1 0 12236 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_127
timestamp 1679235063
transform 1 0 12788 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_139
timestamp 1679235063
transform 1 0 13892 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_160
timestamp 1679235063
transform 1 0 15824 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1679235063
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1679235063
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1679235063
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1679235063
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1679235063
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1679235063
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1679235063
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1679235063
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_249
timestamp 1679235063
transform 1 0 24012 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_259
timestamp 1679235063
transform 1 0 24932 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1679235063
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1679235063
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1679235063
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1679235063
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1679235063
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1679235063
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1679235063
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1679235063
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1679235063
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1679235063
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1679235063
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1679235063
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_109
timestamp 1679235063
transform 1 0 11132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_113
timestamp 1679235063
transform 1 0 11500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_117
timestamp 1679235063
transform 1 0 11868 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_129
timestamp 1679235063
transform 1 0 12972 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1679235063
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1679235063
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1679235063
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1679235063
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1679235063
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1679235063
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1679235063
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1679235063
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1679235063
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1679235063
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1679235063
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1679235063
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1679235063
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1679235063
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_259
timestamp 1679235063
transform 1 0 24932 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_264
timestamp 1679235063
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1679235063
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1679235063
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1679235063
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1679235063
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1679235063
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1679235063
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1679235063
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1679235063
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_81
timestamp 1679235063
transform 1 0 8556 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_89
timestamp 1679235063
transform 1 0 9292 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_96
timestamp 1679235063
transform 1 0 9936 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_100
timestamp 1679235063
transform 1 0 10304 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1679235063
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1679235063
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1679235063
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1679235063
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1679235063
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1679235063
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1679235063
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1679235063
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1679235063
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1679235063
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1679235063
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1679235063
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1679235063
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1679235063
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_249
timestamp 1679235063
transform 1 0 24012 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_255
timestamp 1679235063
transform 1 0 24564 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_258
timestamp 1679235063
transform 1 0 24840 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1679235063
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1679235063
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1679235063
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1679235063
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1679235063
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1679235063
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1679235063
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1679235063
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1679235063
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1679235063
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1679235063
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_97
timestamp 1679235063
transform 1 0 10028 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_103
timestamp 1679235063
transform 1 0 10580 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_115
timestamp 1679235063
transform 1 0 11684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_127
timestamp 1679235063
transform 1 0 12788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1679235063
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1679235063
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1679235063
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1679235063
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1679235063
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1679235063
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1679235063
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1679235063
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1679235063
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1679235063
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_233
timestamp 1679235063
transform 1 0 22540 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_241
timestamp 1679235063
transform 1 0 23276 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_250
timestamp 1679235063
transform 1 0 24104 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_84_253
timestamp 1679235063
transform 1 0 24380 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1679235063
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1679235063
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1679235063
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1679235063
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1679235063
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1679235063
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1679235063
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_57
timestamp 1679235063
transform 1 0 6348 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_80
timestamp 1679235063
transform 1 0 8464 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_86
timestamp 1679235063
transform 1 0 9016 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_98
timestamp 1679235063
transform 1 0 10120 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_110
timestamp 1679235063
transform 1 0 11224 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1679235063
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1679235063
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1679235063
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1679235063
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1679235063
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1679235063
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1679235063
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1679235063
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1679235063
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1679235063
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1679235063
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1679235063
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1679235063
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1679235063
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_249
timestamp 1679235063
transform 1 0 24012 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_255
timestamp 1679235063
transform 1 0 24564 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_258
timestamp 1679235063
transform 1 0 24840 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_264
timestamp 1679235063
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1679235063
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1679235063
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1679235063
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1679235063
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1679235063
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1679235063
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1679235063
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1679235063
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1679235063
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1679235063
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_97
timestamp 1679235063
transform 1 0 10028 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_105
timestamp 1679235063
transform 1 0 10764 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_111
timestamp 1679235063
transform 1 0 11316 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_116
timestamp 1679235063
transform 1 0 11776 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_128
timestamp 1679235063
transform 1 0 12880 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1679235063
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1679235063
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1679235063
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1679235063
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1679235063
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1679235063
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1679235063
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1679235063
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1679235063
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1679235063
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_245
timestamp 1679235063
transform 1 0 23644 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_249
timestamp 1679235063
transform 1 0 24012 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_253
timestamp 1679235063
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1679235063
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1679235063
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1679235063
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1679235063
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1679235063
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1679235063
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1679235063
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1679235063
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1679235063
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1679235063
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1679235063
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1679235063
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1679235063
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1679235063
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1679235063
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1679235063
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1679235063
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1679235063
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1679235063
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1679235063
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1679235063
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1679235063
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1679235063
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1679235063
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1679235063
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1679235063
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_237
timestamp 1679235063
transform 1 0 22908 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_241
timestamp 1679235063
transform 1 0 23276 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_250
timestamp 1679235063
transform 1 0 24104 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1679235063
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1679235063
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1679235063
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1679235063
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1679235063
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1679235063
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1679235063
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_65
timestamp 1679235063
transform 1 0 7084 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_69
timestamp 1679235063
transform 1 0 7452 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_76
timestamp 1679235063
transform 1 0 8096 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_80
timestamp 1679235063
transform 1 0 8464 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_85
timestamp 1679235063
transform 1 0 8924 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_89
timestamp 1679235063
transform 1 0 9292 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_94
timestamp 1679235063
transform 1 0 9752 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_106
timestamp 1679235063
transform 1 0 10856 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_118
timestamp 1679235063
transform 1 0 11960 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_130
timestamp 1679235063
transform 1 0 13064 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_138
timestamp 1679235063
transform 1 0 13800 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1679235063
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1679235063
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1679235063
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1679235063
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1679235063
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1679235063
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1679235063
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1679235063
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1679235063
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1679235063
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1679235063
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1679235063
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_253
timestamp 1679235063
transform 1 0 24380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_88_263
timestamp 1679235063
transform 1 0 25300 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1679235063
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1679235063
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1679235063
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1679235063
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1679235063
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1679235063
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1679235063
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1679235063
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1679235063
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1679235063
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1679235063
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1679235063
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1679235063
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1679235063
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1679235063
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1679235063
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1679235063
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1679235063
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1679235063
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1679235063
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1679235063
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1679235063
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1679235063
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1679235063
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1679235063
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1679235063
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_249
timestamp 1679235063
transform 1 0 24012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_253
timestamp 1679235063
transform 1 0 24380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_256
timestamp 1679235063
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1679235063
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1679235063
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1679235063
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1679235063
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1679235063
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1679235063
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1679235063
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_65
timestamp 1679235063
transform 1 0 7084 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_69
timestamp 1679235063
transform 1 0 7452 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_74
timestamp 1679235063
transform 1 0 7912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1679235063
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_85
timestamp 1679235063
transform 1 0 8924 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_91
timestamp 1679235063
transform 1 0 9476 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_103
timestamp 1679235063
transform 1 0 10580 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_115
timestamp 1679235063
transform 1 0 11684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_127
timestamp 1679235063
transform 1 0 12788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1679235063
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1679235063
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1679235063
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1679235063
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1679235063
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1679235063
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1679235063
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1679235063
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1679235063
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1679235063
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1679235063
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1679235063
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1679235063
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_253
timestamp 1679235063
transform 1 0 24380 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_256
timestamp 1679235063
transform 1 0 24656 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1679235063
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1679235063
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1679235063
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1679235063
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1679235063
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1679235063
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1679235063
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1679235063
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1679235063
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1679235063
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1679235063
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1679235063
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1679235063
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1679235063
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1679235063
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1679235063
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1679235063
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1679235063
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1679235063
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1679235063
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1679235063
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1679235063
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1679235063
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1679235063
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1679235063
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1679235063
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1679235063
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_251
timestamp 1679235063
transform 1 0 24196 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_256
timestamp 1679235063
transform 1 0 24656 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1679235063
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1679235063
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1679235063
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1679235063
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1679235063
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1679235063
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_53
timestamp 1679235063
transform 1 0 5980 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_62
timestamp 1679235063
transform 1 0 6808 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_74
timestamp 1679235063
transform 1 0 7912 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1679235063
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1679235063
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1679235063
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1679235063
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1679235063
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1679235063
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1679235063
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1679235063
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1679235063
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1679235063
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1679235063
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1679235063
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1679235063
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1679235063
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1679235063
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1679235063
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1679235063
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_245
timestamp 1679235063
transform 1 0 23644 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_250
timestamp 1679235063
transform 1 0 24104 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_255
timestamp 1679235063
transform 1 0 24564 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1679235063
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1679235063
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1679235063
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1679235063
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_39
timestamp 1679235063
transform 1 0 4692 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_43
timestamp 1679235063
transform 1 0 5060 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1679235063
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1679235063
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1679235063
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1679235063
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1679235063
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1679235063
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1679235063
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1679235063
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1679235063
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1679235063
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1679235063
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1679235063
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1679235063
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1679235063
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1679235063
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1679235063
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1679235063
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1679235063
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1679235063
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1679235063
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_225
timestamp 1679235063
transform 1 0 21804 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_233
timestamp 1679235063
transform 1 0 22540 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_236
timestamp 1679235063
transform 1 0 22816 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_244
timestamp 1679235063
transform 1 0 23552 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_250
timestamp 1679235063
transform 1 0 24104 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1679235063
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1679235063
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1679235063
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1679235063
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1679235063
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_47
timestamp 1679235063
transform 1 0 5428 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_59
timestamp 1679235063
transform 1 0 6532 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_76
timestamp 1679235063
transform 1 0 8096 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1679235063
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_97
timestamp 1679235063
transform 1 0 10028 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1679235063
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_133
timestamp 1679235063
transform 1 0 13340 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_137
timestamp 1679235063
transform 1 0 13708 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1679235063
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_151
timestamp 1679235063
transform 1 0 14996 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_158
timestamp 1679235063
transform 1 0 15640 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_170
timestamp 1679235063
transform 1 0 16744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_174
timestamp 1679235063
transform 1 0 17112 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_183
timestamp 1679235063
transform 1 0 17940 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_187
timestamp 1679235063
transform 1 0 18308 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1679235063
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1679235063
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1679235063
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_221
timestamp 1679235063
transform 1 0 21436 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_229
timestamp 1679235063
transform 1 0 22172 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_234
timestamp 1679235063
transform 1 0 22632 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1679235063
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1679235063
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_253
timestamp 1679235063
transform 1 0 24380 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1679235063
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1679235063
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1679235063
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1679235063
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1679235063
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1679235063
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1679235063
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1679235063
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1679235063
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1679235063
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_85
timestamp 1679235063
transform 1 0 8924 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_89
timestamp 1679235063
transform 1 0 9292 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_106
timestamp 1679235063
transform 1 0 10856 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1679235063
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_119
timestamp 1679235063
transform 1 0 12052 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_136
timestamp 1679235063
transform 1 0 13616 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_141
timestamp 1679235063
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_146
timestamp 1679235063
transform 1 0 14536 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_150
timestamp 1679235063
transform 1 0 14904 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_159
timestamp 1679235063
transform 1 0 15732 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_163
timestamp 1679235063
transform 1 0 16100 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1679235063
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_179
timestamp 1679235063
transform 1 0 17572 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_191
timestamp 1679235063
transform 1 0 18676 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1679235063
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_209
timestamp 1679235063
transform 1 0 20332 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_217
timestamp 1679235063
transform 1 0 21068 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_221
timestamp 1679235063
transform 1 0 21436 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1679235063
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_231
timestamp 1679235063
transform 1 0 22356 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_235
timestamp 1679235063
transform 1 0 22724 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_240
timestamp 1679235063
transform 1 0 23184 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1679235063
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_253
timestamp 1679235063
transform 1 0 24380 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1679235063
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold2
timestamp 1679235063
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 24656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold6
timestamp 1679235063
transform 1 0 17388 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 3956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 23368 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 23368 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 24656 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 24656 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 24656 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 16836 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7820 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 14996 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold17
timestamp 1679235063
transform 1 0 7452 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 14260 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold19
timestamp 1679235063
transform 1 0 7176 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 17940 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold21
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 24656 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 24656 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 24656 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 24656 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 24656 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 24656 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 24656 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 24656 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 23368 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 6624 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 6348 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 1932 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 24656 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 24656 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 24564 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 24380 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 25116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 24472 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1679235063
transform 1 0 25024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1679235063
transform 1 0 25024 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 25116 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1679235063
transform 1 0 25024 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1679235063
transform 1 0 25024 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1679235063
transform 1 0 25024 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1679235063
transform 1 0 25024 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1679235063
transform 1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 25116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1679235063
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1679235063
transform 1 0 25024 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1679235063
transform 1 0 25024 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1679235063
transform 1 0 24472 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 23828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 23184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1679235063
transform 1 0 5152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1679235063
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1679235063
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1679235063
transform 1 0 7820 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1679235063
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1679235063
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1679235063
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1679235063
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1679235063
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 11040 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1679235063
transform 1 0 2116 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1679235063
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1679235063
transform 1 0 3404 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1679235063
transform 1 0 5152 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 14260 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1679235063
transform 1 0 15364 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1679235063
transform 1 0 16836 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 17664 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 19412 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1679235063
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24840 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1679235063
transform 1 0 24840 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1679235063
transform 1 0 24840 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 25024 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1679235063
transform 1 0 22264 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1679235063
transform 1 0 23736 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1679235063
transform 1 0 24472 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1679235063
transform 1 0 23000 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1679235063
transform 1 0 20700 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1679235063
transform 1 0 21988 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1679235063
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1679235063
transform 1 0 23736 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 17480 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 1564 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 22632 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 22632 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 9752 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 22080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 22080 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 23920 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 18216 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 20056 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 12328 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 23828 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 21712 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 21252 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 17480 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 15272 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 17296 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 20240 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 20056 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 12052 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 3956 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 6624 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform 1 0 9384 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform 1 0 10764 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 12144 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1679235063
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1679235063
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1679235063
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1679235063
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1679235063
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1679235063
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1679235063
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1679235063
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1679235063
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1679235063
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1679235063
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1679235063
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1679235063
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1679235063
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1679235063
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1679235063
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1679235063
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1679235063
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1679235063
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1679235063
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1679235063
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1679235063
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1679235063
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1679235063
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1679235063
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1679235063
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1679235063
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1679235063
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1679235063
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1679235063
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1679235063
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1679235063
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1679235063
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1679235063
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1679235063
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1679235063
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1679235063
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1679235063
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1679235063
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1679235063
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1679235063
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1679235063
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1679235063
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1679235063
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1679235063
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1679235063
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1679235063
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1679235063
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1679235063
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1679235063
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1679235063
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1679235063
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1679235063
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1679235063
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1679235063
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1679235063
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1679235063
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1679235063
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1679235063
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1679235063
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1679235063
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1679235063
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1679235063
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1679235063
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1679235063
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1679235063
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1679235063
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1679235063
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1679235063
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1679235063
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1679235063
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1679235063
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1679235063
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1679235063
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1679235063
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1679235063
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1679235063
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1679235063
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1679235063
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1679235063
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1679235063
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1679235063
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1679235063
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1679235063
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1679235063
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1679235063
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1679235063
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1679235063
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1679235063
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1679235063
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1679235063
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1679235063
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1679235063
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1679235063
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1679235063
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1679235063
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1679235063
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1679235063
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1679235063
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1679235063
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1679235063
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1679235063
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1679235063
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1679235063
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1679235063
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1679235063
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1679235063
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1679235063
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1679235063
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1679235063
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18584 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19872 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22080 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23276 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21528 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21896 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23184 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23552 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23552 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23184 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22080 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19872 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17940 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17020 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16744 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16744 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17388 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20700 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22448 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23276 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23460 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21620 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19504 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19044 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20608 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23460 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20332 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13340 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9108 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10488 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9292 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11132 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11776 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11408 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13340 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13064 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12972 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10856 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8096 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6624 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10672 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12328 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12696 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12512 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11776 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9108 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9016 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10764 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15180 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16100 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16376 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14904 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13156 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13892 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15088 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15916 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19596 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20516 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20424 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20240 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23092 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22632 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22080 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19504 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19596 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18492 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17296 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__198
timestamp 1679235063
transform 1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19504 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20056 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__160
timestamp 1679235063
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22172 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19228 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__162
timestamp 1679235063
transform 1 0 19688 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19504 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22632 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 21988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20240 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__199
timestamp 1679235063
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__200
timestamp 1679235063
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19596 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__201
timestamp 1679235063
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__202
timestamp 1679235063
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20148 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__151
timestamp 1679235063
transform 1 0 18216 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17756 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20056 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17480 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__152
timestamp 1679235063
transform 1 0 18032 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21620 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__154
timestamp 1679235063
transform 1 0 19688 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23000 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22356 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__156
timestamp 1679235063
transform 1 0 24748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22724 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__157
timestamp 1679235063
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__158
timestamp 1679235063
transform 1 0 20056 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19872 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__159
timestamp 1679235063
transform 1 0 19412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18768 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23552 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22264 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__161
timestamp 1679235063
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19964 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12144 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__164
timestamp 1679235063
transform 1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14812 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15180 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9200 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__170
timestamp 1679235063
transform 1 0 9936 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12144 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15456 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10672 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__181
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13524 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15272 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__192
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15640 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13248 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__193
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11224 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__165
timestamp 1679235063
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9936 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 7820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__166
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11500 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15732 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__167
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__168
timestamp 1679235063
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14536 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__169
timestamp 1679235063
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__171
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__172
timestamp 1679235063
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__173
timestamp 1679235063
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__174
timestamp 1679235063
transform 1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20148 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__175
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13708 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19780 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__176
timestamp 1679235063
transform 1 0 15456 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17848 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__177
timestamp 1679235063
transform 1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__178
timestamp 1679235063
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21528 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13340 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__179
timestamp 1679235063
transform 1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14720 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__180
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__182
timestamp 1679235063
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23092 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__183
timestamp 1679235063
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__184
timestamp 1679235063
transform 1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18032 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19596 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19688 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18768 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__185
timestamp 1679235063
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__186
timestamp 1679235063
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21436 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__187
timestamp 1679235063
transform 1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__188
timestamp 1679235063
transform -1 0 12144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20516 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__189
timestamp 1679235063
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17940 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__190
timestamp 1679235063
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17388 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__191
timestamp 1679235063
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1679235063
transform 1 0 11040 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1679235063
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1679235063
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1679235063
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1679235063
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1679235063
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1679235063
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1679235063
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1679235063
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1679235063
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1679235063
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1679235063
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1679235063
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1679235063
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1679235063
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1679235063
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1679235063
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1679235063
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1679235063
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1679235063
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1679235063
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1679235063
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1679235063
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1679235063
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1679235063
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1679235063
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1679235063
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1679235063
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1679235063
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1679235063
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1679235063
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1679235063
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1679235063
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1679235063
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1679235063
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1679235063
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1679235063
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1679235063
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1679235063
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1679235063
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1679235063
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1679235063
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1679235063
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1679235063
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1679235063
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1679235063
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1679235063
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1679235063
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1679235063
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1679235063
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1679235063
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1679235063
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1679235063
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1679235063
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1679235063
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1679235063
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1679235063
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1679235063
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1679235063
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1679235063
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1679235063
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1679235063
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1679235063
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1679235063
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1679235063
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1679235063
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1679235063
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1679235063
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1679235063
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1679235063
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1679235063
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1679235063
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1679235063
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1679235063
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1679235063
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1679235063
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1679235063
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1679235063
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1679235063
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1679235063
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1679235063
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1679235063
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1679235063
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1679235063
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1679235063
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1679235063
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1679235063
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1679235063
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1679235063
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1679235063
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1679235063
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1679235063
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1679235063
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1679235063
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1679235063
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1679235063
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1679235063
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1679235063
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1679235063
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1679235063
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1679235063
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1679235063
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1679235063
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1679235063
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1679235063
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1679235063
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1679235063
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1679235063
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1679235063
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1679235063
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1679235063
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1679235063
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1679235063
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1679235063
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1679235063
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1679235063
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1679235063
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1679235063
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1679235063
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1679235063
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1679235063
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1679235063
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1679235063
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1679235063
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1679235063
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1679235063
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1679235063
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1679235063
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1679235063
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1679235063
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1679235063
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1679235063
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1679235063
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1679235063
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1679235063
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1679235063
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1679235063
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1679235063
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1679235063
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1679235063
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1679235063
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1679235063
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1679235063
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1679235063
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1679235063
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1679235063
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1679235063
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1679235063
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1679235063
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1679235063
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1679235063
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1679235063
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1679235063
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1679235063
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1679235063
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1679235063
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1679235063
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1679235063
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1679235063
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1679235063
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1679235063
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1679235063
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1679235063
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1679235063
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1679235063
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 25870 56200 25926 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1030 56200 1086 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 3790 56200 3846 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 6550 56200 6606 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 14830 56200 14886 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 17590 56200 17646 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 20350 56200 20406 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 23110 56200 23166 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable
port 158 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 9890 35598 9890 35598 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 9706 30906 9706 30906 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9292 42670 9292 42670 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 9154 44302 9154 44302 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 8280 37978 8280 37978 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 8418 16218 8418 16218 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 15778 12750 15778 12750 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 9338 12750 9338 12750 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 9660 15538 9660 15538 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 8050 14586 8050 14586 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 14858 14484 14858 14484 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13570 10098 13570 10098 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 9706 13362 9706 13362 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 8510 21318 8510 21318 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 16376 10574 16376 10574 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 13202 12784 13202 12784 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 13294 18836 13294 18836 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 9936 17714 9936 17714 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 12742 15980 12742 15980 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 10902 21522 10902 21522 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal2 12098 9520 12098 9520 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9200 15674 9200 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9062 30702 9062 30702 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 13938 9826 13938 9826 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14582 10387 14582 10387 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13432 12682 13432 12682 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9660 12954 9660 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11132 14994 11132 14994 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10994 12410 10994 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9154 12954 9154 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10258 12954 10258 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 10166 17238 10166 17238 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 15870 8500 15870 8500 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9016 13498 9016 13498 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 7774 17850 7774 17850 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 16330 8330 16330 8330 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15134 10234 15134 10234 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15318 13158 15318 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14352 14246 14352 14246 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 10718 10574 10718 10574 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10626 11696 10626 11696 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9798 11866 9798 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11592 13158 11592 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8924 16626 8924 16626 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13294 12954 13294 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10304 20570 10304 20570 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9292 33966 9292 33966 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14306 12886 14306 12886 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13432 14314 13432 14314 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12650 11832 12650 11832 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 11638 16456 11638 16456 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12650 17170 12650 17170 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12880 18666 12880 18666 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 10258 18394 10258 18394 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 13662 23222 13662 23222 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 12742 20298 12742 20298 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14030 15334 14030 15334 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10442 26520 10442 26520 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9200 29274 9200 29274 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13294 16150 13294 16150 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12926 11866 12926 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12604 14484 12604 14484 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 13846 18564 13846 18564 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12190 18768 12190 18768 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11362 15674 11362 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10488 23630 10488 23630 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 13846 24752 13846 24752 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10350 21658 10350 21658 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 10718 43146 10718 43146 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 11040 44166 11040 44166 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 11224 49130 11224 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 15766 44778 15766 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9568 44778 9568 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 10212 42670 10212 42670 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 10396 49130 10396 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 15640 45866 15640 45866 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 10212 45050 10212 45050 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 9200 44370 9200 44370 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 9568 50218 9568 50218 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 13662 46818 13662 46818 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 7912 50422 7912 50422 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 8510 48756 8510 48756 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal2 13754 46750 13754 46750 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25300 54162 25300 54162 0 ccff_head
rlabel metal2 1518 2064 1518 2064 0 ccff_head_0
rlabel metal3 25630 748 25630 748 0 ccff_tail
rlabel metal1 1564 53618 1564 53618 0 ccff_tail_0
rlabel metal1 25024 25262 25024 25262 0 chanx_right_in[0]
rlabel metal2 25346 34391 25346 34391 0 chanx_right_in[10]
rlabel metal1 24794 35054 24794 35054 0 chanx_right_in[11]
rlabel metal1 24472 36142 24472 36142 0 chanx_right_in[12]
rlabel metal1 24840 36754 24840 36754 0 chanx_right_in[13]
rlabel metal1 24794 37842 24794 37842 0 chanx_right_in[14]
rlabel metal1 24840 38726 24840 38726 0 chanx_right_in[15]
rlabel metal2 25346 39253 25346 39253 0 chanx_right_in[16]
rlabel metal2 25346 39967 25346 39967 0 chanx_right_in[17]
rlabel metal2 25346 40613 25346 40613 0 chanx_right_in[18]
rlabel metal1 24794 41582 24794 41582 0 chanx_right_in[19]
rlabel metal1 25392 24174 25392 24174 0 chanx_right_in[1]
rlabel metal1 24840 42330 24840 42330 0 chanx_right_in[20]
rlabel metal1 24840 43282 24840 43282 0 chanx_right_in[21]
rlabel metal2 24702 44183 24702 44183 0 chanx_right_in[22]
rlabel metal1 25392 45458 25392 45458 0 chanx_right_in[23]
rlabel metal2 25346 45781 25346 45781 0 chanx_right_in[24]
rlabel metal2 25346 46495 25346 46495 0 chanx_right_in[25]
rlabel metal2 25346 47141 25346 47141 0 chanx_right_in[26]
rlabel metal1 24794 48110 24794 48110 0 chanx_right_in[27]
rlabel metal1 24840 48858 24840 48858 0 chanx_right_in[28]
rlabel metal1 24518 49402 24518 49402 0 chanx_right_in[29]
rlabel metal2 24058 27013 24058 27013 0 chanx_right_in[2]
rlabel metal1 24564 29478 24564 29478 0 chanx_right_in[3]
rlabel metal1 23414 29580 23414 29580 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel via2 25530 30923 25530 30923 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal1 24840 33286 24840 33286 0 chanx_right_in[8]
rlabel metal2 25346 33677 25346 33677 0 chanx_right_in[9]
rlabel metal2 22218 2057 22218 2057 0 chanx_right_out[0]
rlabel metal2 24794 9061 24794 9061 0 chanx_right_out[10]
rlabel metal3 24894 10540 24894 10540 0 chanx_right_out[11]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[12]
rlabel metal3 25676 12172 25676 12172 0 chanx_right_out[13]
rlabel metal3 25768 12988 25768 12988 0 chanx_right_out[14]
rlabel metal2 23874 13549 23874 13549 0 chanx_right_out[15]
rlabel metal1 24380 14450 24380 14450 0 chanx_right_out[16]
rlabel metal2 23322 15249 23322 15249 0 chanx_right_out[17]
rlabel metal2 24794 15589 24794 15589 0 chanx_right_out[18]
rlabel metal2 23874 16813 23874 16813 0 chanx_right_out[19]
rlabel metal2 22126 2091 22126 2091 0 chanx_right_out[1]
rlabel metal1 24380 17714 24380 17714 0 chanx_right_out[20]
rlabel metal1 24104 18326 24104 18326 0 chanx_right_out[21]
rlabel metal1 23460 18802 23460 18802 0 chanx_right_out[22]
rlabel metal2 24702 19261 24702 19261 0 chanx_right_out[23]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[24]
rlabel metal3 24848 21964 24848 21964 0 chanx_right_out[25]
rlabel metal3 25630 22780 25630 22780 0 chanx_right_out[26]
rlabel metal2 25162 23137 25162 23137 0 chanx_right_out[27]
rlabel metal3 25124 24412 25124 24412 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal1 21850 3672 21850 3672 0 chanx_right_out[2]
rlabel metal2 21850 6749 21850 6749 0 chanx_right_out[3]
rlabel metal2 20654 5916 20654 5916 0 chanx_right_out[4]
rlabel metal3 25170 5644 25170 5644 0 chanx_right_out[5]
rlabel metal3 25630 6460 25630 6460 0 chanx_right_out[6]
rlabel metal1 24104 7446 24104 7446 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal3 25676 8908 25676 8908 0 chanx_right_out[9]
rlabel metal2 1886 1588 1886 1588 0 chany_bottom_in_0[0]
rlabel metal1 5842 2278 5842 2278 0 chany_bottom_in_0[10]
rlabel metal1 5658 4114 5658 4114 0 chany_bottom_in_0[11]
rlabel metal1 5980 3502 5980 3502 0 chany_bottom_in_0[12]
rlabel metal2 6670 891 6670 891 0 chany_bottom_in_0[13]
rlabel metal1 7682 3536 7682 3536 0 chany_bottom_in_0[14]
rlabel metal1 7452 4454 7452 4454 0 chany_bottom_in_0[15]
rlabel metal1 7820 3026 7820 3026 0 chany_bottom_in_0[16]
rlabel metal2 8142 1367 8142 1367 0 chany_bottom_in_0[17]
rlabel metal2 8510 1761 8510 1761 0 chany_bottom_in_0[18]
rlabel metal1 5796 2822 5796 2822 0 chany_bottom_in_0[19]
rlabel metal2 2254 2132 2254 2132 0 chany_bottom_in_0[1]
rlabel metal1 10212 4114 10212 4114 0 chany_bottom_in_0[20]
rlabel metal1 9338 2890 9338 2890 0 chany_bottom_in_0[21]
rlabel metal2 7958 2587 7958 2587 0 chany_bottom_in_0[22]
rlabel metal1 9568 1802 9568 1802 0 chany_bottom_in_0[23]
rlabel metal1 10074 3502 10074 3502 0 chany_bottom_in_0[24]
rlabel metal1 10212 1734 10212 1734 0 chany_bottom_in_0[25]
rlabel metal2 11730 3468 11730 3468 0 chany_bottom_in_0[26]
rlabel metal1 9890 2992 9890 2992 0 chany_bottom_in_0[27]
rlabel metal2 12190 1656 12190 1656 0 chany_bottom_in_0[28]
rlabel metal2 12558 3740 12558 3740 0 chany_bottom_in_0[29]
rlabel metal1 2392 2958 2392 2958 0 chany_bottom_in_0[2]
rlabel metal1 2484 2482 2484 2482 0 chany_bottom_in_0[3]
rlabel metal1 3496 3026 3496 3026 0 chany_bottom_in_0[4]
rlabel metal1 3496 4046 3496 4046 0 chany_bottom_in_0[5]
rlabel metal1 4002 3910 4002 3910 0 chany_bottom_in_0[6]
rlabel metal1 4048 3502 4048 3502 0 chany_bottom_in_0[7]
rlabel metal1 4462 3570 4462 3570 0 chany_bottom_in_0[8]
rlabel metal1 4968 2958 4968 2958 0 chany_bottom_in_0[9]
rlabel metal2 12926 1231 12926 1231 0 chany_bottom_out_0[0]
rlabel metal1 17894 2890 17894 2890 0 chany_bottom_out_0[10]
rlabel metal1 22632 2414 22632 2414 0 chany_bottom_out_0[11]
rlabel metal2 17342 1435 17342 1435 0 chany_bottom_out_0[12]
rlabel metal1 18814 2822 18814 2822 0 chany_bottom_out_0[13]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out_0[14]
rlabel metal2 18446 1435 18446 1435 0 chany_bottom_out_0[15]
rlabel metal2 18814 1231 18814 1231 0 chany_bottom_out_0[16]
rlabel metal1 19550 5746 19550 5746 0 chany_bottom_out_0[17]
rlabel metal1 20470 3366 20470 3366 0 chany_bottom_out_0[18]
rlabel metal2 19918 1520 19918 1520 0 chany_bottom_out_0[19]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out_0[1]
rlabel metal2 20286 1010 20286 1010 0 chany_bottom_out_0[20]
rlabel metal2 20654 1520 20654 1520 0 chany_bottom_out_0[21]
rlabel metal2 21022 1761 21022 1761 0 chany_bottom_out_0[22]
rlabel metal2 21390 1761 21390 1761 0 chany_bottom_out_0[23]
rlabel metal1 21528 6222 21528 6222 0 chany_bottom_out_0[24]
rlabel metal2 22126 823 22126 823 0 chany_bottom_out_0[25]
rlabel metal1 22540 8398 22540 8398 0 chany_bottom_out_0[26]
rlabel metal2 22862 823 22862 823 0 chany_bottom_out_0[27]
rlabel metal2 23230 1656 23230 1656 0 chany_bottom_out_0[28]
rlabel metal2 17802 3451 17802 3451 0 chany_bottom_out_0[29]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out_0[2]
rlabel metal1 14398 3570 14398 3570 0 chany_bottom_out_0[3]
rlabel metal2 14398 1622 14398 1622 0 chany_bottom_out_0[4]
rlabel metal1 15042 2958 15042 2958 0 chany_bottom_out_0[5]
rlabel metal1 16238 2822 16238 2822 0 chany_bottom_out_0[6]
rlabel metal1 16054 3570 16054 3570 0 chany_bottom_out_0[7]
rlabel metal1 16606 2958 16606 2958 0 chany_bottom_out_0[8]
rlabel metal1 16790 4046 16790 4046 0 chany_bottom_out_0[9]
rlabel metal1 20148 13294 20148 13294 0 clknet_0_prog_clk
rlabel metal1 9798 14382 9798 14382 0 clknet_4_0_0_prog_clk
rlabel metal1 6670 48790 6670 48790 0 clknet_4_10_0_prog_clk
rlabel metal2 16790 32062 16790 32062 0 clknet_4_11_0_prog_clk
rlabel metal1 18170 20570 18170 20570 0 clknet_4_12_0_prog_clk
rlabel metal2 23046 21794 23046 21794 0 clknet_4_13_0_prog_clk
rlabel metal1 19090 32266 19090 32266 0 clknet_4_14_0_prog_clk
rlabel metal1 20700 34034 20700 34034 0 clknet_4_15_0_prog_clk
rlabel metal2 13478 13600 13478 13600 0 clknet_4_1_0_prog_clk
rlabel metal1 9706 17646 9706 17646 0 clknet_4_2_0_prog_clk
rlabel metal1 12788 21522 12788 21522 0 clknet_4_3_0_prog_clk
rlabel metal1 15548 5678 15548 5678 0 clknet_4_4_0_prog_clk
rlabel metal1 20378 12274 20378 12274 0 clknet_4_5_0_prog_clk
rlabel metal1 17986 16660 17986 16660 0 clknet_4_6_0_prog_clk
rlabel metal1 20056 19890 20056 19890 0 clknet_4_7_0_prog_clk
rlabel metal2 13386 29648 13386 29648 0 clknet_4_8_0_prog_clk
rlabel metal1 16146 28526 16146 28526 0 clknet_4_9_0_prog_clk
rlabel metal1 2484 54094 2484 54094 0 gfpga_pad_io_soc_dir[0]
rlabel metal1 4140 53618 4140 53618 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 5198 55158 5198 55158 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 6578 54920 6578 54920 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 13662 53754 13662 53754 0 gfpga_pad_io_soc_in[0]
rlabel metal1 14950 54162 14950 54162 0 gfpga_pad_io_soc_in[1]
rlabel metal1 16330 54298 16330 54298 0 gfpga_pad_io_soc_in[2]
rlabel metal2 17802 56236 17802 56236 0 gfpga_pad_io_soc_in[3]
rlabel metal2 7958 55711 7958 55711 0 gfpga_pad_io_soc_out[0]
rlabel metal1 9614 54094 9614 54094 0 gfpga_pad_io_soc_out[1]
rlabel metal1 10718 53652 10718 53652 0 gfpga_pad_io_soc_out[2]
rlabel metal2 12282 56236 12282 56236 0 gfpga_pad_io_soc_out[3]
rlabel metal1 19228 54162 19228 54162 0 isol_n
rlabel metal2 24610 51034 24610 51034 0 net1
rlabel metal1 24656 39270 24656 39270 0 net10
rlabel metal2 22126 22780 22126 22780 0 net100
rlabel metal1 22908 20570 22908 20570 0 net101
rlabel metal1 23920 22610 23920 22610 0 net102
rlabel metal1 20838 25160 20838 25160 0 net103
rlabel metal2 22862 25636 22862 25636 0 net104
rlabel metal2 13202 4352 13202 4352 0 net105
rlabel metal1 19205 3706 19205 3706 0 net106
rlabel metal1 13800 5882 13800 5882 0 net107
rlabel metal1 21206 13362 21206 13362 0 net108
rlabel via1 13386 5253 13386 5253 0 net109
rlabel metal1 24242 40154 24242 40154 0 net11
rlabel metal1 24150 15946 24150 15946 0 net110
rlabel metal2 9982 6035 9982 6035 0 net111
rlabel metal2 10074 6647 10074 6647 0 net112
rlabel metal1 17526 14008 17526 14008 0 net113
rlabel metal1 18952 3026 18952 3026 0 net114
rlabel metal1 21022 2618 21022 2618 0 net115
rlabel metal1 18998 4114 18998 4114 0 net116
rlabel metal2 19642 2587 19642 2587 0 net117
rlabel metal2 19458 4097 19458 4097 0 net118
rlabel metal1 12604 4590 12604 4590 0 net119
rlabel metal1 25300 40358 25300 40358 0 net12
rlabel metal1 21022 3502 21022 3502 0 net120
rlabel metal1 20332 5678 20332 5678 0 net121
rlabel metal1 24932 18666 24932 18666 0 net122
rlabel metal1 21988 4590 21988 4590 0 net123
rlabel metal1 13248 2482 13248 2482 0 net124
rlabel metal2 21574 2958 21574 2958 0 net125
rlabel metal2 21298 6018 21298 6018 0 net126
rlabel metal2 17710 8449 17710 8449 0 net127
rlabel metal1 15916 6766 15916 6766 0 net128
rlabel metal1 20332 6290 20332 6290 0 net129
rlabel metal3 23161 38828 23161 38828 0 net13
rlabel metal2 17526 3876 17526 3876 0 net130
rlabel metal2 22310 5780 22310 5780 0 net131
rlabel via2 20470 7837 20470 7837 0 net132
rlabel metal1 20286 8398 20286 8398 0 net133
rlabel metal2 12282 4335 12282 4335 0 net134
rlabel metal1 16560 17034 16560 17034 0 net135
rlabel metal3 17089 15300 17089 15300 0 net136
rlabel metal1 14122 2414 14122 2414 0 net137
rlabel metal1 14766 3026 14766 3026 0 net138
rlabel metal1 16836 2414 16836 2414 0 net139
rlabel metal2 23414 23528 23414 23528 0 net14
rlabel metal1 16836 3502 16836 3502 0 net140
rlabel metal1 17572 13158 17572 13158 0 net141
rlabel metal1 17572 13294 17572 13294 0 net142
rlabel metal1 4646 53210 4646 53210 0 net143
rlabel metal1 5382 52666 5382 52666 0 net144
rlabel metal2 4830 52768 4830 52768 0 net145
rlabel metal1 8556 51510 8556 51510 0 net146
rlabel metal1 7866 51578 7866 51578 0 net147
rlabel metal2 9614 52326 9614 52326 0 net148
rlabel metal2 10718 51442 10718 51442 0 net149
rlabel metal2 16606 14484 16606 14484 0 net15
rlabel metal2 11730 51748 11730 51748 0 net150
rlabel metal1 18262 26010 18262 26010 0 net151
rlabel metal1 18032 27438 18032 27438 0 net152
rlabel metal1 24656 15538 24656 15538 0 net153
rlabel metal2 19734 28288 19734 28288 0 net154
rlabel metal1 22724 26962 22724 26962 0 net155
rlabel metal2 24978 28798 24978 28798 0 net156
rlabel metal1 21850 30226 21850 30226 0 net157
rlabel metal1 20194 30362 20194 30362 0 net158
rlabel metal2 19182 29376 19182 29376 0 net159
rlabel metal1 24886 42772 24886 42772 0 net16
rlabel metal1 21942 19346 21942 19346 0 net160
rlabel metal1 21988 17170 21988 17170 0 net161
rlabel metal1 19688 22746 19688 22746 0 net162
rlabel metal2 22034 21250 22034 21250 0 net163
rlabel metal1 7636 17306 7636 17306 0 net164
rlabel metal1 7222 12274 7222 12274 0 net165
rlabel metal2 8234 12546 8234 12546 0 net166
rlabel metal1 13478 17646 13478 17646 0 net167
rlabel metal2 13202 17408 13202 17408 0 net168
rlabel metal1 15732 16218 15732 16218 0 net169
rlabel via3 16859 18292 16859 18292 0 net17
rlabel metal2 9982 21250 9982 21250 0 net170
rlabel metal1 13524 10710 13524 10710 0 net171
rlabel metal2 12650 7616 12650 7616 0 net172
rlabel metal1 15410 7854 15410 7854 0 net173
rlabel metal1 17296 14314 17296 14314 0 net174
rlabel metal1 14214 15130 14214 15130 0 net175
rlabel metal1 15824 16422 15824 16422 0 net176
rlabel metal1 15870 15130 15870 15130 0 net177
rlabel metal2 13386 8126 13386 8126 0 net178
rlabel metal1 14766 4658 14766 4658 0 net179
rlabel metal1 25208 45254 25208 45254 0 net18
rlabel metal1 15318 5814 15318 5814 0 net180
rlabel metal1 11408 21658 11408 21658 0 net181
rlabel metal3 19412 9792 19412 9792 0 net182
rlabel metal1 21988 9486 21988 9486 0 net183
rlabel metal2 18446 11968 18446 11968 0 net184
rlabel metal1 18952 12274 18952 12274 0 net185
rlabel metal2 20010 11390 20010 11390 0 net186
rlabel metal2 22770 5627 22770 5627 0 net187
rlabel metal2 14214 4896 14214 4896 0 net188
rlabel metal1 21114 3162 21114 3162 0 net189
rlabel metal2 25116 40732 25116 40732 0 net19
rlabel metal1 21574 2346 21574 2346 0 net190
rlabel metal1 11592 7854 11592 7854 0 net191
rlabel metal2 11730 19584 11730 19584 0 net192
rlabel metal2 9430 17408 9430 17408 0 net193
rlabel metal1 10948 12954 10948 12954 0 net194
rlabel metal1 13018 10030 13018 10030 0 net195
rlabel metal1 15410 23086 15410 23086 0 net196
rlabel metal1 15640 25874 15640 25874 0 net197
rlabel metal1 20332 21522 20332 21522 0 net198
rlabel metal1 23230 21896 23230 21896 0 net199
rlabel metal1 1610 4692 1610 4692 0 net2
rlabel metal2 21206 41072 21206 41072 0 net20
rlabel metal1 23552 21998 23552 21998 0 net200
rlabel metal1 20792 23154 20792 23154 0 net201
rlabel metal2 18538 24650 18538 24650 0 net202
rlabel metal1 24932 3366 24932 3366 0 net203
rlabel metal2 22126 4624 22126 4624 0 net204
rlabel metal2 24610 3706 24610 3706 0 net205
rlabel metal1 18814 2380 18814 2380 0 net206
rlabel metal1 23782 3706 23782 3706 0 net207
rlabel metal1 18952 17850 18952 17850 0 net208
rlabel metal1 1978 3536 1978 3536 0 net209
rlabel metal1 25852 47158 25852 47158 0 net21
rlabel metal1 5014 4522 5014 4522 0 net210
rlabel metal2 24702 53754 24702 53754 0 net211
rlabel metal2 24058 45900 24058 45900 0 net212
rlabel metal1 24426 25466 24426 25466 0 net213
rlabel metal1 25024 36006 25024 36006 0 net214
rlabel metal2 25346 35462 25346 35462 0 net215
rlabel metal2 17066 53754 17066 53754 0 net216
rlabel metal1 13018 31994 13018 31994 0 net217
rlabel metal2 15594 53754 15594 53754 0 net218
rlabel metal1 12420 37910 12420 37910 0 net219
rlabel via2 17250 16099 17250 16099 0 net22
rlabel metal1 14720 53754 14720 53754 0 net220
rlabel metal1 9292 27370 9292 27370 0 net221
rlabel metal1 18262 53550 18262 53550 0 net222
rlabel metal1 12282 39610 12282 39610 0 net223
rlabel metal2 25346 37026 25346 37026 0 net224
rlabel metal2 25346 38114 25346 38114 0 net225
rlabel metal2 25162 42398 25162 42398 0 net226
rlabel metal2 25346 43554 25346 43554 0 net227
rlabel metal1 25254 41174 25254 41174 0 net228
rlabel metal2 25346 44642 25346 44642 0 net229
rlabel metal1 18216 17850 18216 17850 0 net23
rlabel metal2 25162 47838 25162 47838 0 net230
rlabel metal2 25162 48926 25162 48926 0 net231
rlabel metal1 24288 49742 24288 49742 0 net232
rlabel metal1 6670 3162 6670 3162 0 net233
rlabel metal2 7038 3910 7038 3910 0 net234
rlabel metal1 7452 2618 7452 2618 0 net235
rlabel metal2 2944 2516 2944 2516 0 net236
rlabel metal1 2208 3706 2208 3706 0 net237
rlabel metal1 3726 4590 3726 4590 0 net238
rlabel metal1 23414 54196 23414 54196 0 net239
rlabel metal1 24794 49844 24794 49844 0 net24
rlabel metal2 24610 52700 24610 52700 0 net240
rlabel metal2 23414 49130 23414 49130 0 net241
rlabel metal1 25300 20910 25300 20910 0 net25
rlabel metal1 25392 23086 25392 23086 0 net26
rlabel metal2 22494 27744 22494 27744 0 net27
rlabel metal1 23000 26282 23000 26282 0 net28
rlabel metal1 25116 26282 25116 26282 0 net29
rlabel metal3 20125 15164 20125 15164 0 net3
rlabel metal1 25116 31926 25116 31926 0 net30
rlabel metal1 24380 33626 24380 33626 0 net31
rlabel metal1 24702 33830 24702 33830 0 net32
rlabel metal2 1702 2176 1702 2176 0 net33
rlabel metal1 14306 14450 14306 14450 0 net34
rlabel metal2 12282 13396 12282 13396 0 net35
rlabel metal2 6578 5134 6578 5134 0 net36
rlabel metal2 5842 3774 5842 3774 0 net37
rlabel metal2 7498 7956 7498 7956 0 net38
rlabel metal1 13800 14926 13800 14926 0 net39
rlabel metal1 25116 31994 25116 31994 0 net4
rlabel metal1 14812 13158 14812 13158 0 net40
rlabel metal1 14122 13362 14122 13362 0 net41
rlabel metal1 13478 7956 13478 7956 0 net42
rlabel metal1 7866 4012 7866 4012 0 net43
rlabel metal1 5336 16966 5336 16966 0 net44
rlabel metal1 13800 5542 13800 5542 0 net45
rlabel metal2 14306 7582 14306 7582 0 net46
rlabel metal2 15686 2315 15686 2315 0 net47
rlabel metal2 14950 2689 14950 2689 0 net48
rlabel metal1 18906 12886 18906 12886 0 net49
rlabel metal1 22034 17748 22034 17748 0 net5
rlabel metal1 17526 8364 17526 8364 0 net50
rlabel metal2 21114 13226 21114 13226 0 net51
rlabel metal1 15778 8806 15778 8806 0 net52
rlabel metal1 16192 7718 16192 7718 0 net53
rlabel metal1 14674 8806 14674 8806 0 net54
rlabel metal2 2438 9826 2438 9826 0 net55
rlabel metal1 6348 2550 6348 2550 0 net56
rlabel metal1 10764 19142 10764 19142 0 net57
rlabel metal2 2530 3774 2530 3774 0 net58
rlabel metal2 4186 7514 4186 7514 0 net59
rlabel metal1 24564 35462 24564 35462 0 net6
rlabel metal1 8096 12750 8096 12750 0 net60
rlabel metal1 13892 18598 13892 18598 0 net61
rlabel metal1 12926 17102 12926 17102 0 net62
rlabel metal1 13938 53958 13938 53958 0 net63
rlabel metal1 15088 53414 15088 53414 0 net64
rlabel metal1 16284 53414 16284 53414 0 net65
rlabel metal1 17112 44914 17112 44914 0 net66
rlabel metal1 18170 54196 18170 54196 0 net67
rlabel metal1 21390 3536 21390 3536 0 net68
rlabel metal1 25024 50694 25024 50694 0 net69
rlabel metal1 25484 37298 25484 37298 0 net7
rlabel metal1 25576 51306 25576 51306 0 net70
rlabel metal2 17618 32164 17618 32164 0 net71
rlabel metal2 25254 49674 25254 49674 0 net72
rlabel metal1 20148 20910 20148 20910 0 net73
rlabel metal2 20102 21760 20102 21760 0 net74
rlabel metal1 21160 20434 21160 20434 0 net75
rlabel metal1 17848 19278 17848 19278 0 net76
rlabel metal1 20608 20842 20608 20842 0 net77
rlabel metal2 20194 21726 20194 21726 0 net78
rlabel metal1 21206 20570 21206 20570 0 net79
rlabel metal1 25576 38182 25576 38182 0 net8
rlabel metal1 17848 19210 17848 19210 0 net80
rlabel metal1 18768 14994 18768 14994 0 net81
rlabel metal1 1794 53516 1794 53516 0 net82
rlabel metal1 15272 6290 15272 6290 0 net83
rlabel metal1 15686 8534 15686 8534 0 net84
rlabel metal1 23092 11118 23092 11118 0 net85
rlabel metal1 24288 9146 24288 9146 0 net86
rlabel metal1 23966 11322 23966 11322 0 net87
rlabel metal1 24564 11730 24564 11730 0 net88
rlabel metal1 22862 13328 22862 13328 0 net89
rlabel metal1 25116 38726 25116 38726 0 net9
rlabel metal1 24288 13498 24288 13498 0 net90
rlabel metal2 22034 13974 22034 13974 0 net91
rlabel metal1 24380 12410 24380 12410 0 net92
rlabel metal1 22034 13804 22034 13804 0 net93
rlabel metal1 12926 4454 12926 4454 0 net94
rlabel metal2 24610 17204 24610 17204 0 net95
rlabel metal2 22126 18428 22126 18428 0 net96
rlabel metal1 23736 18734 23736 18734 0 net97
rlabel metal1 23046 20264 23046 20264 0 net98
rlabel metal1 22678 20978 22678 20978 0 net99
rlabel metal2 18906 23970 18906 23970 0 prog_clk
rlabel metal1 24518 4114 24518 4114 0 prog_reset
rlabel metal1 25024 50898 25024 50898 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 24978 51323 24978 51323 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24978 52275 24978 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel via2 25530 52955 25530 52955 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 23828 53006 23828 53006 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 24932 53210 24932 53210 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25860 55420 25860 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 23437 56100 23437 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 20562 56236 20562 56236 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21896 54162 21896 54162 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 23138 55711 23138 55711 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 24150 52462 24150 52462 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 22310 34918 22310 34918 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21988 34918 21988 34918 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 21298 35734 21298 35734 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 19136 21658 19136 21658 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 18768 13838 18768 13838 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal1 21160 19278 21160 19278 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal1 20056 19754 20056 19754 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 22862 21454 22862 21454 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel viali 25254 22073 25254 22073 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal1 25024 23834 25024 23834 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal2 22402 27608 22402 27608 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal1 25162 27540 25162 27540 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 20700 26418 20700 26418 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal1 23552 28594 23552 28594 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal1 19366 26758 19366 26758 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal2 22586 27438 22586 27438 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal1 18768 29818 18768 29818 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal2 18906 29172 18906 29172 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal1 18124 31858 18124 31858 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal1 17795 31994 17795 31994 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal2 25162 19924 25162 19924 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal1 24058 20026 24058 20026 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal2 21022 29614 21022 29614 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal1 20976 31858 20976 31858 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal1 23552 30294 23552 30294 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal1 23322 31790 23322 31790 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal1 25208 32538 25208 32538 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal1 24518 32334 24518 32334 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal1 23414 33422 23414 33422 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal1 22356 33422 22356 33422 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 20654 33286 20654 33286 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel metal1 23322 33830 23322 33830 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 20884 32198 20884 32198 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal2 21206 33082 21206 33082 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal1 22954 21658 22954 21658 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 25392 20570 25392 20570 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 23966 29070 23966 29070 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 20838 24378 20838 24378 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal1 20240 23630 20240 23630 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 22218 24752 22218 24752 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal1 10994 26418 10994 26418 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal1 19044 33082 19044 33082 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal1 13662 29818 13662 29818 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal1 12558 22032 12558 22032 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 8832 19142 8832 19142 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal2 14858 25126 14858 25126 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 6900 19278 6900 19278 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal2 10902 19244 10902 19244 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 8510 18598 8510 18598 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 13754 21454 13754 21454 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal1 12926 21114 12926 21114 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal2 14490 19754 14490 19754 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal1 14996 21454 14996 21454 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal1 14352 16694 14352 16694 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal1 14214 19142 14214 19142 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal1 11132 26894 11132 26894 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal1 15778 27948 15778 27948 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal1 9476 26894 9476 26894 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal1 12926 10540 12926 10540 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal1 10718 11186 10718 11186 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal1 12834 7276 12834 7276 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel metal2 10994 7514 10994 7514 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal1 12650 6834 12650 6834 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal1 11592 5882 11592 5882 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal1 17066 14484 17066 14484 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel metal1 14260 12750 14260 12750 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 17434 19244 17434 19244 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 15081 20026 15081 20026 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal2 17158 21182 17158 21182 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal1 18032 22066 18032 22066 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal1 18676 18802 18676 18802 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal2 18630 20893 18630 20893 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal2 16698 9282 16698 9282 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal1 17572 18802 17572 18802 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal1 16192 5338 16192 5338 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal1 13938 6290 13938 6290 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 16376 5610 16376 5610 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 15410 5202 15410 5202 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 13662 28594 13662 28594 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal1 15962 29682 15962 29682 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal1 13616 30022 13616 30022 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal1 19136 6630 19136 6630 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal1 17572 6698 17572 6698 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal1 21022 10574 21022 10574 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal1 21298 9146 21298 9146 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal1 20930 15334 20930 15334 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal1 19826 20978 19826 20978 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal1 21620 16014 21620 16014 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 20010 12750 20010 12750 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal1 22770 12886 22770 12886 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal1 21850 20366 21850 20366 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal2 23414 10268 23414 10268 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal1 21390 12716 21390 12716 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal1 23828 7718 23828 7718 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal2 22402 8483 22402 8483 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal2 21298 4964 21298 4964 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal1 21298 7276 21298 7276 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal1 19780 7310 19780 7310 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel metal1 19313 7174 19313 7174 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal2 19090 9248 19090 9248 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal1 13846 24038 13846 24038 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal1 14536 29274 14536 29274 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal1 15870 26860 15870 26860 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal2 14766 25024 14766 25024 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal2 12926 23970 12926 23970 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal1 17894 14790 17894 14790 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 20654 19482 20654 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20010 19482 20010 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19458 19142 19458 19142 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16974 11118 16974 11118 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 24978 22066 24978 22066 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 15028 21022 15028 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19826 17646 19826 17646 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 23046 24786 23046 24786 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19550 17714 19550 17714 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17572 9350 17572 9350 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal1 21436 23834 21436 23834 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 17578 20056 17578 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19136 10166 19136 10166 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal1 19596 24038 19596 24038 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18308 16082 18308 16082 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21298 3026 21298 3026 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal1 18952 25942 18952 25942 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16606 22406 16606 22406 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 14398 6851 14398 6851 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal1 18952 27370 18952 27370 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 19346 16284 19346 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21298 7412 21298 7412 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal2 25070 19380 25070 19380 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22402 10642 22402 10642 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17388 18156 17388 18156 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal1 21252 31926 21252 31926 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19320 19822 19320 19822 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 20907 13804 20907 13804 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal1 22908 31926 22908 31926 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21298 18292 21298 18292 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20608 18598 20608 18598 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal2 24932 32572 24932 32572 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 18700 21482 18700 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19550 20230 19550 20230 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal1 22632 34918 22632 34918 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20148 20434 20148 20434 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 17986 10676 17986 10676 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal1 21344 35530 21344 35530 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19228 20434 19228 20434 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15548 21318 15548 21318 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 19780 35530 19780 35530 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15732 21522 15732 21522 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21298 13838 21298 13838 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 23092 19482 23092 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21252 13906 21252 13906 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13340 5678 13340 5678 0 sb_0__8_.mux_bottom_track_51.out
rlabel metal2 22770 17680 22770 17680 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21022 12988 21022 12988 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22080 3026 22080 3026 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal1 20838 23086 20838 23086 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19918 23290 19918 23290 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18216 17238 18216 17238 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20056 14246 20056 14246 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 22540 21658 22540 21658 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21988 18972 21988 18972 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21758 25330 21758 25330 0 sb_0__8_.mux_right_track_0.out
rlabel metal1 14122 32742 14122 32742 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14076 31926 14076 31926 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12236 24786 12236 24786 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7682 17068 7682 17068 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14674 24616 14674 24616 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 21022 21148 21022 21148 0 sb_0__8_.mux_right_track_10.out
rlabel metal2 11730 24310 11730 24310 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14306 23137 14306 23137 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10626 18394 10626 18394 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7222 12954 7222 12954 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14122 19448 14122 19448 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16974 19788 16974 19788 0 sb_0__8_.mux_right_track_12.out
rlabel metal1 12052 18666 12052 18666 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9614 12614 9614 12614 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 19312 12558 19312 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18722 21216 18722 21216 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 15456 22134 15456 22134 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15226 19822 15226 19822 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17733 21522 17733 21522 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18998 19448 18998 19448 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 15732 20570 15732 20570 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14122 16966 14122 16966 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18170 20264 18170 20264 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18906 16422 18906 16422 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 14812 16218 14812 16218 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17733 16558 17733 16558 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 25296 21022 25296 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 14168 27438 14168 27438 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13616 27370 13616 27370 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12650 26656 12650 26656 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12650 21403 12650 21403 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13846 25976 13846 25976 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19734 13328 19734 13328 0 sb_0__8_.mux_right_track_20.out
rlabel metal2 12834 11016 12834 11016 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18308 12818 18308 12818 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17526 10778 17526 10778 0 sb_0__8_.mux_right_track_22.out
rlabel metal1 10810 6426 10810 6426 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 9401 12466 9401 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22034 12767 22034 12767 0 sb_0__8_.mux_right_track_24.out
rlabel metal2 12834 7106 12834 7106 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14582 8058 14582 8058 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23414 13634 23414 13634 0 sb_0__8_.mux_right_track_26.out
rlabel metal1 14398 12954 14398 12954 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19642 14076 19642 14076 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25254 16014 25254 16014 0 sb_0__8_.mux_right_track_28.out
rlabel metal1 17112 23494 17112 23494 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17250 19686 17250 19686 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20010 18768 20010 18768 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20930 17544 20930 17544 0 sb_0__8_.mux_right_track_30.out
rlabel metal1 17940 19890 17940 19890 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17480 19754 17480 19754 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21114 17680 21114 17680 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21804 15334 21804 15334 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 18492 18598 18492 18598 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18768 18666 18768 18666 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19918 18870 19918 18870 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22494 10098 22494 10098 0 sb_0__8_.mux_right_track_34.out
rlabel metal1 16974 18598 16974 18598 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12972 7718 12972 7718 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20194 11458 20194 11458 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13524 6630 13524 6630 0 sb_0__8_.mux_right_track_36.out
rlabel metal1 15364 6426 15364 6426 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15318 6154 15318 6154 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 6834 12558 6834 0 sb_0__8_.mux_right_track_38.out
rlabel metal2 14766 6256 14766 6256 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 5202 12926 5202 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22310 24582 22310 24582 0 sb_0__8_.mux_right_track_4.out
rlabel metal1 15640 29274 15640 29274 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15962 29614 15962 29614 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15410 29002 15410 29002 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13984 24820 13984 24820 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17710 25262 17710 25262 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10166 3162 10166 3162 0 sb_0__8_.mux_right_track_40.out
rlabel metal2 17802 6528 17802 6528 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17250 3094 17250 3094 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12834 5457 12834 5457 0 sb_0__8_.mux_right_track_42.out
rlabel metal2 21206 10829 21206 10829 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19090 10574 19090 10574 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24564 16014 24564 16014 0 sb_0__8_.mux_right_track_44.out
rlabel metal1 19780 21046 19780 21046 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18078 11832 18078 11832 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22172 14858 22172 14858 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23500 9350 23500 9350 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 20562 21930 20562 21930 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19366 12614 19366 12614 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20746 15776 20746 15776 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21390 13005 21390 13005 0 sb_0__8_.mux_right_track_48.out
rlabel metal1 21022 20298 21022 20298 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20746 11254 20746 11254 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21988 14518 21988 14518 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13754 5644 13754 5644 0 sb_0__8_.mux_right_track_50.out
rlabel metal1 21574 12614 21574 12614 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18630 5389 18630 5389 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18400 3570 18400 3570 0 sb_0__8_.mux_right_track_52.out
rlabel metal2 19550 10268 19550 10268 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 2074 21988 2074 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21298 2108 21298 2108 0 sb_0__8_.mux_right_track_54.out
rlabel metal1 20884 4046 20884 4046 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 2414 21022 2414 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14030 4896 14030 4896 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 18492 5746 18492 5746 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18262 3417 18262 3417 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24656 3162 24656 3162 0 sb_0__8_.mux_right_track_58.out
rlabel metal1 17388 12954 17388 12954 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11546 8058 11546 8058 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20148 12886 20148 12886 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21206 22032 21206 22032 0 sb_0__8_.mux_right_track_6.out
rlabel metal1 16192 27030 16192 27030 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 27098 16284 27098 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 25296 14950 25296 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14536 23698 14536 23698 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 23732 18262 23732 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 16882 22882 16882 22882 0 sb_0__8_.mux_right_track_8.out
rlabel metal2 13754 25500 13754 25500 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13984 23766 13984 23766 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12650 22134 12650 22134 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8740 17306 8740 17306 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16192 22610 16192 22610 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
