magic
tech sky130A
magscale 1 2
timestamp 1625785872
<< locali >>
rect 17417 13175 17451 13277
rect 15577 12835 15611 12937
rect 8401 12631 8435 12733
rect 18981 12495 19015 13413
rect 11529 11679 11563 11849
rect 18981 11271 19015 12257
rect 8769 7735 8803 7905
<< viali >>
rect 2697 14569 2731 14603
rect 4077 14569 4111 14603
rect 8033 14569 8067 14603
rect 1869 14501 1903 14535
rect 2237 14501 2271 14535
rect 3617 14501 3651 14535
rect 5549 14501 5583 14535
rect 9965 14501 9999 14535
rect 12173 14501 12207 14535
rect 14565 14501 14599 14535
rect 16037 14501 16071 14535
rect 16957 14501 16991 14535
rect 17877 14501 17911 14535
rect 18061 14501 18095 14535
rect 1501 14433 1535 14467
rect 2605 14433 2639 14467
rect 3065 14433 3099 14467
rect 3341 14433 3375 14467
rect 3893 14433 3927 14467
rect 4169 14433 4203 14467
rect 5733 14433 5767 14467
rect 7941 14433 7975 14467
rect 10149 14433 10183 14467
rect 12357 14433 12391 14467
rect 14749 14433 14783 14467
rect 15209 14433 15243 14467
rect 15577 14433 15611 14467
rect 17233 14433 17267 14467
rect 17693 14433 17727 14467
rect 18429 14433 18463 14467
rect 15945 14365 15979 14399
rect 16221 14365 16255 14399
rect 1685 14297 1719 14331
rect 2053 14297 2087 14331
rect 2881 14297 2915 14331
rect 15117 14297 15151 14331
rect 16773 14297 16807 14331
rect 17509 14297 17543 14331
rect 18245 14297 18279 14331
rect 2329 14229 2363 14263
rect 3433 14229 3467 14263
rect 7757 14229 7791 14263
rect 15393 14229 15427 14263
rect 15669 14229 15703 14263
rect 17417 14229 17451 14263
rect 1961 14025 1995 14059
rect 3341 14025 3375 14059
rect 3525 14025 3559 14059
rect 12817 14025 12851 14059
rect 13185 14025 13219 14059
rect 15025 14025 15059 14059
rect 15209 14025 15243 14059
rect 15393 14025 15427 14059
rect 15577 14025 15611 14059
rect 2789 13957 2823 13991
rect 17049 13957 17083 13991
rect 2605 13889 2639 13923
rect 3065 13889 3099 13923
rect 15761 13889 15795 13923
rect 16313 13889 16347 13923
rect 17141 13889 17175 13923
rect 1501 13821 1535 13855
rect 2145 13821 2179 13855
rect 2421 13821 2455 13855
rect 3157 13821 3191 13855
rect 12725 13821 12759 13855
rect 17509 13821 17543 13855
rect 17693 13821 17727 13855
rect 17877 13821 17911 13855
rect 18061 13821 18095 13855
rect 18429 13821 18463 13855
rect 1869 13753 1903 13787
rect 15853 13753 15887 13787
rect 17325 13753 17359 13787
rect 1593 13685 1627 13719
rect 2329 13685 2363 13719
rect 18337 13685 18371 13719
rect 2513 13481 2547 13515
rect 8493 13481 8527 13515
rect 9505 13481 9539 13515
rect 15301 13481 15335 13515
rect 15761 13481 15795 13515
rect 15991 13481 16025 13515
rect 16313 13481 16347 13515
rect 16589 13481 16623 13515
rect 1869 13413 1903 13447
rect 2329 13413 2363 13447
rect 2973 13413 3007 13447
rect 17049 13413 17083 13447
rect 18981 13413 19015 13447
rect 1501 13345 1535 13379
rect 2053 13345 2087 13379
rect 4721 13345 4755 13379
rect 4813 13345 4847 13379
rect 7030 13345 7064 13379
rect 8401 13345 8435 13379
rect 9873 13345 9907 13379
rect 14749 13345 14783 13379
rect 16094 13345 16128 13379
rect 16497 13345 16531 13379
rect 16957 13345 16991 13379
rect 17693 13345 17727 13379
rect 18061 13345 18095 13379
rect 18429 13345 18463 13379
rect 2145 13277 2179 13311
rect 2789 13277 2823 13311
rect 4905 13277 4939 13311
rect 7297 13277 7331 13311
rect 8677 13277 8711 13311
rect 9965 13277 9999 13311
rect 10057 13277 10091 13311
rect 14473 13277 14507 13311
rect 14657 13277 14691 13311
rect 17141 13277 17175 13311
rect 17417 13277 17451 13311
rect 18245 13277 18279 13311
rect 4261 13209 4295 13243
rect 15117 13209 15151 13243
rect 15393 13209 15427 13243
rect 17877 13209 17911 13243
rect 1593 13141 1627 13175
rect 3433 13141 3467 13175
rect 4353 13141 4387 13175
rect 5273 13141 5307 13175
rect 5917 13141 5951 13175
rect 8033 13141 8067 13175
rect 9229 13141 9263 13175
rect 11529 13141 11563 13175
rect 15669 13141 15703 13175
rect 17417 13141 17451 13175
rect 17601 13141 17635 13175
rect 1961 12937 1995 12971
rect 4813 12937 4847 12971
rect 6653 12937 6687 12971
rect 8493 12937 8527 12971
rect 11897 12937 11931 12971
rect 14657 12937 14691 12971
rect 15577 12937 15611 12971
rect 15853 12937 15887 12971
rect 18337 12937 18371 12971
rect 1685 12869 1719 12903
rect 8125 12869 8159 12903
rect 2145 12801 2179 12835
rect 4629 12801 4663 12835
rect 5457 12801 5491 12835
rect 8033 12801 8067 12835
rect 10793 12801 10827 12835
rect 13829 12801 13863 12835
rect 14105 12801 14139 12835
rect 15393 12801 15427 12835
rect 15577 12801 15611 12835
rect 16405 12801 16439 12835
rect 16773 12801 16807 12835
rect 17141 12801 17175 12835
rect 17785 12801 17819 12835
rect 2513 12733 2547 12767
rect 2973 12733 3007 12767
rect 7766 12733 7800 12767
rect 8401 12733 8435 12767
rect 9873 12733 9907 12767
rect 11713 12733 11747 12767
rect 13205 12733 13239 12767
rect 13461 12733 13495 12767
rect 16221 12733 16255 12767
rect 17601 12733 17635 12767
rect 18153 12733 18187 12767
rect 18521 12733 18555 12767
rect 1501 12665 1535 12699
rect 1869 12665 1903 12699
rect 2697 12665 2731 12699
rect 3240 12665 3274 12699
rect 5181 12665 5215 12699
rect 5641 12665 5675 12699
rect 6193 12665 6227 12699
rect 9606 12665 9640 12699
rect 11069 12665 11103 12699
rect 13645 12665 13679 12699
rect 14197 12665 14231 12699
rect 15117 12665 15151 12699
rect 16313 12665 16347 12699
rect 17693 12665 17727 12699
rect 2329 12597 2363 12631
rect 4353 12597 4387 12631
rect 5273 12597 5307 12631
rect 5917 12597 5951 12631
rect 6561 12597 6595 12631
rect 8401 12597 8435 12631
rect 10517 12597 10551 12631
rect 10977 12597 11011 12631
rect 11437 12597 11471 12631
rect 12081 12597 12115 12631
rect 14289 12597 14323 12631
rect 14749 12597 14783 12631
rect 15209 12597 15243 12631
rect 15669 12597 15703 12631
rect 17233 12597 17267 12631
rect 18981 12461 19015 12495
rect 3525 12393 3559 12427
rect 5089 12393 5123 12427
rect 5181 12393 5215 12427
rect 6009 12393 6043 12427
rect 6561 12393 6595 12427
rect 7665 12393 7699 12427
rect 8217 12393 8251 12427
rect 8585 12393 8619 12427
rect 9597 12393 9631 12427
rect 11897 12393 11931 12427
rect 12357 12393 12391 12427
rect 12817 12393 12851 12427
rect 18153 12393 18187 12427
rect 5641 12325 5675 12359
rect 7757 12325 7791 12359
rect 10692 12325 10726 12359
rect 13952 12325 13986 12359
rect 15976 12325 16010 12359
rect 1501 12257 1535 12291
rect 1869 12257 1903 12291
rect 2412 12257 2446 12291
rect 4261 12257 4295 12291
rect 6469 12257 6503 12291
rect 7021 12257 7055 12291
rect 9965 12257 9999 12291
rect 12265 12257 12299 12291
rect 16405 12257 16439 12291
rect 17621 12257 17655 12291
rect 18429 12257 18463 12291
rect 18981 12257 19015 12291
rect 2145 12189 2179 12223
rect 3617 12189 3651 12223
rect 4353 12189 4387 12223
rect 4537 12189 4571 12223
rect 5273 12189 5307 12223
rect 6653 12189 6687 12223
rect 7573 12189 7607 12223
rect 8677 12189 8711 12223
rect 8861 12189 8895 12223
rect 9321 12189 9355 12223
rect 10057 12189 10091 12223
rect 10241 12189 10275 12223
rect 10425 12189 10459 12223
rect 12449 12189 12483 12223
rect 14197 12189 14231 12223
rect 14749 12189 14783 12223
rect 16221 12189 16255 12223
rect 17877 12189 17911 12223
rect 4721 12121 4755 12155
rect 8125 12121 8159 12155
rect 9413 12121 9447 12155
rect 11805 12121 11839 12155
rect 14841 12121 14875 12155
rect 16497 12121 16531 12155
rect 1593 12053 1627 12087
rect 1961 12053 1995 12087
rect 3893 12053 3927 12087
rect 5825 12053 5859 12087
rect 6101 12053 6135 12087
rect 7205 12053 7239 12087
rect 14381 12053 14415 12087
rect 18337 12053 18371 12087
rect 3525 11849 3559 11883
rect 4721 11849 4755 11883
rect 5549 11849 5583 11883
rect 8861 11849 8895 11883
rect 8953 11849 8987 11883
rect 9873 11849 9907 11883
rect 10701 11849 10735 11883
rect 11529 11849 11563 11883
rect 11989 11849 12023 11883
rect 13461 11849 13495 11883
rect 14381 11849 14415 11883
rect 15945 11849 15979 11883
rect 16773 11849 16807 11883
rect 2237 11713 2271 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 5365 11713 5399 11747
rect 6101 11713 6135 11747
rect 7021 11713 7055 11747
rect 9505 11713 9539 11747
rect 10517 11713 10551 11747
rect 11253 11713 11287 11747
rect 13921 11781 13955 11815
rect 13001 11713 13035 11747
rect 14841 11713 14875 11747
rect 15025 11713 15059 11747
rect 15301 11713 15335 11747
rect 16221 11713 16255 11747
rect 17601 11713 17635 11747
rect 18337 11713 18371 11747
rect 3801 11645 3835 11679
rect 5917 11645 5951 11679
rect 6837 11645 6871 11679
rect 7481 11645 7515 11679
rect 7748 11645 7782 11679
rect 9321 11645 9355 11679
rect 10241 11645 10275 11679
rect 11069 11645 11103 11679
rect 11529 11645 11563 11679
rect 12265 11645 12299 11679
rect 14749 11645 14783 11679
rect 15577 11645 15611 11679
rect 18245 11645 18279 11679
rect 1777 11577 1811 11611
rect 2053 11577 2087 11611
rect 3065 11577 3099 11611
rect 4261 11577 4295 11611
rect 15485 11577 15519 11611
rect 1685 11509 1719 11543
rect 2329 11509 2363 11543
rect 2605 11509 2639 11543
rect 2881 11509 2915 11543
rect 3341 11509 3375 11543
rect 4629 11509 4663 11543
rect 5089 11509 5123 11543
rect 5181 11509 5215 11543
rect 6009 11509 6043 11543
rect 6469 11509 6503 11543
rect 6929 11509 6963 11543
rect 7389 11509 7423 11543
rect 9413 11509 9447 11543
rect 10333 11509 10367 11543
rect 11161 11509 11195 11543
rect 11713 11509 11747 11543
rect 12173 11509 12207 11543
rect 12449 11509 12483 11543
rect 12817 11509 12851 11543
rect 12909 11509 12943 11543
rect 13277 11509 13311 11543
rect 13645 11509 13679 11543
rect 14013 11509 14047 11543
rect 14289 11509 14323 11543
rect 16313 11509 16347 11543
rect 16405 11509 16439 11543
rect 16957 11509 16991 11543
rect 17325 11509 17359 11543
rect 17417 11509 17451 11543
rect 17785 11509 17819 11543
rect 18153 11509 18187 11543
rect 6009 11305 6043 11339
rect 7573 11305 7607 11339
rect 10885 11305 10919 11339
rect 11529 11305 11563 11339
rect 13461 11305 13495 11339
rect 13921 11305 13955 11339
rect 15117 11305 15151 11339
rect 16773 11305 16807 11339
rect 17601 11305 17635 11339
rect 4160 11237 4194 11271
rect 5457 11237 5491 11271
rect 9382 11237 9416 11271
rect 10701 11237 10735 11271
rect 15301 11237 15335 11271
rect 17049 11237 17083 11271
rect 18981 11237 19015 11271
rect 1869 11169 1903 11203
rect 3442 11169 3476 11203
rect 6377 11169 6411 11203
rect 7205 11169 7239 11203
rect 8033 11169 8067 11203
rect 8493 11169 8527 11203
rect 11069 11169 11103 11203
rect 11437 11169 11471 11203
rect 12245 11169 12279 11203
rect 13829 11169 13863 11203
rect 14933 11169 14967 11203
rect 15649 11169 15683 11203
rect 17233 11169 17267 11203
rect 17417 11169 17451 11203
rect 17969 11169 18003 11203
rect 1685 11101 1719 11135
rect 1777 11101 1811 11135
rect 3709 11101 3743 11135
rect 3893 11101 3927 11135
rect 5917 11101 5951 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 7021 11101 7055 11135
rect 7113 11101 7147 11135
rect 7757 11101 7791 11135
rect 7941 11101 7975 11135
rect 9137 11101 9171 11135
rect 11345 11101 11379 11135
rect 11989 11101 12023 11135
rect 14013 11101 14047 11135
rect 14381 11101 14415 11135
rect 15393 11101 15427 11135
rect 18061 11101 18095 11135
rect 18245 11101 18279 11135
rect 2237 11033 2271 11067
rect 8677 11033 8711 11067
rect 10517 11033 10551 11067
rect 16865 11033 16899 11067
rect 18521 11033 18555 11067
rect 2329 10965 2363 10999
rect 5273 10965 5307 10999
rect 5641 10965 5675 10999
rect 8401 10965 8435 10999
rect 8861 10965 8895 10999
rect 11897 10965 11931 10999
rect 13369 10965 13403 10999
rect 14749 10965 14783 10999
rect 2237 10761 2271 10795
rect 2329 10761 2363 10795
rect 7849 10761 7883 10795
rect 10793 10761 10827 10795
rect 18337 10761 18371 10795
rect 4169 10693 4203 10727
rect 9321 10693 9355 10727
rect 10885 10693 10919 10727
rect 11713 10693 11747 10727
rect 14841 10693 14875 10727
rect 1685 10625 1719 10659
rect 2973 10625 3007 10659
rect 3985 10625 4019 10659
rect 16221 10625 16255 10659
rect 16405 10625 16439 10659
rect 16957 10625 16991 10659
rect 1869 10557 1903 10591
rect 2697 10557 2731 10591
rect 3709 10557 3743 10591
rect 5549 10557 5583 10591
rect 6469 10557 6503 10591
rect 7941 10557 7975 10591
rect 8197 10557 8231 10591
rect 9413 10557 9447 10591
rect 11437 10557 11471 10591
rect 13093 10557 13127 10591
rect 13369 10557 13403 10591
rect 16681 10557 16715 10591
rect 5282 10489 5316 10523
rect 5825 10489 5859 10523
rect 6101 10489 6135 10523
rect 6736 10489 6770 10523
rect 9658 10489 9692 10523
rect 11161 10489 11195 10523
rect 11253 10489 11287 10523
rect 12826 10489 12860 10523
rect 13614 10489 13648 10523
rect 15965 10489 15999 10523
rect 16497 10489 16531 10523
rect 17224 10489 17258 10523
rect 1777 10421 1811 10455
rect 2789 10421 2823 10455
rect 3157 10421 3191 10455
rect 3341 10421 3375 10455
rect 3801 10421 3835 10455
rect 5733 10421 5767 10455
rect 6193 10421 6227 10455
rect 13277 10421 13311 10455
rect 14749 10421 14783 10455
rect 18521 10421 18555 10455
rect 3341 10217 3375 10251
rect 4445 10217 4479 10251
rect 4905 10217 4939 10251
rect 6193 10217 6227 10251
rect 6469 10217 6503 10251
rect 7021 10217 7055 10251
rect 7389 10217 7423 10251
rect 7665 10217 7699 10251
rect 9505 10217 9539 10251
rect 9597 10217 9631 10251
rect 10517 10217 10551 10251
rect 10977 10217 11011 10251
rect 11805 10217 11839 10251
rect 13185 10217 13219 10251
rect 13553 10217 13587 10251
rect 14933 10217 14967 10251
rect 15301 10217 15335 10251
rect 15669 10217 15703 10251
rect 16129 10217 16163 10251
rect 16497 10217 16531 10251
rect 17417 10217 17451 10251
rect 17877 10217 17911 10251
rect 4813 10149 4847 10183
rect 8033 10149 8067 10183
rect 8861 10149 8895 10183
rect 10425 10149 10459 10183
rect 14841 10149 14875 10183
rect 1676 10081 1710 10115
rect 4077 10081 4111 10115
rect 4353 10081 4387 10115
rect 5641 10081 5675 10115
rect 8125 10081 8159 10115
rect 11345 10081 11379 10115
rect 12173 10081 12207 10115
rect 12909 10081 12943 10115
rect 13645 10081 13679 10115
rect 14197 10081 14231 10115
rect 17325 10081 17359 10115
rect 17785 10081 17819 10115
rect 18521 10081 18555 10115
rect 1409 10013 1443 10047
rect 3433 10013 3467 10047
rect 3525 10013 3559 10047
rect 5089 10013 5123 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 6745 10013 6779 10047
rect 6929 10013 6963 10047
rect 8309 10013 8343 10047
rect 8677 10013 8711 10047
rect 9689 10013 9723 10047
rect 10333 10013 10367 10047
rect 11437 10013 11471 10047
rect 11621 10013 11655 10047
rect 12265 10013 12299 10047
rect 12449 10013 12483 10047
rect 12817 10013 12851 10047
rect 13737 10013 13771 10047
rect 15025 10013 15059 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16589 10013 16623 10047
rect 16773 10013 16807 10047
rect 18061 10013 18095 10047
rect 4169 9945 4203 9979
rect 5273 9945 5307 9979
rect 10057 9945 10091 9979
rect 10885 9945 10919 9979
rect 2789 9877 2823 9911
rect 2973 9877 3007 9911
rect 3893 9877 3927 9911
rect 6377 9877 6411 9911
rect 7573 9877 7607 9911
rect 9137 9877 9171 9911
rect 13093 9877 13127 9911
rect 14473 9877 14507 9911
rect 17141 9877 17175 9911
rect 18337 9877 18371 9911
rect 3801 9673 3835 9707
rect 13737 9673 13771 9707
rect 16037 9673 16071 9707
rect 1685 9605 1719 9639
rect 2881 9605 2915 9639
rect 5273 9605 5307 9639
rect 5365 9605 5399 9639
rect 6469 9605 6503 9639
rect 6837 9605 6871 9639
rect 7665 9605 7699 9639
rect 8493 9605 8527 9639
rect 11253 9605 11287 9639
rect 11529 9605 11563 9639
rect 15761 9605 15795 9639
rect 2053 9537 2087 9571
rect 2145 9537 2179 9571
rect 4353 9537 4387 9571
rect 4721 9537 4755 9571
rect 6009 9537 6043 9571
rect 7297 9537 7331 9571
rect 7481 9537 7515 9571
rect 8217 9537 8251 9571
rect 9045 9537 9079 9571
rect 9413 9537 9447 9571
rect 10977 9537 11011 9571
rect 12357 9537 12391 9571
rect 16681 9537 16715 9571
rect 2237 9469 2271 9503
rect 3065 9469 3099 9503
rect 3985 9469 4019 9503
rect 4261 9469 4295 9503
rect 5825 9469 5859 9503
rect 6653 9469 6687 9503
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 10710 9469 10744 9503
rect 11897 9469 11931 9503
rect 14197 9469 14231 9503
rect 14464 9469 14498 9503
rect 16957 9469 16991 9503
rect 1501 9401 1535 9435
rect 3341 9401 3375 9435
rect 7205 9401 7239 9435
rect 8033 9401 8067 9435
rect 12624 9401 12658 9435
rect 13829 9401 13863 9435
rect 15853 9401 15887 9435
rect 17224 9401 17258 9435
rect 2605 9333 2639 9367
rect 3617 9333 3651 9367
rect 4077 9333 4111 9367
rect 4813 9333 4847 9367
rect 4905 9333 4939 9367
rect 5733 9333 5767 9367
rect 6193 9333 6227 9367
rect 8125 9333 8159 9367
rect 9597 9333 9631 9367
rect 11161 9333 11195 9367
rect 11713 9333 11747 9367
rect 12081 9333 12115 9367
rect 12265 9333 12299 9367
rect 14013 9333 14047 9367
rect 15577 9333 15611 9367
rect 16405 9333 16439 9367
rect 16497 9333 16531 9367
rect 18337 9333 18371 9367
rect 18521 9333 18555 9367
rect 3617 9129 3651 9163
rect 6377 9129 6411 9163
rect 8217 9129 8251 9163
rect 8861 9129 8895 9163
rect 9137 9129 9171 9163
rect 9965 9129 9999 9163
rect 10885 9129 10919 9163
rect 11345 9129 11379 9163
rect 11713 9129 11747 9163
rect 12173 9129 12207 9163
rect 12541 9129 12575 9163
rect 13001 9129 13035 9163
rect 13369 9129 13403 9163
rect 15761 9129 15795 9163
rect 17509 9129 17543 9163
rect 17877 9129 17911 9163
rect 18337 9129 18371 9163
rect 2504 9061 2538 9095
rect 4138 9061 4172 9095
rect 6009 9061 6043 9095
rect 12633 9061 12667 9095
rect 16282 9061 16316 9095
rect 1501 8993 1535 9027
rect 2145 8993 2179 9027
rect 2237 8993 2271 9027
rect 3893 8993 3927 9027
rect 5457 8993 5491 9027
rect 6837 8993 6871 9027
rect 7104 8993 7138 9027
rect 10793 8993 10827 9027
rect 14841 8993 14875 9027
rect 15393 8993 15427 9027
rect 16037 8993 16071 9027
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 6469 8925 6503 8959
rect 9413 8925 9447 8959
rect 10057 8925 10091 8959
rect 10241 8925 10275 8959
rect 10977 8925 11011 8959
rect 11805 8925 11839 8959
rect 11989 8925 12023 8959
rect 12817 8925 12851 8959
rect 13461 8925 13495 8959
rect 13553 8925 13587 8959
rect 14933 8925 14967 8959
rect 15025 8925 15059 8959
rect 17969 8925 18003 8959
rect 18061 8925 18095 8959
rect 1777 8857 1811 8891
rect 8677 8857 8711 8891
rect 14013 8857 14047 8891
rect 17417 8857 17451 8891
rect 1961 8789 1995 8823
rect 5273 8789 5307 8823
rect 6745 8789 6779 8823
rect 8309 8789 8343 8823
rect 8493 8789 8527 8823
rect 9597 8789 9631 8823
rect 10425 8789 10459 8823
rect 14105 8789 14139 8823
rect 14473 8789 14507 8823
rect 15669 8789 15703 8823
rect 6285 8585 6319 8619
rect 7849 8585 7883 8619
rect 10977 8585 11011 8619
rect 17049 8585 17083 8619
rect 3249 8517 3283 8551
rect 4261 8517 4295 8551
rect 5181 8517 5215 8551
rect 14289 8517 14323 8551
rect 15117 8517 15151 8551
rect 15945 8517 15979 8551
rect 17325 8517 17359 8551
rect 2789 8449 2823 8483
rect 3709 8449 3743 8483
rect 3801 8449 3835 8483
rect 4813 8449 4847 8483
rect 4905 8449 4939 8483
rect 5733 8449 5767 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13921 8449 13955 8483
rect 14105 8449 14139 8483
rect 14749 8449 14783 8483
rect 14933 8449 14967 8483
rect 15669 8449 15703 8483
rect 16497 8449 16531 8483
rect 2533 8381 2567 8415
rect 3065 8381 3099 8415
rect 3433 8381 3467 8415
rect 5365 8381 5399 8415
rect 6469 8381 6503 8415
rect 9341 8381 9375 8415
rect 9597 8381 9631 8415
rect 12909 8381 12943 8415
rect 13829 8381 13863 8415
rect 15485 8381 15519 8415
rect 16313 8381 16347 8415
rect 17141 8381 17175 8415
rect 17417 8381 17451 8415
rect 17785 8381 17819 8415
rect 18061 8381 18095 8415
rect 18429 8381 18463 8415
rect 2881 8313 2915 8347
rect 4721 8313 4755 8347
rect 5917 8313 5951 8347
rect 6714 8313 6748 8347
rect 8125 8313 8159 8347
rect 9689 8313 9723 8347
rect 12173 8313 12207 8347
rect 16405 8313 16439 8347
rect 17969 8313 18003 8347
rect 1409 8245 1443 8279
rect 3893 8245 3927 8279
rect 4353 8245 4387 8279
rect 5825 8245 5859 8279
rect 8217 8245 8251 8279
rect 11805 8245 11839 8279
rect 12265 8245 12299 8279
rect 13001 8245 13035 8279
rect 13369 8245 13403 8279
rect 13461 8245 13495 8279
rect 14657 8245 14691 8279
rect 15577 8245 15611 8279
rect 17601 8245 17635 8279
rect 2053 8041 2087 8075
rect 2605 8041 2639 8075
rect 2973 8041 3007 8075
rect 3893 8041 3927 8075
rect 4353 8041 4387 8075
rect 6285 8041 6319 8075
rect 6377 8041 6411 8075
rect 6837 8041 6871 8075
rect 8309 8041 8343 8075
rect 8677 8041 8711 8075
rect 9505 8041 9539 8075
rect 10701 8041 10735 8075
rect 12725 8041 12759 8075
rect 13461 8041 13495 8075
rect 17233 8041 17267 8075
rect 17601 8041 17635 8075
rect 3433 7973 3467 8007
rect 3617 7973 3651 8007
rect 10241 7973 10275 8007
rect 11590 7973 11624 8007
rect 16098 7973 16132 8007
rect 17785 7973 17819 8007
rect 18429 7973 18463 8007
rect 1593 7905 1627 7939
rect 2145 7905 2179 7939
rect 4261 7905 4295 7939
rect 5172 7905 5206 7939
rect 6561 7905 6595 7939
rect 7021 7905 7055 7939
rect 7481 7905 7515 7939
rect 8217 7905 8251 7939
rect 8769 7905 8803 7939
rect 10333 7905 10367 7939
rect 13829 7905 13863 7939
rect 15494 7905 15528 7939
rect 15761 7905 15795 7939
rect 15853 7905 15887 7939
rect 17417 7905 17451 7939
rect 1961 7837 1995 7871
rect 3065 7837 3099 7871
rect 3157 7837 3191 7871
rect 4445 7837 4479 7871
rect 4905 7837 4939 7871
rect 6745 7837 6779 7871
rect 7205 7837 7239 7871
rect 7389 7837 7423 7871
rect 8125 7837 8159 7871
rect 7849 7769 7883 7803
rect 9597 7837 9631 7871
rect 9689 7837 9723 7871
rect 10149 7837 10183 7871
rect 10885 7837 10919 7871
rect 11345 7837 11379 7871
rect 13093 7837 13127 7871
rect 13921 7837 13955 7871
rect 14105 7837 14139 7871
rect 14381 7769 14415 7803
rect 17969 7769 18003 7803
rect 1501 7701 1535 7735
rect 2513 7701 2547 7735
rect 4721 7701 4755 7735
rect 8769 7701 8803 7735
rect 8953 7701 8987 7735
rect 9137 7701 9171 7735
rect 11253 7701 11287 7735
rect 13277 7701 13311 7735
rect 18153 7701 18187 7735
rect 1409 7497 1443 7531
rect 2973 7497 3007 7531
rect 3525 7497 3559 7531
rect 4905 7497 4939 7531
rect 6469 7497 6503 7531
rect 12357 7497 12391 7531
rect 13185 7497 13219 7531
rect 14565 7497 14599 7531
rect 15393 7497 15427 7531
rect 16773 7497 16807 7531
rect 17325 7497 17359 7531
rect 17509 7497 17543 7531
rect 3065 7429 3099 7463
rect 8493 7429 8527 7463
rect 12173 7429 12207 7463
rect 14381 7429 14415 7463
rect 16497 7429 16531 7463
rect 4261 7361 4295 7395
rect 7113 7361 7147 7395
rect 7757 7361 7791 7395
rect 7941 7361 7975 7395
rect 10149 7361 10183 7395
rect 11897 7361 11931 7395
rect 13001 7361 13035 7395
rect 13737 7361 13771 7395
rect 15209 7361 15243 7395
rect 15945 7361 15979 7395
rect 17141 7361 17175 7395
rect 18521 7361 18555 7395
rect 1593 7293 1627 7327
rect 1849 7293 1883 7327
rect 4077 7293 4111 7327
rect 6029 7293 6063 7327
rect 6285 7293 6319 7327
rect 8117 7293 8151 7327
rect 8585 7293 8619 7327
rect 8841 7293 8875 7327
rect 12817 7293 12851 7327
rect 13553 7293 13587 7327
rect 14933 7293 14967 7327
rect 17601 7293 17635 7327
rect 17877 7293 17911 7327
rect 3249 7225 3283 7259
rect 7665 7225 7699 7259
rect 10416 7225 10450 7259
rect 12725 7225 12759 7259
rect 14197 7225 14231 7259
rect 15025 7225 15059 7259
rect 16221 7225 16255 7259
rect 18337 7225 18371 7259
rect 3617 7157 3651 7191
rect 3985 7157 4019 7191
rect 4445 7157 4479 7191
rect 4813 7157 4847 7191
rect 6837 7157 6871 7191
rect 6929 7157 6963 7191
rect 7297 7157 7331 7191
rect 8309 7157 8343 7191
rect 9965 7157 9999 7191
rect 11529 7157 11563 7191
rect 11805 7157 11839 7191
rect 13645 7157 13679 7191
rect 14105 7157 14139 7191
rect 15761 7157 15795 7191
rect 15853 7157 15887 7191
rect 17785 7157 17819 7191
rect 18061 7157 18095 7191
rect 2145 6953 2179 6987
rect 4261 6953 4295 6987
rect 6009 6953 6043 6987
rect 8861 6953 8895 6987
rect 9505 6953 9539 6987
rect 15393 6953 15427 6987
rect 17233 6953 17267 6987
rect 17509 6953 17543 6987
rect 17785 6953 17819 6987
rect 1961 6885 1995 6919
rect 2574 6885 2608 6919
rect 4353 6885 4387 6919
rect 5181 6885 5215 6919
rect 6837 6885 6871 6919
rect 7748 6885 7782 6919
rect 11437 6885 11471 6919
rect 11713 6885 11747 6919
rect 12173 6885 12207 6919
rect 14749 6885 14783 6919
rect 17969 6885 18003 6919
rect 1593 6817 1627 6851
rect 1777 6817 1811 6851
rect 2329 6817 2363 6851
rect 5089 6817 5123 6851
rect 6101 6817 6135 6851
rect 7481 6817 7515 6851
rect 11089 6817 11123 6851
rect 13001 6817 13035 6851
rect 13829 6817 13863 6851
rect 15669 6817 15703 6851
rect 18153 6817 18187 6851
rect 18337 6817 18371 6851
rect 4537 6749 4571 6783
rect 5273 6749 5307 6783
rect 6285 6749 6319 6783
rect 6929 6749 6963 6783
rect 7113 6749 7147 6783
rect 7389 6749 7423 6783
rect 9321 6749 9355 6783
rect 9413 6749 9447 6783
rect 11345 6749 11379 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 12725 6749 12759 6783
rect 12909 6749 12943 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 14841 6749 14875 6783
rect 15025 6749 15059 6783
rect 3893 6681 3927 6715
rect 5641 6681 5675 6715
rect 9965 6681 9999 6715
rect 12541 6681 12575 6715
rect 13461 6681 13495 6715
rect 15945 6681 15979 6715
rect 18521 6681 18555 6715
rect 1501 6613 1535 6647
rect 3709 6613 3743 6647
rect 4721 6613 4755 6647
rect 6469 6613 6503 6647
rect 9873 6613 9907 6647
rect 13369 6613 13403 6647
rect 14381 6613 14415 6647
rect 15485 6613 15519 6647
rect 16957 6613 16991 6647
rect 2605 6409 2639 6443
rect 2973 6409 3007 6443
rect 7941 6409 7975 6443
rect 10517 6409 10551 6443
rect 11529 6409 11563 6443
rect 11989 6409 12023 6443
rect 12817 6409 12851 6443
rect 13645 6409 13679 6443
rect 17417 6409 17451 6443
rect 17785 6409 17819 6443
rect 2697 6341 2731 6375
rect 7849 6341 7883 6375
rect 10425 6341 10459 6375
rect 11713 6341 11747 6375
rect 3525 6273 3559 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 8493 6273 8527 6307
rect 10977 6273 11011 6307
rect 12449 6273 12483 6307
rect 12633 6273 12667 6307
rect 13369 6273 13403 6307
rect 1593 6205 1627 6239
rect 2145 6205 2179 6239
rect 2421 6205 2455 6239
rect 2881 6205 2915 6239
rect 3341 6205 3375 6239
rect 3433 6205 3467 6239
rect 3985 6205 4019 6239
rect 5190 6205 5224 6239
rect 5457 6205 5491 6239
rect 5917 6205 5951 6239
rect 6469 6205 6503 6239
rect 8769 6205 8803 6239
rect 9045 6205 9079 6239
rect 10701 6205 10735 6239
rect 11069 6205 11103 6239
rect 11161 6205 11195 6239
rect 11897 6205 11931 6239
rect 13277 6205 13311 6239
rect 14758 6205 14792 6239
rect 15025 6205 15059 6239
rect 15117 6205 15151 6239
rect 17233 6205 17267 6239
rect 17601 6205 17635 6239
rect 17877 6205 17911 6239
rect 1961 6137 1995 6171
rect 6714 6137 6748 6171
rect 9312 6137 9346 6171
rect 13185 6137 13219 6171
rect 15577 6137 15611 6171
rect 18337 6137 18371 6171
rect 18521 6137 18555 6171
rect 1501 6069 1535 6103
rect 1869 6069 1903 6103
rect 2329 6069 2363 6103
rect 3801 6069 3835 6103
rect 4077 6069 4111 6103
rect 6285 6069 6319 6103
rect 8309 6069 8343 6103
rect 8401 6069 8435 6103
rect 8953 6069 8987 6103
rect 12357 6069 12391 6103
rect 15301 6069 15335 6103
rect 15485 6069 15519 6103
rect 18061 6069 18095 6103
rect 3709 5865 3743 5899
rect 4353 5865 4387 5899
rect 4721 5865 4755 5899
rect 5089 5865 5123 5899
rect 5549 5865 5583 5899
rect 7205 5865 7239 5899
rect 9413 5865 9447 5899
rect 11437 5865 11471 5899
rect 13553 5865 13587 5899
rect 14841 5865 14875 5899
rect 15669 5865 15703 5899
rect 16129 5865 16163 5899
rect 17785 5865 17819 5899
rect 1860 5797 1894 5831
rect 6684 5797 6718 5831
rect 8953 5797 8987 5831
rect 12440 5797 12474 5831
rect 17417 5797 17451 5831
rect 18337 5797 18371 5831
rect 1501 5729 1535 5763
rect 3065 5729 3099 5763
rect 3525 5729 3559 5763
rect 4261 5729 4295 5763
rect 5181 5729 5215 5763
rect 6929 5729 6963 5763
rect 7113 5729 7147 5763
rect 8329 5729 8363 5763
rect 9505 5729 9539 5763
rect 9965 5729 9999 5763
rect 10232 5729 10266 5763
rect 11805 5729 11839 5763
rect 12173 5729 12207 5763
rect 14749 5729 14783 5763
rect 15577 5729 15611 5763
rect 17325 5729 17359 5763
rect 17601 5729 17635 5763
rect 17877 5729 17911 5763
rect 1593 5661 1627 5695
rect 4537 5661 4571 5695
rect 5273 5661 5307 5695
rect 8585 5661 8619 5695
rect 9321 5661 9355 5695
rect 13737 5661 13771 5695
rect 15025 5661 15059 5695
rect 15761 5661 15795 5695
rect 3341 5593 3375 5627
rect 11621 5593 11655 5627
rect 11989 5593 12023 5627
rect 18521 5593 18555 5627
rect 2973 5525 3007 5559
rect 3249 5525 3283 5559
rect 3893 5525 3927 5559
rect 9873 5525 9907 5559
rect 11345 5525 11379 5559
rect 13829 5525 13863 5559
rect 14105 5525 14139 5559
rect 14381 5525 14415 5559
rect 15209 5525 15243 5559
rect 18061 5525 18095 5559
rect 6561 5321 6595 5355
rect 8217 5321 8251 5355
rect 8493 5321 8527 5355
rect 9321 5321 9355 5355
rect 10149 5321 10183 5355
rect 5917 5253 5951 5287
rect 14105 5253 14139 5287
rect 17693 5253 17727 5287
rect 2789 5185 2823 5219
rect 3709 5185 3743 5219
rect 4445 5185 4479 5219
rect 4629 5185 4663 5219
rect 5365 5185 5399 5219
rect 6193 5185 6227 5219
rect 7205 5185 7239 5219
rect 8033 5185 8067 5219
rect 8953 5185 8987 5219
rect 9137 5185 9171 5219
rect 9873 5185 9907 5219
rect 10977 5185 11011 5219
rect 13829 5185 13863 5219
rect 15577 5185 15611 5219
rect 15945 5185 15979 5219
rect 18521 5185 18555 5219
rect 3065 5117 3099 5151
rect 3617 5117 3651 5151
rect 4353 5117 4387 5151
rect 6101 5117 6135 5151
rect 6929 5117 6963 5151
rect 8401 5117 8435 5151
rect 9689 5117 9723 5151
rect 10793 5117 10827 5151
rect 12837 5117 12871 5151
rect 13093 5117 13127 5151
rect 13737 5117 13771 5151
rect 15485 5117 15519 5151
rect 17877 5117 17911 5151
rect 18337 5117 18371 5151
rect 2544 5049 2578 5083
rect 3525 5049 3559 5083
rect 5181 5049 5215 5083
rect 5641 5049 5675 5083
rect 9781 5049 9815 5083
rect 11253 5049 11287 5083
rect 11437 5049 11471 5083
rect 13645 5049 13679 5083
rect 15218 5049 15252 5083
rect 1409 4981 1443 5015
rect 2881 4981 2915 5015
rect 3157 4981 3191 5015
rect 3985 4981 4019 5015
rect 4813 4981 4847 5015
rect 5273 4981 5307 5015
rect 7021 4981 7055 5015
rect 7389 4981 7423 5015
rect 7757 4981 7791 5015
rect 7849 4981 7883 5015
rect 8861 4981 8895 5015
rect 10425 4981 10459 5015
rect 10885 4981 10919 5015
rect 11713 4981 11747 5015
rect 13277 4981 13311 5015
rect 18061 4981 18095 5015
rect 1869 4777 1903 4811
rect 2513 4777 2547 4811
rect 2973 4777 3007 4811
rect 3433 4777 3467 4811
rect 7113 4777 7147 4811
rect 7481 4777 7515 4811
rect 9229 4777 9263 4811
rect 9781 4777 9815 4811
rect 12173 4777 12207 4811
rect 12633 4777 12667 4811
rect 12725 4777 12759 4811
rect 13093 4777 13127 4811
rect 13461 4777 13495 4811
rect 14381 4777 14415 4811
rect 14841 4777 14875 4811
rect 15301 4777 15335 4811
rect 1409 4709 1443 4743
rect 1593 4709 1627 4743
rect 2421 4709 2455 4743
rect 3341 4709 3375 4743
rect 7849 4709 7883 4743
rect 10916 4709 10950 4743
rect 14105 4709 14139 4743
rect 14749 4709 14783 4743
rect 17417 4709 17451 4743
rect 17969 4709 18003 4743
rect 18337 4709 18371 4743
rect 1961 4641 1995 4675
rect 3893 4641 3927 4675
rect 4160 4641 4194 4675
rect 5733 4641 5767 4675
rect 6193 4641 6227 4675
rect 7021 4641 7055 4675
rect 8585 4641 8619 4675
rect 9321 4641 9355 4675
rect 11621 4641 11655 4675
rect 13553 4641 13587 4675
rect 18153 4641 18187 4675
rect 2237 4573 2271 4607
rect 3525 4573 3559 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 6469 4573 6503 4607
rect 7297 4573 7331 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 9597 4573 9631 4607
rect 11161 4573 11195 4607
rect 11713 4573 11747 4607
rect 11805 4573 11839 4607
rect 12817 4573 12851 4607
rect 13737 4573 13771 4607
rect 14013 4573 14047 4607
rect 15025 4573 15059 4607
rect 6377 4505 6411 4539
rect 6653 4505 6687 4539
rect 8677 4505 8711 4539
rect 9505 4505 9539 4539
rect 11253 4505 11287 4539
rect 18521 4505 18555 4539
rect 2881 4437 2915 4471
rect 5273 4437 5307 4471
rect 6101 4437 6135 4471
rect 8309 4437 8343 4471
rect 8861 4437 8895 4471
rect 12265 4437 12299 4471
rect 7665 4233 7699 4267
rect 9137 4233 9171 4267
rect 10977 4233 11011 4267
rect 14473 4233 14507 4267
rect 15485 4233 15519 4267
rect 4905 4165 4939 4199
rect 13553 4165 13587 4199
rect 14381 4165 14415 4199
rect 17509 4165 17543 4199
rect 3525 4097 3559 4131
rect 5273 4097 5307 4131
rect 6009 4097 6043 4131
rect 7021 4097 7055 4131
rect 9689 4097 9723 4131
rect 9781 4097 9815 4131
rect 10517 4097 10551 4131
rect 10609 4097 10643 4131
rect 11713 4097 11747 4131
rect 13829 4097 13863 4131
rect 13921 4097 13955 4131
rect 14933 4097 14967 4131
rect 15117 4097 15151 4131
rect 16681 4097 16715 4131
rect 1777 4029 1811 4063
rect 2053 4029 2087 4063
rect 5089 4029 5123 4063
rect 5549 4029 5583 4063
rect 6837 4029 6871 4063
rect 7297 4029 7331 4063
rect 7757 4029 7791 4063
rect 10425 4029 10459 4063
rect 11069 4029 11103 4063
rect 11980 4029 12014 4063
rect 14013 4029 14047 4063
rect 16589 4029 16623 4063
rect 17049 4029 17083 4063
rect 17325 4029 17359 4063
rect 17601 4029 17635 4063
rect 18337 4029 18371 4063
rect 1593 3961 1627 3995
rect 2298 3961 2332 3995
rect 3770 3961 3804 3995
rect 6929 3961 6963 3995
rect 8024 3961 8058 3995
rect 17969 3961 18003 3995
rect 18153 3961 18187 3995
rect 18521 3961 18555 3995
rect 1501 3893 1535 3927
rect 1961 3893 1995 3927
rect 3433 3893 3467 3927
rect 5457 3893 5491 3927
rect 5917 3893 5951 3927
rect 6469 3893 6503 3927
rect 7481 3893 7515 3927
rect 9229 3893 9263 3927
rect 9597 3893 9631 3927
rect 10057 3893 10091 3927
rect 11345 3893 11379 3927
rect 13093 3893 13127 3927
rect 13277 3893 13311 3927
rect 14841 3893 14875 3927
rect 15393 3893 15427 3927
rect 17233 3893 17267 3927
rect 17785 3893 17819 3927
rect 3341 3689 3375 3723
rect 4721 3689 4755 3723
rect 7481 3689 7515 3723
rect 7941 3689 7975 3723
rect 8861 3689 8895 3723
rect 9137 3689 9171 3723
rect 9597 3689 9631 3723
rect 10885 3689 10919 3723
rect 11253 3689 11287 3723
rect 11989 3689 12023 3723
rect 13461 3689 13495 3723
rect 13921 3689 13955 3723
rect 15761 3689 15795 3723
rect 1593 3621 1627 3655
rect 2329 3621 2363 3655
rect 2881 3621 2915 3655
rect 3065 3621 3099 3655
rect 3433 3621 3467 3655
rect 7297 3621 7331 3655
rect 9505 3621 9539 3655
rect 10149 3621 10183 3655
rect 14626 3621 14660 3655
rect 16405 3621 16439 3655
rect 17969 3621 18003 3655
rect 1961 3553 1995 3587
rect 2697 3553 2731 3587
rect 4261 3553 4295 3587
rect 4905 3553 4939 3587
rect 5181 3553 5215 3587
rect 5529 3553 5563 3587
rect 6929 3553 6963 3587
rect 7205 3553 7239 3587
rect 7849 3553 7883 3587
rect 8309 3553 8343 3587
rect 8585 3553 8619 3587
rect 11713 3553 11747 3587
rect 12337 3553 12371 3587
rect 16221 3553 16255 3587
rect 16957 3553 16991 3587
rect 17233 3553 17267 3587
rect 17601 3553 17635 3587
rect 18337 3553 18371 3587
rect 2513 3485 2547 3519
rect 3709 3485 3743 3519
rect 4077 3485 4111 3519
rect 4169 3485 4203 3519
rect 5273 3485 5307 3519
rect 8033 3485 8067 3519
rect 9689 3485 9723 3519
rect 10609 3485 10643 3519
rect 10793 3485 10827 3519
rect 11437 3485 11471 3519
rect 12081 3485 12115 3519
rect 14381 3485 14415 3519
rect 16681 3485 16715 3519
rect 18521 3485 18555 3519
rect 4997 3417 5031 3451
rect 8769 3417 8803 3451
rect 9965 3417 9999 3451
rect 11529 3417 11563 3451
rect 17785 3417 17819 3451
rect 18153 3417 18187 3451
rect 1501 3349 1535 3383
rect 1869 3349 1903 3383
rect 2237 3349 2271 3383
rect 4629 3349 4663 3383
rect 6653 3349 6687 3383
rect 6745 3349 6779 3383
rect 7021 3349 7055 3383
rect 8493 3349 8527 3383
rect 10425 3349 10459 3383
rect 13645 3349 13679 3383
rect 13737 3349 13771 3383
rect 16865 3349 16899 3383
rect 17141 3349 17175 3383
rect 17417 3349 17451 3383
rect 3893 3145 3927 3179
rect 3985 3145 4019 3179
rect 7941 3145 7975 3179
rect 8953 3145 8987 3179
rect 9781 3145 9815 3179
rect 10057 3145 10091 3179
rect 13553 3145 13587 3179
rect 13737 3145 13771 3179
rect 15577 3145 15611 3179
rect 2881 3077 2915 3111
rect 5641 3077 5675 3111
rect 13185 3077 13219 3111
rect 13921 3077 13955 3111
rect 17785 3077 17819 3111
rect 3341 3009 3375 3043
rect 4629 3009 4663 3043
rect 5273 3009 5307 3043
rect 5365 3009 5399 3043
rect 9229 3009 9263 3043
rect 10609 3009 10643 3043
rect 10793 3009 10827 3043
rect 11805 3009 11839 3043
rect 11989 3009 12023 3043
rect 16037 3009 16071 3043
rect 18521 3009 18555 3043
rect 1593 2941 1627 2975
rect 1961 2941 1995 2975
rect 3065 2941 3099 2975
rect 3525 2941 3559 2975
rect 4353 2941 4387 2975
rect 5181 2941 5215 2975
rect 5825 2941 5859 2975
rect 6101 2941 6135 2975
rect 6561 2941 6595 2975
rect 8217 2941 8251 2975
rect 8493 2941 8527 2975
rect 8769 2941 8803 2975
rect 9413 2941 9447 2975
rect 11529 2941 11563 2975
rect 13093 2941 13127 2975
rect 13369 2941 13403 2975
rect 14105 2941 14139 2975
rect 16313 2941 16347 2975
rect 16773 2941 16807 2975
rect 17141 2941 17175 2975
rect 17233 2941 17267 2975
rect 17601 2941 17635 2975
rect 17969 2941 18003 2975
rect 18337 2941 18371 2975
rect 1409 2873 1443 2907
rect 1777 2873 1811 2907
rect 2329 2873 2363 2907
rect 2697 2873 2731 2907
rect 6806 2873 6840 2907
rect 9321 2873 9355 2907
rect 10977 2873 11011 2907
rect 11161 2873 11195 2907
rect 12541 2873 12575 2907
rect 12725 2873 12759 2907
rect 16497 2873 16531 2907
rect 2237 2805 2271 2839
rect 2605 2805 2639 2839
rect 3433 2805 3467 2839
rect 4445 2805 4479 2839
rect 4813 2805 4847 2839
rect 5917 2805 5951 2839
rect 6193 2805 6227 2839
rect 8033 2805 8067 2839
rect 8309 2805 8343 2839
rect 8585 2805 8619 2839
rect 10149 2805 10183 2839
rect 10517 2805 10551 2839
rect 11345 2805 11379 2839
rect 12081 2805 12115 2839
rect 12449 2805 12483 2839
rect 12909 2805 12943 2839
rect 15761 2805 15795 2839
rect 16129 2805 16163 2839
rect 16957 2805 16991 2839
rect 17417 2805 17451 2839
rect 18061 2805 18095 2839
rect 4261 2601 4295 2635
rect 4721 2601 4755 2635
rect 5181 2601 5215 2635
rect 5917 2601 5951 2635
rect 9597 2601 9631 2635
rect 9873 2601 9907 2635
rect 10241 2601 10275 2635
rect 10333 2601 10367 2635
rect 11069 2601 11103 2635
rect 11437 2601 11471 2635
rect 11713 2601 11747 2635
rect 11897 2601 11931 2635
rect 12357 2601 12391 2635
rect 13461 2601 13495 2635
rect 14565 2601 14599 2635
rect 15209 2601 15243 2635
rect 15669 2601 15703 2635
rect 16221 2601 16255 2635
rect 2145 2533 2179 2567
rect 2329 2533 2363 2567
rect 4169 2533 4203 2567
rect 6745 2533 6779 2567
rect 8217 2533 8251 2567
rect 8401 2533 8435 2567
rect 8585 2533 8619 2567
rect 8953 2533 8987 2567
rect 9413 2533 9447 2567
rect 10977 2533 11011 2567
rect 12265 2533 12299 2567
rect 13277 2533 13311 2567
rect 14105 2533 14139 2567
rect 15025 2533 15059 2567
rect 16405 2533 16439 2567
rect 17601 2533 17635 2567
rect 18337 2533 18371 2567
rect 2053 2465 2087 2499
rect 2697 2465 2731 2499
rect 3249 2465 3283 2499
rect 3525 2465 3559 2499
rect 5089 2465 5123 2499
rect 5825 2465 5859 2499
rect 6929 2465 6963 2499
rect 11529 2465 11563 2499
rect 12909 2465 12943 2499
rect 13645 2465 13679 2499
rect 14749 2465 14783 2499
rect 15393 2465 15427 2499
rect 15485 2465 15519 2499
rect 15761 2465 15795 2499
rect 16037 2465 16071 2499
rect 16865 2465 16899 2499
rect 17233 2465 17267 2499
rect 17969 2465 18003 2499
rect 1869 2397 1903 2431
rect 4077 2397 4111 2431
rect 5273 2397 5307 2431
rect 5733 2397 5767 2431
rect 7757 2397 7791 2431
rect 9229 2397 9263 2431
rect 10517 2397 10551 2431
rect 10885 2397 10919 2431
rect 12449 2397 12483 2431
rect 1501 2329 1535 2363
rect 2513 2329 2547 2363
rect 3065 2329 3099 2363
rect 3709 2329 3743 2363
rect 4629 2329 4663 2363
rect 6561 2329 6595 2363
rect 8769 2329 8803 2363
rect 12725 2329 12759 2363
rect 13093 2329 13127 2363
rect 13921 2329 13955 2363
rect 14841 2329 14875 2363
rect 15945 2329 15979 2363
rect 16589 2329 16623 2363
rect 17417 2329 17451 2363
rect 18521 2329 18555 2363
rect 2973 2261 3007 2295
rect 6285 2261 6319 2295
rect 8125 2261 8159 2295
rect 16773 2261 16807 2295
rect 17693 2261 17727 2295
rect 18061 2261 18095 2295
<< metal1 >>
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 17770 14940 17776 14952
rect 15344 14912 17776 14940
rect 15344 14900 15350 14912
rect 17770 14900 17776 14912
rect 17828 14900 17834 14952
rect 2314 14832 2320 14884
rect 2372 14872 2378 14884
rect 12710 14872 12716 14884
rect 2372 14844 12716 14872
rect 2372 14832 2378 14844
rect 12710 14832 12716 14844
rect 12768 14832 12774 14884
rect 15470 14832 15476 14884
rect 15528 14872 15534 14884
rect 16390 14872 16396 14884
rect 15528 14844 16396 14872
rect 15528 14832 15534 14844
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 17218 14804 17224 14816
rect 4120 14776 17224 14804
rect 4120 14764 4126 14776
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 2590 14560 2596 14612
rect 2648 14600 2654 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2648 14572 2697 14600
rect 2648 14560 2654 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 4062 14600 4068 14612
rect 4023 14572 4068 14600
rect 2685 14563 2743 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7800 14572 8033 14600
rect 7800 14560 7806 14572
rect 1854 14532 1860 14544
rect 1815 14504 1860 14532
rect 1854 14492 1860 14504
rect 1912 14492 1918 14544
rect 2222 14532 2228 14544
rect 2183 14504 2228 14532
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 3602 14532 3608 14544
rect 3563 14504 3608 14532
rect 3602 14492 3608 14504
rect 3660 14492 3666 14544
rect 5534 14532 5540 14544
rect 5495 14504 5540 14532
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 1872 14396 1900 14492
rect 2498 14424 2504 14476
rect 2556 14464 2562 14476
rect 2593 14467 2651 14473
rect 2593 14464 2605 14467
rect 2556 14436 2605 14464
rect 2556 14424 2562 14436
rect 2593 14433 2605 14436
rect 2639 14464 2651 14467
rect 2866 14464 2872 14476
rect 2639 14436 2872 14464
rect 2639 14433 2651 14436
rect 2593 14427 2651 14433
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 2958 14424 2964 14476
rect 3016 14464 3022 14476
rect 3053 14467 3111 14473
rect 3053 14464 3065 14467
rect 3016 14436 3065 14464
rect 3016 14424 3022 14436
rect 3053 14433 3065 14436
rect 3099 14464 3111 14467
rect 3329 14467 3387 14473
rect 3099 14436 3280 14464
rect 3099 14433 3111 14436
rect 3053 14427 3111 14433
rect 3252 14408 3280 14436
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 2682 14396 2688 14408
rect 1872 14368 2688 14396
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 3344 14396 3372 14427
rect 3418 14424 3424 14476
rect 3476 14464 3482 14476
rect 7944 14473 7972 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 16574 14600 16580 14612
rect 8021 14563 8079 14569
rect 15212 14572 16580 14600
rect 9950 14532 9956 14544
rect 9911 14504 9956 14532
rect 9950 14492 9956 14504
rect 10008 14492 10014 14544
rect 12158 14532 12164 14544
rect 12119 14504 12164 14532
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 14553 14535 14611 14541
rect 14553 14532 14565 14535
rect 14424 14504 14565 14532
rect 14424 14492 14430 14504
rect 14553 14501 14565 14504
rect 14599 14501 14611 14535
rect 14553 14495 14611 14501
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3476 14436 3893 14464
rect 3476 14424 3482 14436
rect 3881 14433 3893 14436
rect 3927 14464 3939 14467
rect 4157 14467 4215 14473
rect 4157 14464 4169 14467
rect 3927 14436 4169 14464
rect 3927 14433 3939 14436
rect 3881 14427 3939 14433
rect 4157 14433 4169 14436
rect 4203 14433 4215 14467
rect 4157 14427 4215 14433
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14433 5779 14467
rect 5721 14427 5779 14433
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14433 7987 14467
rect 7929 14427 7987 14433
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 11514 14464 11520 14476
rect 10183 14436 11520 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 3510 14396 3516 14408
rect 3344 14368 3516 14396
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 5736 14396 5764 14427
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 12342 14464 12348 14476
rect 12303 14436 12348 14464
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 14734 14464 14740 14476
rect 14695 14436 14740 14464
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 15212 14473 15240 14572
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 16025 14535 16083 14541
rect 16025 14532 16037 14535
rect 15304 14504 16037 14532
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 15068 14436 15209 14464
rect 15068 14424 15074 14436
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 14752 14396 14780 14424
rect 15304 14396 15332 14504
rect 16025 14501 16037 14504
rect 16071 14532 16083 14535
rect 16206 14532 16212 14544
rect 16071 14504 16212 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 16390 14492 16396 14544
rect 16448 14532 16454 14544
rect 16945 14535 17003 14541
rect 16945 14532 16957 14535
rect 16448 14504 16957 14532
rect 16448 14492 16454 14504
rect 16945 14501 16957 14504
rect 16991 14501 17003 14535
rect 16945 14495 17003 14501
rect 17402 14492 17408 14544
rect 17460 14532 17466 14544
rect 17865 14535 17923 14541
rect 17865 14532 17877 14535
rect 17460 14504 17877 14532
rect 17460 14492 17466 14504
rect 17865 14501 17877 14504
rect 17911 14501 17923 14535
rect 18046 14532 18052 14544
rect 18007 14504 18052 14532
rect 17865 14495 17923 14501
rect 18046 14492 18052 14504
rect 18104 14492 18110 14544
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14433 15623 14467
rect 17218 14464 17224 14476
rect 17179 14436 17224 14464
rect 15565 14427 15623 14433
rect 5736 14368 12434 14396
rect 14752 14368 15332 14396
rect 1670 14328 1676 14340
rect 1631 14300 1676 14328
rect 1670 14288 1676 14300
rect 1728 14288 1734 14340
rect 2041 14331 2099 14337
rect 2041 14297 2053 14331
rect 2087 14328 2099 14331
rect 2498 14328 2504 14340
rect 2087 14300 2504 14328
rect 2087 14297 2099 14300
rect 2041 14291 2099 14297
rect 2498 14288 2504 14300
rect 2556 14288 2562 14340
rect 2869 14331 2927 14337
rect 2869 14297 2881 14331
rect 2915 14328 2927 14331
rect 3602 14328 3608 14340
rect 2915 14300 3608 14328
rect 2915 14297 2927 14300
rect 2869 14291 2927 14297
rect 3602 14288 3608 14300
rect 3660 14288 3666 14340
rect 8202 14328 8208 14340
rect 7576 14300 8208 14328
rect 2317 14263 2375 14269
rect 2317 14229 2329 14263
rect 2363 14260 2375 14263
rect 3326 14260 3332 14272
rect 2363 14232 3332 14260
rect 2363 14229 2375 14232
rect 2317 14223 2375 14229
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14260 3479 14263
rect 7576 14260 7604 14300
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 7742 14260 7748 14272
rect 3467 14232 7604 14260
rect 7703 14232 7748 14260
rect 3467 14229 3479 14232
rect 3421 14223 3479 14229
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 12406 14260 12434 14368
rect 15105 14331 15163 14337
rect 15105 14297 15117 14331
rect 15151 14328 15163 14331
rect 15194 14328 15200 14340
rect 15151 14300 15200 14328
rect 15151 14297 15163 14300
rect 15105 14291 15163 14297
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15580 14328 15608 14427
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 17678 14464 17684 14476
rect 17639 14436 17684 14464
rect 17678 14424 17684 14436
rect 17736 14424 17742 14476
rect 18414 14464 18420 14476
rect 18375 14436 18420 14464
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16114 14396 16120 14408
rect 15979 14368 16120 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14365 16267 14399
rect 18782 14396 18788 14408
rect 16209 14359 16267 14365
rect 17052 14368 18788 14396
rect 16224 14328 16252 14359
rect 15580 14300 16252 14328
rect 16666 14288 16672 14340
rect 16724 14328 16730 14340
rect 16761 14331 16819 14337
rect 16761 14328 16773 14331
rect 16724 14300 16773 14328
rect 16724 14288 16730 14300
rect 16761 14297 16773 14300
rect 16807 14297 16819 14331
rect 16761 14291 16819 14297
rect 14918 14260 14924 14272
rect 12406 14232 14924 14260
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 15378 14260 15384 14272
rect 15339 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 15657 14263 15715 14269
rect 15657 14229 15669 14263
rect 15703 14260 15715 14263
rect 17052 14260 17080 14368
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 17218 14288 17224 14340
rect 17276 14328 17282 14340
rect 17497 14331 17555 14337
rect 17497 14328 17509 14331
rect 17276 14300 17509 14328
rect 17276 14288 17282 14300
rect 17497 14297 17509 14300
rect 17543 14297 17555 14331
rect 17497 14291 17555 14297
rect 18046 14288 18052 14340
rect 18104 14328 18110 14340
rect 18233 14331 18291 14337
rect 18233 14328 18245 14331
rect 18104 14300 18245 14328
rect 18104 14288 18110 14300
rect 18233 14297 18245 14300
rect 18279 14297 18291 14331
rect 18233 14291 18291 14297
rect 15703 14232 17080 14260
rect 17405 14263 17463 14269
rect 15703 14229 15715 14232
rect 15657 14223 15715 14229
rect 17405 14229 17417 14263
rect 17451 14260 17463 14263
rect 18138 14260 18144 14272
rect 17451 14232 18144 14260
rect 17451 14229 17463 14232
rect 17405 14223 17463 14229
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 1486 14016 1492 14068
rect 1544 14016 1550 14068
rect 1949 14059 2007 14065
rect 1949 14025 1961 14059
rect 1995 14056 2007 14059
rect 1995 14028 3096 14056
rect 1995 14025 2007 14028
rect 1949 14019 2007 14025
rect 1504 13988 1532 14016
rect 2777 13991 2835 13997
rect 2777 13988 2789 13991
rect 1504 13960 2789 13988
rect 2777 13957 2789 13960
rect 2823 13957 2835 13991
rect 3068 13988 3096 14028
rect 3234 14016 3240 14068
rect 3292 14056 3298 14068
rect 3329 14059 3387 14065
rect 3329 14056 3341 14059
rect 3292 14028 3341 14056
rect 3292 14016 3298 14028
rect 3329 14025 3341 14028
rect 3375 14025 3387 14059
rect 3510 14056 3516 14068
rect 3471 14028 3516 14056
rect 3329 14019 3387 14025
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 12066 14056 12072 14068
rect 11572 14028 12072 14056
rect 11572 14016 11578 14028
rect 12066 14016 12072 14028
rect 12124 14056 12130 14068
rect 12805 14059 12863 14065
rect 12805 14056 12817 14059
rect 12124 14028 12817 14056
rect 12124 14016 12130 14028
rect 12805 14025 12817 14028
rect 12851 14025 12863 14059
rect 12805 14019 12863 14025
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 14734 14056 14740 14068
rect 13219 14028 14740 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 15010 14056 15016 14068
rect 14971 14028 15016 14056
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 15197 14059 15255 14065
rect 15197 14025 15209 14059
rect 15243 14056 15255 14059
rect 15286 14056 15292 14068
rect 15243 14028 15292 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 15381 14059 15439 14065
rect 15381 14025 15393 14059
rect 15427 14056 15439 14059
rect 15470 14056 15476 14068
rect 15427 14028 15476 14056
rect 15427 14025 15439 14028
rect 15381 14019 15439 14025
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 17954 14056 17960 14068
rect 15611 14028 17960 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 8110 13988 8116 14000
rect 3068 13960 8116 13988
rect 2777 13951 2835 13957
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 14918 13948 14924 14000
rect 14976 13988 14982 14000
rect 16390 13988 16396 14000
rect 14976 13960 16396 13988
rect 14976 13948 14982 13960
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 16482 13948 16488 14000
rect 16540 13948 16546 14000
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 17083 13960 18460 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 1504 13892 2605 13920
rect 1504 13864 1532 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 2682 13880 2688 13932
rect 2740 13920 2746 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2740 13892 3065 13920
rect 2740 13880 2746 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 3053 13883 3111 13889
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 10502 13920 10508 13932
rect 5684 13892 10508 13920
rect 5684 13880 5690 13892
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 15436 13892 15761 13920
rect 15436 13880 15442 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 16298 13920 16304 13932
rect 16259 13892 16304 13920
rect 15749 13883 15807 13889
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 16500 13920 16528 13948
rect 17129 13923 17187 13929
rect 16500 13892 16896 13920
rect 1486 13852 1492 13864
rect 1447 13824 1492 13852
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 2133 13855 2191 13861
rect 2133 13852 2145 13855
rect 1596 13824 2145 13852
rect 1118 13744 1124 13796
rect 1176 13784 1182 13796
rect 1596 13784 1624 13824
rect 2133 13821 2145 13824
rect 2179 13852 2191 13855
rect 2409 13855 2467 13861
rect 2409 13852 2421 13855
rect 2179 13824 2421 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2409 13821 2421 13824
rect 2455 13821 2467 13855
rect 2409 13815 2467 13821
rect 2516 13824 2774 13852
rect 1176 13756 1624 13784
rect 1857 13787 1915 13793
rect 1176 13744 1182 13756
rect 1857 13753 1869 13787
rect 1903 13784 1915 13787
rect 1946 13784 1952 13796
rect 1903 13756 1952 13784
rect 1903 13753 1915 13756
rect 1857 13747 1915 13753
rect 1946 13744 1952 13756
rect 2004 13744 2010 13796
rect 2516 13784 2544 13824
rect 2240 13756 2544 13784
rect 2746 13784 2774 13824
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 3145 13855 3203 13861
rect 3145 13852 3157 13855
rect 2924 13824 3157 13852
rect 2924 13812 2930 13824
rect 3145 13821 3157 13824
rect 3191 13821 3203 13855
rect 11698 13852 11704 13864
rect 3145 13815 3203 13821
rect 3804 13824 11704 13852
rect 3804 13784 3832 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 12710 13852 12716 13864
rect 12671 13824 12716 13852
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 2746 13756 3832 13784
rect 1581 13719 1639 13725
rect 1581 13685 1593 13719
rect 1627 13716 1639 13719
rect 2240 13716 2268 13756
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 15068 13756 15424 13784
rect 15068 13744 15074 13756
rect 1627 13688 2268 13716
rect 1627 13685 1639 13688
rect 1581 13679 1639 13685
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 2372 13688 2417 13716
rect 2372 13676 2378 13688
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 5074 13716 5080 13728
rect 2648 13688 5080 13716
rect 2648 13676 2654 13688
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 15286 13716 15292 13728
rect 5224 13688 15292 13716
rect 5224 13676 5230 13688
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15396 13716 15424 13756
rect 15838 13744 15844 13796
rect 15896 13784 15902 13796
rect 15896 13756 15941 13784
rect 15896 13744 15902 13756
rect 16022 13744 16028 13796
rect 16080 13784 16086 13796
rect 16592 13784 16620 13892
rect 16080 13756 16620 13784
rect 16868 13784 16896 13892
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17310 13920 17316 13932
rect 17175 13892 17316 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17770 13920 17776 13932
rect 17696 13892 17776 13920
rect 16942 13812 16948 13864
rect 17000 13852 17006 13864
rect 17696 13861 17724 13892
rect 17770 13880 17776 13892
rect 17828 13880 17834 13932
rect 18432 13864 18460 13960
rect 17497 13855 17555 13861
rect 17497 13852 17509 13855
rect 17000 13824 17509 13852
rect 17000 13812 17006 13824
rect 17497 13821 17509 13824
rect 17543 13821 17555 13855
rect 17497 13815 17555 13821
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13821 17739 13855
rect 17862 13852 17868 13864
rect 17823 13824 17868 13852
rect 17681 13815 17739 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 18012 13824 18061 13852
rect 18012 13812 18018 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18414 13852 18420 13864
rect 18375 13824 18420 13852
rect 18049 13815 18107 13821
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 17313 13787 17371 13793
rect 17313 13784 17325 13787
rect 16868 13756 17325 13784
rect 16080 13744 16086 13756
rect 17313 13753 17325 13756
rect 17359 13753 17371 13787
rect 17313 13747 17371 13753
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 17972 13784 18000 13812
rect 17644 13756 18000 13784
rect 17644 13744 17650 13756
rect 18325 13719 18383 13725
rect 18325 13716 18337 13719
rect 15396 13688 18337 13716
rect 18325 13685 18337 13688
rect 18371 13685 18383 13719
rect 18325 13679 18383 13685
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2501 13515 2559 13521
rect 2501 13512 2513 13515
rect 2004 13484 2513 13512
rect 2004 13472 2010 13484
rect 2501 13481 2513 13484
rect 2547 13512 2559 13515
rect 3050 13512 3056 13524
rect 2547 13484 3056 13512
rect 2547 13481 2559 13484
rect 2501 13475 2559 13481
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 3694 13512 3700 13524
rect 3384 13484 3700 13512
rect 3384 13472 3390 13484
rect 3694 13472 3700 13484
rect 3752 13472 3758 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 8527 13484 9505 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 13814 13512 13820 13524
rect 9493 13475 9551 13481
rect 9646 13484 13820 13512
rect 1854 13444 1860 13456
rect 1815 13416 1860 13444
rect 1854 13404 1860 13416
rect 1912 13444 1918 13456
rect 2317 13447 2375 13453
rect 2317 13444 2329 13447
rect 1912 13416 2329 13444
rect 1912 13404 1918 13416
rect 2317 13413 2329 13416
rect 2363 13413 2375 13447
rect 2317 13407 2375 13413
rect 2961 13447 3019 13453
rect 2961 13413 2973 13447
rect 3007 13444 3019 13447
rect 6362 13444 6368 13456
rect 3007 13416 6368 13444
rect 3007 13413 3019 13416
rect 2961 13407 3019 13413
rect 6362 13404 6368 13416
rect 6420 13404 6426 13456
rect 9646 13444 9674 13484
rect 13814 13472 13820 13484
rect 13872 13512 13878 13524
rect 14366 13512 14372 13524
rect 13872 13484 14372 13512
rect 13872 13472 13878 13484
rect 14366 13472 14372 13484
rect 14424 13512 14430 13524
rect 15102 13512 15108 13524
rect 14424 13484 15108 13512
rect 14424 13472 14430 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 15746 13512 15752 13524
rect 15707 13484 15752 13512
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 15838 13472 15844 13524
rect 15896 13512 15902 13524
rect 15979 13515 16037 13521
rect 15979 13512 15991 13515
rect 15896 13484 15991 13512
rect 15896 13472 15902 13484
rect 15979 13481 15991 13484
rect 16025 13481 16037 13515
rect 15979 13475 16037 13481
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13512 16359 13515
rect 16390 13512 16396 13524
rect 16347 13484 16396 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16574 13512 16580 13524
rect 16535 13484 16580 13512
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 17586 13512 17592 13524
rect 16816 13484 17592 13512
rect 16816 13472 16822 13484
rect 17586 13472 17592 13484
rect 17644 13472 17650 13524
rect 6472 13416 9674 13444
rect 1486 13376 1492 13388
rect 1447 13348 1492 13376
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 3326 13376 3332 13388
rect 2087 13348 3332 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 3326 13336 3332 13348
rect 3384 13336 3390 13388
rect 4706 13376 4712 13388
rect 4667 13348 4712 13376
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13376 4859 13379
rect 4982 13376 4988 13388
rect 4847 13348 4988 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5074 13336 5080 13388
rect 5132 13376 5138 13388
rect 6472 13376 6500 13416
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 11572 13416 15148 13444
rect 11572 13404 11578 13416
rect 5132 13348 6500 13376
rect 5132 13336 5138 13348
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 7018 13379 7076 13385
rect 7018 13376 7030 13379
rect 6696 13348 7030 13376
rect 6696 13336 6702 13348
rect 7018 13345 7030 13348
rect 7064 13345 7076 13379
rect 8386 13376 8392 13388
rect 8347 13348 8392 13376
rect 7018 13339 7076 13345
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13376 9919 13379
rect 11882 13376 11888 13388
rect 9907 13348 11888 13376
rect 9907 13345 9919 13348
rect 9861 13339 9919 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 14734 13376 14740 13388
rect 14695 13348 14740 13376
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 15120 13376 15148 13416
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 15252 13416 16536 13444
rect 15252 13404 15258 13416
rect 16082 13379 16140 13385
rect 15120 13348 15884 13376
rect 1504 13308 1532 13336
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 1504 13280 2145 13308
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 2133 13271 2191 13277
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13308 2835 13311
rect 3050 13308 3056 13320
rect 2823 13280 3056 13308
rect 2823 13277 2835 13280
rect 2777 13271 2835 13277
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 7285 13311 7343 13317
rect 4948 13280 4993 13308
rect 4948 13268 4954 13280
rect 7285 13277 7297 13311
rect 7331 13308 7343 13311
rect 7466 13308 7472 13320
rect 7331 13280 7472 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7466 13268 7472 13280
rect 7524 13308 7530 13320
rect 8018 13308 8024 13320
rect 7524 13280 8024 13308
rect 7524 13268 7530 13280
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8846 13308 8852 13320
rect 8711 13280 8852 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 9640 13280 9965 13308
rect 9640 13268 9646 13280
rect 9953 13277 9965 13280
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 3234 13240 3240 13252
rect 2746 13212 3240 13240
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2746 13172 2774 13212
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 4249 13243 4307 13249
rect 4249 13209 4261 13243
rect 4295 13240 4307 13243
rect 4614 13240 4620 13252
rect 4295 13212 4620 13240
rect 4295 13209 4307 13212
rect 4249 13203 4307 13209
rect 4614 13200 4620 13212
rect 4672 13200 4678 13252
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 10060 13240 10088 13271
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 13412 13280 14473 13308
rect 13412 13268 13418 13280
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13308 14703 13311
rect 15654 13308 15660 13320
rect 14691 13280 15660 13308
rect 14691 13277 14703 13280
rect 14645 13271 14703 13277
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 8536 13212 10088 13240
rect 10244 13212 12434 13240
rect 8536 13200 8542 13212
rect 3418 13172 3424 13184
rect 1627 13144 2774 13172
rect 3379 13144 3424 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 4338 13172 4344 13184
rect 4299 13144 4344 13172
rect 4338 13132 4344 13144
rect 4396 13132 4402 13184
rect 5258 13172 5264 13184
rect 5219 13144 5264 13172
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5902 13172 5908 13184
rect 5863 13144 5908 13172
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 8021 13175 8079 13181
rect 8021 13141 8033 13175
rect 8067 13172 8079 13175
rect 8938 13172 8944 13184
rect 8067 13144 8944 13172
rect 8067 13141 8079 13144
rect 8021 13135 8079 13141
rect 8938 13132 8944 13144
rect 8996 13132 9002 13184
rect 9214 13172 9220 13184
rect 9127 13144 9220 13172
rect 9214 13132 9220 13144
rect 9272 13172 9278 13184
rect 10244 13172 10272 13212
rect 11514 13172 11520 13184
rect 9272 13144 10272 13172
rect 11475 13144 11520 13172
rect 9272 13132 9278 13144
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 12406 13172 12434 13212
rect 14090 13200 14096 13252
rect 14148 13240 14154 13252
rect 14550 13240 14556 13252
rect 14148 13212 14556 13240
rect 14148 13200 14154 13212
rect 14550 13200 14556 13212
rect 14608 13240 14614 13252
rect 14826 13240 14832 13252
rect 14608 13212 14832 13240
rect 14608 13200 14614 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 15105 13243 15163 13249
rect 15105 13209 15117 13243
rect 15151 13240 15163 13243
rect 15286 13240 15292 13252
rect 15151 13212 15292 13240
rect 15151 13209 15163 13212
rect 15105 13203 15163 13209
rect 15286 13200 15292 13212
rect 15344 13200 15350 13252
rect 15378 13200 15384 13252
rect 15436 13240 15442 13252
rect 15856 13240 15884 13348
rect 16082 13345 16094 13379
rect 16128 13376 16140 13379
rect 16206 13376 16212 13388
rect 16128 13348 16212 13376
rect 16128 13345 16140 13348
rect 16082 13339 16140 13345
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 16508 13385 16536 13416
rect 17034 13404 17040 13456
rect 17092 13444 17098 13456
rect 18969 13447 19027 13453
rect 18969 13444 18981 13447
rect 17092 13416 17137 13444
rect 18064 13416 18981 13444
rect 17092 13404 17098 13416
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13345 16543 13379
rect 16485 13339 16543 13345
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13345 17003 13379
rect 17678 13376 17684 13388
rect 17639 13348 17684 13376
rect 16945 13339 17003 13345
rect 16390 13268 16396 13320
rect 16448 13308 16454 13320
rect 16960 13308 16988 13339
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 18064 13385 18092 13416
rect 18969 13413 18981 13416
rect 19015 13413 19027 13447
rect 18969 13407 19027 13413
rect 18049 13379 18107 13385
rect 18049 13376 18061 13379
rect 17788 13348 18061 13376
rect 17126 13308 17132 13320
rect 16448 13280 16988 13308
rect 17087 13280 17132 13308
rect 16448 13268 16454 13280
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13308 17463 13311
rect 17788 13308 17816 13348
rect 18049 13345 18061 13348
rect 18095 13345 18107 13379
rect 18414 13376 18420 13388
rect 18375 13348 18420 13376
rect 18049 13339 18107 13345
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 17451 13280 17816 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18233 13311 18291 13317
rect 18233 13308 18245 13311
rect 18012 13280 18245 13308
rect 18012 13268 18018 13280
rect 18233 13277 18245 13280
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 17865 13243 17923 13249
rect 17865 13240 17877 13243
rect 15436 13212 15481 13240
rect 15856 13212 17877 13240
rect 15436 13200 15442 13212
rect 17865 13209 17877 13212
rect 17911 13209 17923 13243
rect 17865 13203 17923 13209
rect 15010 13172 15016 13184
rect 12406 13144 15016 13172
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 15657 13175 15715 13181
rect 15657 13141 15669 13175
rect 15703 13172 15715 13175
rect 17405 13175 17463 13181
rect 17405 13172 17417 13175
rect 15703 13144 17417 13172
rect 15703 13141 15715 13144
rect 15657 13135 15715 13141
rect 17405 13141 17417 13144
rect 17451 13141 17463 13175
rect 17586 13172 17592 13184
rect 17547 13144 17592 13172
rect 17405 13135 17463 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 1995 12940 4660 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12900 1731 12903
rect 4632 12900 4660 12940
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4764 12940 4813 12968
rect 4764 12928 4770 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 6638 12968 6644 12980
rect 6599 12940 6644 12968
rect 4801 12931 4859 12937
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 8294 12968 8300 12980
rect 6748 12940 8300 12968
rect 6748 12900 6776 12940
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8478 12968 8484 12980
rect 8439 12940 8484 12968
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 12342 12968 12348 12980
rect 11931 12940 12348 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 14645 12971 14703 12977
rect 12544 12940 13860 12968
rect 8110 12900 8116 12912
rect 1719 12872 2774 12900
rect 4632 12872 6776 12900
rect 8071 12872 8116 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 2133 12835 2191 12841
rect 2133 12832 2145 12835
rect 1452 12804 2145 12832
rect 1452 12792 1458 12804
rect 2133 12801 2145 12804
rect 2179 12801 2191 12835
rect 2746 12832 2774 12872
rect 8110 12860 8116 12872
rect 8168 12900 8174 12912
rect 8570 12900 8576 12912
rect 8168 12872 8576 12900
rect 8168 12860 8174 12872
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 11146 12860 11152 12912
rect 11204 12900 11210 12912
rect 12544 12900 12572 12940
rect 11204 12872 12572 12900
rect 13832 12900 13860 12940
rect 14645 12937 14657 12971
rect 14691 12968 14703 12971
rect 14734 12968 14740 12980
rect 14691 12940 14740 12968
rect 14691 12937 14703 12940
rect 14645 12931 14703 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 14884 12940 15577 12968
rect 14884 12928 14890 12940
rect 15565 12937 15577 12940
rect 15611 12937 15623 12971
rect 15565 12931 15623 12937
rect 15654 12928 15660 12980
rect 15712 12968 15718 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15712 12940 15853 12968
rect 15712 12928 15718 12940
rect 15841 12937 15853 12940
rect 15887 12937 15899 12971
rect 15841 12931 15899 12937
rect 16206 12928 16212 12980
rect 16264 12968 16270 12980
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 16264 12940 18337 12968
rect 16264 12928 16270 12940
rect 18325 12937 18337 12940
rect 18371 12937 18383 12971
rect 18325 12931 18383 12937
rect 13832 12872 13952 12900
rect 11204 12860 11210 12872
rect 4617 12835 4675 12841
rect 2746 12804 3096 12832
rect 2133 12795 2191 12801
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 1504 12736 2513 12764
rect 1504 12708 1532 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 2924 12736 2973 12764
rect 2924 12724 2930 12736
rect 2961 12733 2973 12736
rect 3007 12733 3019 12767
rect 3068 12764 3096 12804
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5074 12832 5080 12844
rect 4663 12804 5080 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 5534 12832 5540 12844
rect 5491 12804 5540 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5534 12792 5540 12804
rect 5592 12832 5598 12844
rect 5902 12832 5908 12844
rect 5592 12804 5908 12832
rect 5592 12792 5598 12804
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 8018 12832 8024 12844
rect 7979 12804 8024 12832
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 3068 12736 7696 12764
rect 2961 12727 3019 12733
rect 1486 12696 1492 12708
rect 1447 12668 1492 12696
rect 1486 12656 1492 12668
rect 1544 12656 1550 12708
rect 1854 12696 1860 12708
rect 1815 12668 1860 12696
rect 1854 12656 1860 12668
rect 1912 12696 1918 12708
rect 2685 12699 2743 12705
rect 2685 12696 2697 12699
rect 1912 12668 2697 12696
rect 1912 12656 1918 12668
rect 2685 12665 2697 12668
rect 2731 12665 2743 12699
rect 2685 12659 2743 12665
rect 3228 12699 3286 12705
rect 3228 12665 3240 12699
rect 3274 12696 3286 12699
rect 3510 12696 3516 12708
rect 3274 12668 3516 12696
rect 3274 12665 3286 12668
rect 3228 12659 3286 12665
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 5169 12699 5227 12705
rect 5169 12665 5181 12699
rect 5215 12696 5227 12699
rect 5629 12699 5687 12705
rect 5629 12696 5641 12699
rect 5215 12668 5641 12696
rect 5215 12665 5227 12668
rect 5169 12659 5227 12665
rect 5629 12665 5641 12668
rect 5675 12665 5687 12699
rect 5629 12659 5687 12665
rect 5810 12656 5816 12708
rect 5868 12696 5874 12708
rect 6181 12699 6239 12705
rect 6181 12696 6193 12699
rect 5868 12668 6193 12696
rect 5868 12656 5874 12668
rect 6181 12665 6193 12668
rect 6227 12665 6239 12699
rect 6181 12659 6239 12665
rect 6362 12656 6368 12708
rect 6420 12696 6426 12708
rect 7668 12696 7696 12736
rect 7742 12724 7748 12776
rect 7800 12773 7806 12776
rect 7800 12764 7812 12773
rect 8389 12767 8447 12773
rect 7800 12736 7845 12764
rect 7800 12727 7812 12736
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 9861 12767 9919 12773
rect 8435 12736 9720 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 7800 12724 7806 12727
rect 6420 12668 7604 12696
rect 7668 12668 8708 12696
rect 6420 12656 6426 12668
rect 2222 12588 2228 12640
rect 2280 12628 2286 12640
rect 2317 12631 2375 12637
rect 2317 12628 2329 12631
rect 2280 12600 2329 12628
rect 2280 12588 2286 12600
rect 2317 12597 2329 12600
rect 2363 12597 2375 12631
rect 2317 12591 2375 12597
rect 4341 12631 4399 12637
rect 4341 12597 4353 12631
rect 4387 12628 4399 12631
rect 4430 12628 4436 12640
rect 4387 12600 4436 12628
rect 4387 12597 4399 12600
rect 4341 12591 4399 12597
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5718 12628 5724 12640
rect 5307 12600 5724 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5718 12588 5724 12600
rect 5776 12628 5782 12640
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5776 12600 5917 12628
rect 5776 12588 5782 12600
rect 5905 12597 5917 12600
rect 5951 12597 5963 12631
rect 6546 12628 6552 12640
rect 6507 12600 6552 12628
rect 5905 12591 5963 12597
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 7576 12628 7604 12668
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 7576 12600 8401 12628
rect 8389 12597 8401 12600
rect 8435 12597 8447 12631
rect 8680 12628 8708 12668
rect 9490 12656 9496 12708
rect 9548 12696 9554 12708
rect 9594 12699 9652 12705
rect 9594 12696 9606 12699
rect 9548 12668 9606 12696
rect 9548 12656 9554 12668
rect 9594 12665 9606 12668
rect 9640 12665 9652 12699
rect 9692 12696 9720 12736
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 10410 12764 10416 12776
rect 9907 12736 10416 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 11701 12767 11759 12773
rect 11701 12764 11713 12767
rect 10744 12736 11713 12764
rect 10744 12724 10750 12736
rect 11701 12733 11713 12736
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 13193 12767 13251 12773
rect 13193 12733 13205 12767
rect 13239 12764 13251 12767
rect 13354 12764 13360 12776
rect 13239 12736 13360 12764
rect 13239 12733 13251 12736
rect 13193 12727 13251 12733
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13449 12767 13507 12773
rect 13449 12733 13461 12767
rect 13495 12733 13507 12767
rect 13924 12764 13952 12872
rect 13998 12860 14004 12912
rect 14056 12900 14062 12912
rect 14056 12872 17632 12900
rect 14056 12860 14062 12872
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 15611 12804 16405 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 16393 12801 16405 12804
rect 16439 12801 16451 12835
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16393 12795 16451 12801
rect 15396 12764 15424 12795
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12832 17187 12835
rect 17494 12832 17500 12844
rect 17175 12804 17500 12832
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 15654 12764 15660 12776
rect 13924 12736 15332 12764
rect 15396 12736 15660 12764
rect 13449 12727 13507 12733
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 9692 12668 11069 12696
rect 9594 12659 9652 12665
rect 11057 12665 11069 12668
rect 11103 12696 11115 12699
rect 11514 12696 11520 12708
rect 11103 12668 11520 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 8680 12600 10517 12628
rect 8389 12591 8447 12597
rect 10505 12597 10517 12600
rect 10551 12628 10563 12631
rect 10594 12628 10600 12640
rect 10551 12600 10600 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 10594 12588 10600 12600
rect 10652 12628 10658 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10652 12600 10977 12628
rect 10652 12588 10658 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 11422 12628 11428 12640
rect 11383 12600 11428 12628
rect 10965 12591 11023 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 12066 12628 12072 12640
rect 12027 12600 12072 12628
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 13464 12628 13492 12727
rect 13633 12699 13691 12705
rect 13633 12665 13645 12699
rect 13679 12696 13691 12699
rect 13998 12696 14004 12708
rect 13679 12668 14004 12696
rect 13679 12665 13691 12668
rect 13633 12659 13691 12665
rect 13998 12656 14004 12668
rect 14056 12656 14062 12708
rect 14185 12699 14243 12705
rect 14185 12665 14197 12699
rect 14231 12696 14243 12699
rect 15102 12696 15108 12708
rect 14231 12668 14780 12696
rect 15063 12668 15108 12696
rect 14231 12665 14243 12668
rect 14185 12659 14243 12665
rect 14090 12628 14096 12640
rect 13464 12600 14096 12628
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 14752 12637 14780 12668
rect 15102 12656 15108 12668
rect 15160 12656 15166 12708
rect 14737 12631 14795 12637
rect 14332 12600 14377 12628
rect 14332 12588 14338 12600
rect 14737 12597 14749 12631
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 14918 12588 14924 12640
rect 14976 12628 14982 12640
rect 15197 12631 15255 12637
rect 15197 12628 15209 12631
rect 14976 12600 15209 12628
rect 14976 12588 14982 12600
rect 15197 12597 15209 12600
rect 15243 12597 15255 12631
rect 15304 12628 15332 12736
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 16209 12767 16267 12773
rect 16209 12733 16221 12767
rect 16255 12764 16267 12767
rect 16574 12764 16580 12776
rect 16255 12736 16580 12764
rect 16255 12733 16267 12736
rect 16209 12727 16267 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 17604 12773 17632 12872
rect 17770 12832 17776 12844
rect 17731 12804 17776 12832
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 17589 12767 17647 12773
rect 17589 12733 17601 12767
rect 17635 12733 17647 12767
rect 17589 12727 17647 12733
rect 18141 12767 18199 12773
rect 18141 12733 18153 12767
rect 18187 12764 18199 12767
rect 18506 12764 18512 12776
rect 18187 12736 18512 12764
rect 18187 12733 18199 12736
rect 18141 12727 18199 12733
rect 18506 12724 18512 12736
rect 18564 12724 18570 12776
rect 15470 12656 15476 12708
rect 15528 12696 15534 12708
rect 16301 12699 16359 12705
rect 16301 12696 16313 12699
rect 15528 12668 16313 12696
rect 15528 12656 15534 12668
rect 16301 12665 16313 12668
rect 16347 12665 16359 12699
rect 17681 12699 17739 12705
rect 17681 12696 17693 12699
rect 16301 12659 16359 12665
rect 16408 12668 17693 12696
rect 15657 12631 15715 12637
rect 15657 12628 15669 12631
rect 15304 12600 15669 12628
rect 15197 12591 15255 12597
rect 15657 12597 15669 12600
rect 15703 12628 15715 12631
rect 16408 12628 16436 12668
rect 17681 12665 17693 12668
rect 17727 12665 17739 12699
rect 17681 12659 17739 12665
rect 15703 12600 16436 12628
rect 15703 12597 15715 12600
rect 15657 12591 15715 12597
rect 16482 12588 16488 12640
rect 16540 12628 16546 12640
rect 17221 12631 17279 12637
rect 17221 12628 17233 12631
rect 16540 12600 17233 12628
rect 16540 12588 16546 12600
rect 17221 12597 17233 12600
rect 17267 12597 17279 12631
rect 17221 12591 17279 12597
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 18966 12492 18972 12504
rect 1104 12464 18860 12486
rect 18927 12464 18972 12492
rect 18966 12452 18972 12464
rect 19024 12452 19030 12504
rect 3510 12424 3516 12436
rect 3423 12396 3516 12424
rect 3510 12384 3516 12396
rect 3568 12424 3574 12436
rect 4890 12424 4896 12436
rect 3568 12396 4896 12424
rect 3568 12384 3574 12396
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 5074 12424 5080 12436
rect 5035 12396 5080 12424
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 5169 12427 5227 12433
rect 5169 12393 5181 12427
rect 5215 12424 5227 12427
rect 5997 12427 6055 12433
rect 5215 12396 5672 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5644 12365 5672 12396
rect 5997 12393 6009 12427
rect 6043 12424 6055 12427
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 6043 12396 6561 12424
rect 6043 12393 6055 12396
rect 5997 12387 6055 12393
rect 6549 12393 6561 12396
rect 6595 12424 6607 12427
rect 6730 12424 6736 12436
rect 6595 12396 6736 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 7653 12427 7711 12433
rect 7653 12393 7665 12427
rect 7699 12424 7711 12427
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 7699 12396 8217 12424
rect 7699 12393 7711 12396
rect 7653 12387 7711 12393
rect 8205 12393 8217 12396
rect 8251 12393 8263 12427
rect 8570 12424 8576 12436
rect 8531 12396 8576 12424
rect 8205 12387 8263 12393
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9582 12424 9588 12436
rect 9543 12396 9588 12424
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12345 12427 12403 12433
rect 12345 12424 12357 12427
rect 11992 12396 12357 12424
rect 5629 12359 5687 12365
rect 2746 12328 5304 12356
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 1489 12291 1547 12297
rect 1489 12288 1501 12291
rect 1452 12260 1501 12288
rect 1452 12248 1458 12260
rect 1489 12257 1501 12260
rect 1535 12257 1547 12291
rect 1489 12251 1547 12257
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 2222 12288 2228 12300
rect 1903 12260 2228 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 2400 12291 2458 12297
rect 2400 12257 2412 12291
rect 2446 12288 2458 12291
rect 2746 12288 2774 12328
rect 2446 12260 2774 12288
rect 2446 12257 2458 12260
rect 2400 12251 2458 12257
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 3694 12288 3700 12300
rect 3568 12260 3700 12288
rect 3568 12248 3574 12260
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12288 4307 12291
rect 4706 12288 4712 12300
rect 4295 12260 4712 12288
rect 4295 12257 4307 12260
rect 4249 12251 4307 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 3878 12220 3884 12232
rect 3651 12192 3884 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2148 12084 2176 12183
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 4890 12220 4896 12232
rect 4571 12192 4896 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 2866 12084 2872 12096
rect 2148 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12084 2930 12096
rect 3694 12084 3700 12096
rect 2924 12056 3700 12084
rect 2924 12044 2930 12056
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4246 12084 4252 12096
rect 3927 12056 4252 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4356 12084 4384 12183
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5276 12229 5304 12328
rect 5629 12325 5641 12359
rect 5675 12356 5687 12359
rect 7282 12356 7288 12368
rect 5675 12328 7288 12356
rect 5675 12325 5687 12328
rect 5629 12319 5687 12325
rect 7282 12316 7288 12328
rect 7340 12316 7346 12368
rect 7742 12356 7748 12368
rect 7703 12328 7748 12356
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 9398 12356 9404 12368
rect 8404 12328 9404 12356
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12288 6515 12291
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6503 12260 7021 12288
rect 6503 12257 6515 12260
rect 6457 12251 6515 12257
rect 7009 12257 7021 12260
rect 7055 12288 7067 12291
rect 8404 12288 8432 12328
rect 9398 12316 9404 12328
rect 9456 12316 9462 12368
rect 9490 12316 9496 12368
rect 9548 12356 9554 12368
rect 10680 12359 10738 12365
rect 9548 12328 10272 12356
rect 9548 12316 9554 12328
rect 9508 12288 9536 12316
rect 7055 12260 8432 12288
rect 8864 12260 9536 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12220 5319 12223
rect 5534 12220 5540 12232
rect 5307 12192 5540 12220
rect 5307 12189 5319 12192
rect 5261 12183 5319 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 7561 12223 7619 12229
rect 6696 12192 6741 12220
rect 6696 12180 6702 12192
rect 7561 12189 7573 12223
rect 7607 12220 7619 12223
rect 8478 12220 8484 12232
rect 7607 12192 8484 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8662 12220 8668 12232
rect 8623 12192 8668 12220
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8864 12229 8892 12260
rect 9766 12248 9772 12300
rect 9824 12288 9830 12300
rect 9953 12291 10011 12297
rect 9953 12288 9965 12291
rect 9824 12260 9965 12288
rect 9824 12248 9830 12260
rect 9953 12257 9965 12260
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 10244 12288 10272 12328
rect 10680 12325 10692 12359
rect 10726 12356 10738 12359
rect 10778 12356 10784 12368
rect 10726 12328 10784 12356
rect 10726 12325 10738 12328
rect 10680 12319 10738 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11422 12316 11428 12368
rect 11480 12356 11486 12368
rect 11992 12356 12020 12396
rect 12345 12393 12357 12396
rect 12391 12393 12403 12427
rect 12345 12387 12403 12393
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 13354 12424 13360 12436
rect 12851 12396 13360 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 17862 12424 17868 12436
rect 13832 12396 17868 12424
rect 11480 12328 12020 12356
rect 11480 12316 11486 12328
rect 12066 12316 12072 12368
rect 12124 12356 12130 12368
rect 13262 12356 13268 12368
rect 12124 12328 13268 12356
rect 12124 12316 12130 12328
rect 13262 12316 13268 12328
rect 13320 12356 13326 12368
rect 13832 12356 13860 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18141 12427 18199 12433
rect 18141 12393 18153 12427
rect 18187 12424 18199 12427
rect 18414 12424 18420 12436
rect 18187 12396 18420 12424
rect 18187 12393 18199 12396
rect 18141 12387 18199 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 13320 12328 13860 12356
rect 13940 12359 13998 12365
rect 13320 12316 13326 12328
rect 13940 12325 13952 12359
rect 13986 12356 13998 12359
rect 14550 12356 14556 12368
rect 13986 12328 14556 12356
rect 13986 12325 13998 12328
rect 13940 12319 13998 12325
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 15286 12316 15292 12368
rect 15344 12356 15350 12368
rect 15654 12356 15660 12368
rect 15344 12328 15660 12356
rect 15344 12316 15350 12328
rect 15654 12316 15660 12328
rect 15712 12356 15718 12368
rect 15964 12359 16022 12365
rect 15964 12356 15976 12359
rect 15712 12328 15976 12356
rect 15712 12316 15718 12328
rect 15964 12325 15976 12328
rect 16010 12356 16022 12359
rect 16574 12356 16580 12368
rect 16010 12328 16580 12356
rect 16010 12325 16022 12328
rect 15964 12319 16022 12325
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 16850 12316 16856 12368
rect 16908 12356 16914 12368
rect 17310 12356 17316 12368
rect 16908 12328 17316 12356
rect 16908 12316 16914 12328
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 17512 12328 18460 12356
rect 10244 12260 11836 12288
rect 8849 12223 8907 12229
rect 8849 12189 8861 12223
rect 8895 12189 8907 12223
rect 9306 12220 9312 12232
rect 9267 12192 9312 12220
rect 8849 12183 8907 12189
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 10244 12229 10272 12260
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 10229 12183 10287 12189
rect 4709 12155 4767 12161
rect 4709 12121 4721 12155
rect 4755 12152 4767 12155
rect 4982 12152 4988 12164
rect 4755 12124 4988 12152
rect 4755 12121 4767 12124
rect 4709 12115 4767 12121
rect 4982 12112 4988 12124
rect 5040 12112 5046 12164
rect 6178 12112 6184 12164
rect 6236 12152 6242 12164
rect 8113 12155 8171 12161
rect 6236 12124 7328 12152
rect 6236 12112 6242 12124
rect 5442 12084 5448 12096
rect 4356 12056 5448 12084
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5810 12084 5816 12096
rect 5771 12056 5816 12084
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6089 12087 6147 12093
rect 6089 12084 6101 12087
rect 6052 12056 6101 12084
rect 6052 12044 6058 12056
rect 6089 12053 6101 12056
rect 6135 12053 6147 12087
rect 6089 12047 6147 12053
rect 6822 12044 6828 12096
rect 6880 12084 6886 12096
rect 7193 12087 7251 12093
rect 7193 12084 7205 12087
rect 6880 12056 7205 12084
rect 6880 12044 6886 12056
rect 7193 12053 7205 12056
rect 7239 12053 7251 12087
rect 7300 12084 7328 12124
rect 8113 12121 8125 12155
rect 8159 12152 8171 12155
rect 8386 12152 8392 12164
rect 8159 12124 8392 12152
rect 8159 12121 8171 12124
rect 8113 12115 8171 12121
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 9401 12155 9459 12161
rect 8496 12124 9352 12152
rect 8496 12084 8524 12124
rect 7300 12056 8524 12084
rect 7193 12047 7251 12053
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 9214 12084 9220 12096
rect 8720 12056 9220 12084
rect 8720 12044 8726 12056
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9324 12084 9352 12124
rect 9401 12121 9413 12155
rect 9447 12152 9459 12155
rect 9582 12152 9588 12164
rect 9447 12124 9588 12152
rect 9447 12121 9459 12124
rect 9401 12115 9459 12121
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 10060 12152 10088 12183
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 11808 12220 11836 12260
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 12253 12291 12311 12297
rect 12253 12288 12265 12291
rect 11940 12260 12265 12288
rect 11940 12248 11946 12260
rect 12253 12257 12265 12260
rect 12299 12257 12311 12291
rect 12253 12251 12311 12257
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 16393 12291 16451 12297
rect 12584 12260 16344 12288
rect 12584 12248 12590 12260
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 11808 12192 12449 12220
rect 10318 12152 10324 12164
rect 10060 12124 10324 12152
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 11808 12161 11836 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 14182 12220 14188 12232
rect 14143 12192 14188 12220
rect 12437 12183 12495 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 14734 12220 14740 12232
rect 14695 12192 14740 12220
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16316 12220 16344 12260
rect 16393 12257 16405 12291
rect 16439 12288 16451 12291
rect 17512 12288 17540 12328
rect 16439 12260 17540 12288
rect 17609 12291 17667 12297
rect 16439 12257 16451 12260
rect 16393 12251 16451 12257
rect 17609 12257 17621 12291
rect 17655 12288 17667 12291
rect 17770 12288 17776 12300
rect 17655 12260 17776 12288
rect 17655 12257 17667 12260
rect 17609 12251 17667 12257
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 18432 12297 18460 12328
rect 18417 12291 18475 12297
rect 18417 12257 18429 12291
rect 18463 12288 18475 12291
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 18463 12260 18981 12288
rect 18463 12257 18475 12260
rect 18417 12251 18475 12257
rect 18969 12257 18981 12260
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 16850 12220 16856 12232
rect 16316 12192 16856 12220
rect 16209 12183 16267 12189
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12121 11851 12155
rect 11793 12115 11851 12121
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 14829 12155 14887 12161
rect 14829 12152 14841 12155
rect 14608 12124 14841 12152
rect 14608 12112 14614 12124
rect 14829 12121 14841 12124
rect 14875 12121 14887 12155
rect 14829 12115 14887 12121
rect 16224 12096 16252 12183
rect 16850 12180 16856 12192
rect 16908 12180 16914 12232
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 16485 12155 16543 12161
rect 16485 12121 16497 12155
rect 16531 12152 16543 12155
rect 16574 12152 16580 12164
rect 16531 12124 16580 12152
rect 16531 12121 16543 12124
rect 16485 12115 16543 12121
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 12066 12084 12072 12096
rect 9324 12056 12072 12084
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 13906 12044 13912 12096
rect 13964 12084 13970 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 13964 12056 14381 12084
rect 13964 12044 13970 12056
rect 14369 12053 14381 12056
rect 14415 12084 14427 12087
rect 14918 12084 14924 12096
rect 14415 12056 14924 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15102 12044 15108 12096
rect 15160 12084 15166 12096
rect 16206 12084 16212 12096
rect 15160 12056 16212 12084
rect 15160 12044 15166 12056
rect 16206 12044 16212 12056
rect 16264 12084 16270 12096
rect 17880 12084 17908 12183
rect 18322 12084 18328 12096
rect 16264 12056 17908 12084
rect 18283 12056 18328 12084
rect 16264 12044 16270 12056
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 1946 11840 1952 11892
rect 2004 11880 2010 11892
rect 3513 11883 3571 11889
rect 2004 11852 2774 11880
rect 2004 11840 2010 11852
rect 2746 11812 2774 11852
rect 3513 11849 3525 11883
rect 3559 11880 3571 11883
rect 3602 11880 3608 11892
rect 3559 11852 3608 11880
rect 3559 11849 3571 11852
rect 3513 11843 3571 11849
rect 3602 11840 3608 11852
rect 3660 11880 3666 11892
rect 4706 11880 4712 11892
rect 3660 11852 4568 11880
rect 4667 11852 4712 11880
rect 3660 11840 3666 11852
rect 4430 11812 4436 11824
rect 2746 11784 3188 11812
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2774 11744 2780 11756
rect 2271 11716 2780 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 1762 11608 1768 11620
rect 1723 11580 1768 11608
rect 1762 11568 1768 11580
rect 1820 11568 1826 11620
rect 2038 11608 2044 11620
rect 1999 11580 2044 11608
rect 2038 11568 2044 11580
rect 2096 11608 2102 11620
rect 3053 11611 3111 11617
rect 3053 11608 3065 11611
rect 2096 11580 3065 11608
rect 2096 11568 2102 11580
rect 3053 11577 3065 11580
rect 3099 11577 3111 11611
rect 3160 11608 3188 11784
rect 4080 11784 4436 11812
rect 4080 11753 4108 11784
rect 4430 11772 4436 11784
rect 4488 11772 4494 11824
rect 4540 11812 4568 11852
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 5500 11852 5549 11880
rect 5500 11840 5506 11852
rect 5537 11849 5549 11852
rect 5583 11849 5595 11883
rect 8846 11880 8852 11892
rect 5537 11843 5595 11849
rect 5644 11852 8432 11880
rect 8807 11852 8852 11880
rect 5644 11812 5672 11852
rect 4540 11784 5672 11812
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6730 11812 6736 11824
rect 6420 11784 6736 11812
rect 6420 11772 6426 11784
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 8404 11812 8432 11852
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 8996 11852 9041 11880
rect 8996 11840 9002 11852
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9824 11852 9873 11880
rect 9824 11840 9830 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 10376 11852 10701 11880
rect 10376 11840 10382 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11563 11852 11989 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11977 11849 11989 11852
rect 12023 11880 12035 11883
rect 12023 11852 12480 11880
rect 12023 11849 12035 11852
rect 11977 11843 12035 11849
rect 11882 11812 11888 11824
rect 8404 11784 11888 11812
rect 11882 11772 11888 11784
rect 11940 11772 11946 11824
rect 12452 11812 12480 11852
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 12584 11852 13461 11880
rect 12584 11840 12590 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13449 11843 13507 11849
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14332 11852 14381 11880
rect 14332 11840 14338 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14826 11880 14832 11892
rect 14369 11843 14427 11849
rect 14476 11852 14832 11880
rect 13814 11812 13820 11824
rect 12452 11784 13820 11812
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 13909 11815 13967 11821
rect 13909 11781 13921 11815
rect 13955 11812 13967 11815
rect 14090 11812 14096 11824
rect 13955 11784 14096 11812
rect 13955 11781 13967 11784
rect 13909 11775 13967 11781
rect 14090 11772 14096 11784
rect 14148 11812 14154 11824
rect 14476 11812 14504 11852
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 15528 11852 15945 11880
rect 15528 11840 15534 11852
rect 15933 11849 15945 11852
rect 15979 11849 15991 11883
rect 16666 11880 16672 11892
rect 15933 11843 15991 11849
rect 16132 11852 16672 11880
rect 14148 11784 14504 11812
rect 14148 11772 14154 11784
rect 14550 11772 14556 11824
rect 14608 11812 14614 11824
rect 16022 11812 16028 11824
rect 14608 11784 16028 11812
rect 14608 11772 14614 11784
rect 16022 11772 16028 11784
rect 16080 11772 16086 11824
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4246 11744 4252 11756
rect 4203 11716 4252 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11744 5411 11747
rect 5534 11744 5540 11756
rect 5399 11716 5540 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 5534 11704 5540 11716
rect 5592 11744 5598 11756
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5592 11716 6101 11744
rect 5592 11704 5598 11716
rect 6089 11713 6101 11716
rect 6135 11713 6147 11747
rect 6089 11707 6147 11713
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6696 11716 7021 11744
rect 6696 11704 6702 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 9490 11744 9496 11756
rect 9451 11716 9496 11744
rect 7009 11707 7067 11713
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 10778 11744 10784 11756
rect 10551 11716 10784 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 10778 11704 10784 11716
rect 10836 11744 10842 11756
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 10836 11716 11253 11744
rect 10836 11704 10842 11716
rect 11241 11713 11253 11716
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12124 11716 13001 11744
rect 12124 11704 12130 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 14829 11747 14887 11753
rect 14829 11744 14841 11747
rect 13688 11716 14841 11744
rect 13688 11704 13694 11716
rect 14829 11713 14841 11716
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 15286 11744 15292 11756
rect 15059 11716 15292 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3292 11648 3801 11676
rect 3292 11636 3298 11648
rect 3789 11645 3801 11648
rect 3835 11676 3847 11679
rect 4798 11676 4804 11688
rect 3835 11648 4804 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 5994 11676 6000 11688
rect 5951 11648 6000 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 6822 11676 6828 11688
rect 6420 11648 6828 11676
rect 6420 11636 6426 11648
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7466 11676 7472 11688
rect 7427 11648 7472 11676
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 7736 11679 7794 11685
rect 7736 11645 7748 11679
rect 7782 11676 7794 11679
rect 8478 11676 8484 11688
rect 7782 11648 8484 11676
rect 7782 11645 7794 11648
rect 7736 11639 7794 11645
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 9306 11676 9312 11688
rect 9267 11648 9312 11676
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 10226 11676 10232 11688
rect 9456 11648 10232 11676
rect 9456 11636 9462 11648
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11103 11648 11529 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 12250 11676 12256 11688
rect 12211 11648 12256 11676
rect 11517 11639 11575 11645
rect 12250 11636 12256 11648
rect 12308 11676 12314 11688
rect 14550 11676 14556 11688
rect 12308 11648 14556 11676
rect 12308 11636 12314 11648
rect 14550 11636 14556 11648
rect 14608 11636 14614 11688
rect 14734 11676 14740 11688
rect 14695 11648 14740 11676
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 14844 11676 14872 11707
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 16132 11744 16160 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 16761 11883 16819 11889
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 17034 11880 17040 11892
rect 16807 11852 17040 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17494 11880 17500 11892
rect 17368 11852 17500 11880
rect 17368 11840 17374 11852
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 18046 11880 18052 11892
rect 17644 11852 18052 11880
rect 17644 11840 17650 11852
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 15488 11716 16160 11744
rect 16209 11747 16267 11753
rect 15488 11676 15516 11716
rect 16209 11713 16221 11747
rect 16255 11744 16267 11747
rect 16758 11744 16764 11756
rect 16255 11716 16764 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 17586 11744 17592 11756
rect 17547 11716 17592 11744
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 17770 11704 17776 11756
rect 17828 11744 17834 11756
rect 18325 11747 18383 11753
rect 18325 11744 18337 11747
rect 17828 11716 18337 11744
rect 17828 11704 17834 11716
rect 18325 11713 18337 11716
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 14844 11648 15516 11676
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11676 15623 11679
rect 16482 11676 16488 11688
rect 15611 11648 16488 11676
rect 15611 11645 15623 11648
rect 15565 11639 15623 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 16574 11636 16580 11688
rect 16632 11676 16638 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 16632 11648 18245 11676
rect 16632 11636 16638 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 4154 11608 4160 11620
rect 3160 11580 4160 11608
rect 3053 11571 3111 11577
rect 4154 11568 4160 11580
rect 4212 11568 4218 11620
rect 4249 11611 4307 11617
rect 4249 11577 4261 11611
rect 4295 11608 4307 11611
rect 4338 11608 4344 11620
rect 4295 11580 4344 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 4338 11568 4344 11580
rect 4396 11568 4402 11620
rect 10686 11608 10692 11620
rect 4632 11580 10692 11608
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 1780 11540 1808 11568
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 1780 11512 2329 11540
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2590 11540 2596 11552
rect 2551 11512 2596 11540
rect 2317 11503 2375 11509
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 2866 11540 2872 11552
rect 2827 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 3326 11540 3332 11552
rect 3239 11512 3332 11540
rect 3326 11500 3332 11512
rect 3384 11540 3390 11552
rect 3786 11540 3792 11552
rect 3384 11512 3792 11540
rect 3384 11500 3390 11512
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4632 11549 4660 11580
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 13354 11608 13360 11620
rect 11072 11580 13360 11608
rect 11072 11552 11100 11580
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 15473 11611 15531 11617
rect 14016 11580 14964 11608
rect 14016 11552 14044 11580
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 5074 11540 5080 11552
rect 4856 11512 5080 11540
rect 4856 11500 4862 11512
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5997 11543 6055 11549
rect 5224 11512 5269 11540
rect 5224 11500 5230 11512
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6457 11543 6515 11549
rect 6457 11540 6469 11543
rect 6043 11512 6469 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6457 11509 6469 11512
rect 6503 11509 6515 11543
rect 6457 11503 6515 11509
rect 6917 11543 6975 11549
rect 6917 11509 6929 11543
rect 6963 11540 6975 11543
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 6963 11512 7389 11540
rect 6963 11509 6975 11512
rect 6917 11503 6975 11509
rect 7377 11509 7389 11512
rect 7423 11540 7435 11543
rect 8110 11540 8116 11552
rect 7423 11512 8116 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9030 11540 9036 11552
rect 8352 11512 9036 11540
rect 8352 11500 8358 11512
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9398 11540 9404 11552
rect 9359 11512 9404 11540
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 9640 11512 10333 11540
rect 9640 11500 9646 11512
rect 10321 11509 10333 11512
rect 10367 11540 10379 11543
rect 10962 11540 10968 11552
rect 10367 11512 10968 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11054 11500 11060 11552
rect 11112 11500 11118 11552
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 11238 11540 11244 11552
rect 11195 11512 11244 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11698 11540 11704 11552
rect 11659 11512 11704 11540
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12158 11540 12164 11552
rect 12119 11512 12164 11540
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12492 11512 12537 11540
rect 12492 11500 12498 11512
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12768 11512 12817 11540
rect 12768 11500 12774 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13170 11540 13176 11552
rect 12943 11512 13176 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13265 11543 13323 11549
rect 13265 11509 13277 11543
rect 13311 11540 13323 11543
rect 13446 11540 13452 11552
rect 13311 11512 13452 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13998 11540 14004 11552
rect 13959 11512 14004 11540
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 14274 11540 14280 11552
rect 14235 11512 14280 11540
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14936 11540 14964 11580
rect 15473 11577 15485 11611
rect 15519 11608 15531 11611
rect 15519 11580 17816 11608
rect 15519 11577 15531 11580
rect 15473 11571 15531 11577
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 14936 11512 16313 11540
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 16393 11543 16451 11549
rect 16393 11509 16405 11543
rect 16439 11540 16451 11543
rect 16482 11540 16488 11552
rect 16439 11512 16488 11540
rect 16439 11509 16451 11512
rect 16393 11503 16451 11509
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 16942 11540 16948 11552
rect 16903 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17310 11540 17316 11552
rect 17271 11512 17316 11540
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 17788 11549 17816 11580
rect 17773 11543 17831 11549
rect 17460 11512 17505 11540
rect 17460 11500 17466 11512
rect 17773 11509 17785 11543
rect 17819 11509 17831 11543
rect 18138 11540 18144 11552
rect 18099 11512 18144 11540
rect 17773 11503 17831 11509
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 1578 11296 1584 11348
rect 1636 11336 1642 11348
rect 4062 11336 4068 11348
rect 1636 11308 4068 11336
rect 1636 11296 1642 11308
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 4890 11336 4896 11348
rect 4304 11308 4896 11336
rect 4304 11296 4310 11308
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5224 11308 6009 11336
rect 5224 11296 5230 11308
rect 5997 11305 6009 11308
rect 6043 11305 6055 11339
rect 5997 11299 6055 11305
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 9582 11336 9588 11348
rect 7607 11308 9588 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10468 11308 10885 11336
rect 10468 11296 10474 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 10873 11299 10931 11305
rect 4148 11271 4206 11277
rect 4148 11237 4160 11271
rect 4194 11268 4206 11271
rect 4430 11268 4436 11280
rect 4194 11240 4436 11268
rect 4194 11237 4206 11240
rect 4148 11231 4206 11237
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 5445 11271 5503 11277
rect 5445 11237 5457 11271
rect 5491 11268 5503 11271
rect 5534 11268 5540 11280
rect 5491 11240 5540 11268
rect 5491 11237 5503 11240
rect 5445 11231 5503 11237
rect 5534 11228 5540 11240
rect 5592 11268 5598 11280
rect 5718 11268 5724 11280
rect 5592 11240 5724 11268
rect 5592 11228 5598 11240
rect 5718 11228 5724 11240
rect 5776 11268 5782 11280
rect 5776 11240 8616 11268
rect 5776 11228 5782 11240
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 3418 11160 3424 11212
rect 3476 11209 3482 11212
rect 3476 11200 3488 11209
rect 3476 11172 3521 11200
rect 3476 11163 3488 11172
rect 3476 11160 3482 11163
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 6144 11172 6377 11200
rect 6144 11160 6150 11172
rect 6365 11169 6377 11172
rect 6411 11200 6423 11203
rect 6546 11200 6552 11212
rect 6411 11172 6552 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11200 7251 11203
rect 7650 11200 7656 11212
rect 7239 11172 7656 11200
rect 7239 11169 7251 11172
rect 7193 11163 7251 11169
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11200 8079 11203
rect 8294 11200 8300 11212
rect 8067 11172 8300 11200
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8478 11200 8484 11212
rect 8439 11172 8484 11200
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 8588 11200 8616 11240
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 9370 11271 9428 11277
rect 9370 11268 9382 11271
rect 8904 11240 9382 11268
rect 8904 11228 8910 11240
rect 9370 11237 9382 11240
rect 9416 11237 9428 11271
rect 10686 11268 10692 11280
rect 10647 11240 10692 11268
rect 9370 11231 9428 11237
rect 10686 11228 10692 11240
rect 10744 11228 10750 11280
rect 10888 11268 10916 11299
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11146 11336 11152 11348
rect 11020 11308 11152 11336
rect 11020 11296 11026 11308
rect 11146 11296 11152 11308
rect 11204 11336 11210 11348
rect 11422 11336 11428 11348
rect 11204 11308 11428 11336
rect 11204 11296 11210 11308
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 11517 11339 11575 11345
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 12434 11336 12440 11348
rect 11563 11308 12440 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 13228 11308 13461 11336
rect 13228 11296 13234 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13449 11299 13507 11305
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14090 11336 14096 11348
rect 13955 11308 14096 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 15102 11336 15108 11348
rect 14240 11308 15108 11336
rect 14240 11296 14246 11308
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 16758 11336 16764 11348
rect 16671 11308 16764 11336
rect 16758 11296 16764 11308
rect 16816 11336 16822 11348
rect 16816 11308 17264 11336
rect 16816 11296 16822 11308
rect 10888 11240 11560 11268
rect 11054 11200 11060 11212
rect 8588 11172 10180 11200
rect 11015 11172 11060 11200
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 2314 11132 2320 11144
rect 1811 11104 2320 11132
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 1688 11064 1716 11095
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 3694 11132 3700 11144
rect 3655 11104 3700 11132
rect 3694 11092 3700 11104
rect 3752 11132 3758 11144
rect 3881 11135 3939 11141
rect 3881 11132 3893 11135
rect 3752 11104 3893 11132
rect 3752 11092 3758 11104
rect 3881 11101 3893 11104
rect 3927 11101 3939 11135
rect 3881 11095 3939 11101
rect 5626 11092 5632 11144
rect 5684 11132 5690 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5684 11104 5917 11132
rect 5684 11092 5690 11104
rect 5905 11101 5917 11104
rect 5951 11132 5963 11135
rect 6454 11132 6460 11144
rect 5951 11104 6460 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6638 11132 6644 11144
rect 6599 11104 6644 11132
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7374 11132 7380 11144
rect 7147 11104 7380 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 2222 11064 2228 11076
rect 1688 11036 1808 11064
rect 2183 11036 2228 11064
rect 1780 10996 1808 11036
rect 2222 11024 2228 11036
rect 2280 11024 2286 11076
rect 7024 11064 7052 11095
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11101 7803 11135
rect 7926 11132 7932 11144
rect 7887 11104 7932 11132
rect 7745 11095 7803 11101
rect 7760 11064 7788 11095
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 10152 11132 10180 11172
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11204 11172 11437 11200
rect 11204 11160 11210 11172
rect 11425 11169 11437 11172
rect 11471 11169 11483 11203
rect 11532 11200 11560 11240
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 12526 11268 12532 11280
rect 11940 11240 12532 11268
rect 11940 11228 11946 11240
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 13354 11228 13360 11280
rect 13412 11268 13418 11280
rect 15289 11271 15347 11277
rect 13412 11240 14964 11268
rect 13412 11228 13418 11240
rect 11532 11172 12020 11200
rect 11425 11163 11483 11169
rect 11992 11144 12020 11172
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12233 11203 12291 11209
rect 12233 11200 12245 11203
rect 12124 11172 12245 11200
rect 12124 11160 12130 11172
rect 12233 11169 12245 11172
rect 12279 11169 12291 11203
rect 12233 11163 12291 11169
rect 12618 11160 12624 11212
rect 12676 11200 12682 11212
rect 12676 11172 13216 11200
rect 12676 11160 12682 11172
rect 13188 11144 13216 11172
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 14936 11209 14964 11240
rect 15289 11237 15301 11271
rect 15335 11268 15347 11271
rect 17034 11268 17040 11280
rect 15335 11240 17040 11268
rect 15335 11237 15347 11240
rect 15289 11231 15347 11237
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 17236 11268 17264 11308
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17589 11339 17647 11345
rect 17589 11336 17601 11339
rect 17368 11308 17601 11336
rect 17368 11296 17374 11308
rect 17589 11305 17601 11308
rect 17635 11305 17647 11339
rect 17589 11299 17647 11305
rect 17678 11268 17684 11280
rect 17236 11240 17684 11268
rect 17678 11228 17684 11240
rect 17736 11228 17742 11280
rect 18966 11268 18972 11280
rect 18927 11240 18972 11268
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 13817 11203 13875 11209
rect 13817 11200 13829 11203
rect 13504 11172 13829 11200
rect 13504 11160 13510 11172
rect 13817 11169 13829 11172
rect 13863 11200 13875 11203
rect 14921 11203 14979 11209
rect 13863 11172 14872 11200
rect 13863 11169 13875 11172
rect 13817 11163 13875 11169
rect 11238 11132 11244 11144
rect 10152 11104 11244 11132
rect 9125 11095 9183 11101
rect 7834 11064 7840 11076
rect 7024 11036 7840 11064
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8665 11067 8723 11073
rect 8665 11064 8677 11067
rect 7944 11036 8677 11064
rect 2317 10999 2375 11005
rect 2317 10996 2329 10999
rect 1780 10968 2329 10996
rect 2317 10965 2329 10968
rect 2363 10996 2375 10999
rect 2406 10996 2412 11008
rect 2363 10968 2412 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 4246 10996 4252 11008
rect 2556 10968 4252 10996
rect 2556 10956 2562 10968
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5261 10999 5319 11005
rect 5261 10996 5273 10999
rect 5132 10968 5273 10996
rect 5132 10956 5138 10968
rect 5261 10965 5273 10968
rect 5307 10965 5319 10999
rect 5261 10959 5319 10965
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10996 5687 10999
rect 6178 10996 6184 11008
rect 5675 10968 6184 10996
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 6178 10956 6184 10968
rect 6236 10956 6242 11008
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 7944 10996 7972 11036
rect 8665 11033 8677 11036
rect 8711 11064 8723 11067
rect 9140 11064 9168 11095
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 8711 11036 9168 11064
rect 10505 11067 10563 11073
rect 8711 11033 8723 11036
rect 8665 11027 8723 11033
rect 10505 11033 10517 11067
rect 10551 11064 10563 11067
rect 10686 11064 10692 11076
rect 10551 11036 10692 11064
rect 10551 11033 10563 11036
rect 10505 11027 10563 11033
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 11348 11064 11376 11095
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 11790 11132 11796 11144
rect 11572 11104 11796 11132
rect 11572 11092 11578 11104
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12032 11104 12125 11132
rect 12032 11092 12038 11104
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13630 11132 13636 11144
rect 13228 11104 13636 11132
rect 13228 11092 13234 11104
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 14001 11135 14059 11141
rect 14001 11101 14013 11135
rect 14047 11101 14059 11135
rect 14366 11132 14372 11144
rect 14327 11104 14372 11132
rect 14001 11095 14059 11101
rect 11348 11036 12020 11064
rect 8386 10996 8392 11008
rect 7524 10968 7972 10996
rect 8347 10968 8392 10996
rect 7524 10956 7530 10968
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 8849 10999 8907 11005
rect 8849 10965 8861 10999
rect 8895 10996 8907 10999
rect 9122 10996 9128 11008
rect 8895 10968 9128 10996
rect 8895 10965 8907 10968
rect 8849 10959 8907 10965
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 11882 10996 11888 11008
rect 11843 10968 11888 10996
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 11992 10996 12020 11036
rect 13722 11024 13728 11076
rect 13780 11064 13786 11076
rect 14016 11064 14044 11095
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 13780 11036 14044 11064
rect 13780 11024 13786 11036
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 11992 10968 13369 10996
rect 13357 10965 13369 10968
rect 13403 10996 13415 10999
rect 13538 10996 13544 11008
rect 13403 10968 13544 10996
rect 13403 10965 13415 10968
rect 13357 10959 13415 10965
rect 13538 10956 13544 10968
rect 13596 10956 13602 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14734 10996 14740 11008
rect 13872 10968 14740 10996
rect 13872 10956 13878 10968
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 14844 10996 14872 11172
rect 14921 11169 14933 11203
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 15637 11203 15695 11209
rect 15637 11200 15649 11203
rect 15068 11172 15649 11200
rect 15068 11160 15074 11172
rect 15637 11169 15649 11172
rect 15683 11169 15695 11203
rect 15637 11163 15695 11169
rect 16022 11160 16028 11212
rect 16080 11200 16086 11212
rect 16482 11200 16488 11212
rect 16080 11172 16488 11200
rect 16080 11160 16086 11172
rect 16482 11160 16488 11172
rect 16540 11200 16546 11212
rect 17221 11203 17279 11209
rect 17221 11200 17233 11203
rect 16540 11172 17233 11200
rect 16540 11160 16546 11172
rect 17221 11169 17233 11172
rect 17267 11169 17279 11203
rect 17221 11163 17279 11169
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17405 11163 17463 11169
rect 15102 11092 15108 11144
rect 15160 11132 15166 11144
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 15160 11104 15393 11132
rect 15160 11092 15166 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 16850 11064 16856 11076
rect 16811 11036 16856 11064
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 17420 11064 17448 11163
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 17552 11104 18061 11132
rect 17552 11092 17558 11104
rect 18049 11101 18061 11104
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 18414 11132 18420 11144
rect 18279 11104 18420 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18506 11064 18512 11076
rect 17420 11036 18512 11064
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 16574 10996 16580 11008
rect 14844 10968 16580 10996
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 2225 10795 2283 10801
rect 2225 10792 2237 10795
rect 1912 10764 2237 10792
rect 1912 10752 1918 10764
rect 2225 10761 2237 10764
rect 2271 10761 2283 10795
rect 2225 10755 2283 10761
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 5350 10792 5356 10804
rect 2372 10764 2417 10792
rect 4632 10764 5356 10792
rect 2372 10752 2378 10764
rect 4157 10727 4215 10733
rect 4157 10724 4169 10727
rect 3988 10696 4169 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2961 10659 3019 10665
rect 2961 10656 2973 10659
rect 1719 10628 2973 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2961 10625 2973 10628
rect 3007 10656 3019 10659
rect 3418 10656 3424 10668
rect 3007 10628 3424 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3418 10616 3424 10628
rect 3476 10656 3482 10668
rect 3988 10665 4016 10696
rect 4157 10693 4169 10696
rect 4203 10724 4215 10727
rect 4632 10724 4660 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 7558 10792 7564 10804
rect 5552 10764 7564 10792
rect 4203 10696 4660 10724
rect 4203 10693 4215 10696
rect 4157 10687 4215 10693
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3476 10628 3985 10656
rect 3476 10616 3482 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 5552 10656 5580 10764
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 7834 10792 7840 10804
rect 7795 10764 7840 10792
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 16850 10792 16856 10804
rect 11572 10764 16856 10792
rect 11572 10752 11578 10764
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 18325 10795 18383 10801
rect 18325 10792 18337 10795
rect 17644 10764 18337 10792
rect 17644 10752 17650 10764
rect 18325 10761 18337 10764
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 3973 10619 4031 10625
rect 5460 10628 5580 10656
rect 7852 10656 7880 10752
rect 9309 10727 9367 10733
rect 9309 10693 9321 10727
rect 9355 10693 9367 10727
rect 9309 10687 9367 10693
rect 7852 10628 8064 10656
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2590 10588 2596 10600
rect 1903 10560 2596 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10588 2743 10591
rect 3602 10588 3608 10600
rect 2731 10560 3608 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 3786 10588 3792 10600
rect 3743 10560 3792 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 3786 10548 3792 10560
rect 3844 10588 3850 10600
rect 5460 10588 5488 10628
rect 3844 10560 5488 10588
rect 5537 10591 5595 10597
rect 3844 10548 3850 10560
rect 5537 10557 5549 10591
rect 5583 10588 5595 10591
rect 6362 10588 6368 10600
rect 5583 10560 6368 10588
rect 5583 10557 5595 10560
rect 5537 10551 5595 10557
rect 6362 10548 6368 10560
rect 6420 10588 6426 10600
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 6420 10560 6469 10588
rect 6420 10548 6426 10560
rect 6457 10557 6469 10560
rect 6503 10588 6515 10591
rect 7466 10588 7472 10600
rect 6503 10560 7472 10588
rect 6503 10557 6515 10560
rect 6457 10551 6515 10557
rect 7466 10548 7472 10560
rect 7524 10588 7530 10600
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7524 10560 7941 10588
rect 7524 10548 7530 10560
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 8036 10588 8064 10628
rect 8185 10591 8243 10597
rect 8185 10588 8197 10591
rect 8036 10560 8197 10588
rect 7929 10551 7987 10557
rect 8185 10557 8197 10560
rect 8231 10557 8243 10591
rect 9324 10588 9352 10687
rect 10502 10684 10508 10736
rect 10560 10724 10566 10736
rect 10873 10727 10931 10733
rect 10873 10724 10885 10727
rect 10560 10696 10885 10724
rect 10560 10684 10566 10696
rect 10873 10693 10885 10696
rect 10919 10693 10931 10727
rect 10873 10687 10931 10693
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 11701 10727 11759 10733
rect 11701 10724 11713 10727
rect 11296 10696 11713 10724
rect 11296 10684 11302 10696
rect 11701 10693 11713 10696
rect 11747 10724 11759 10727
rect 12066 10724 12072 10736
rect 11747 10696 12072 10724
rect 11747 10693 11759 10696
rect 11701 10687 11759 10693
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 15010 10724 15016 10736
rect 14875 10696 15016 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 16224 10696 16988 10724
rect 16224 10668 16252 10696
rect 16206 10656 16212 10668
rect 16167 10628 16212 10656
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10656 16451 10659
rect 16482 10656 16488 10668
rect 16439 10628 16488 10656
rect 16439 10625 16451 10628
rect 16393 10619 16451 10625
rect 16482 10616 16488 10628
rect 16540 10656 16546 10668
rect 16960 10665 16988 10696
rect 16945 10659 17003 10665
rect 16540 10628 16712 10656
rect 16540 10616 16546 10628
rect 8185 10551 8243 10557
rect 9232 10560 9352 10588
rect 9401 10591 9459 10597
rect 2792 10492 5028 10520
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 1854 10452 1860 10464
rect 1811 10424 1860 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2792 10461 2820 10492
rect 2777 10455 2835 10461
rect 2777 10452 2789 10455
rect 2188 10424 2789 10452
rect 2188 10412 2194 10424
rect 2777 10421 2789 10424
rect 2823 10421 2835 10455
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 2777 10415 2835 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 5000 10452 5028 10492
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 6730 10529 6736 10532
rect 5270 10523 5328 10529
rect 5270 10520 5282 10523
rect 5132 10492 5282 10520
rect 5132 10480 5138 10492
rect 5270 10489 5282 10492
rect 5316 10489 5328 10523
rect 5813 10523 5871 10529
rect 5813 10520 5825 10523
rect 5270 10483 5328 10489
rect 5644 10492 5825 10520
rect 5644 10452 5672 10492
rect 5813 10489 5825 10492
rect 5859 10520 5871 10523
rect 6089 10523 6147 10529
rect 6089 10520 6101 10523
rect 5859 10492 6101 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6089 10489 6101 10492
rect 6135 10520 6147 10523
rect 6135 10492 6684 10520
rect 6135 10489 6147 10492
rect 6089 10483 6147 10489
rect 3844 10424 3889 10452
rect 5000 10424 5672 10452
rect 5721 10455 5779 10461
rect 3844 10412 3850 10424
rect 5721 10421 5733 10455
rect 5767 10452 5779 10455
rect 5994 10452 6000 10464
rect 5767 10424 6000 10452
rect 5767 10421 5779 10424
rect 5721 10415 5779 10421
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6656 10452 6684 10492
rect 6724 10483 6736 10529
rect 6788 10520 6794 10532
rect 6788 10492 6824 10520
rect 6730 10480 6736 10483
rect 6788 10480 6794 10492
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 9232 10520 9260 10560
rect 9401 10557 9413 10591
rect 9447 10588 9459 10591
rect 10410 10588 10416 10600
rect 9447 10560 10416 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 10410 10548 10416 10560
rect 10468 10588 10474 10600
rect 10962 10588 10968 10600
rect 10468 10560 10968 10588
rect 10468 10548 10474 10560
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11425 10591 11483 10597
rect 11425 10588 11437 10591
rect 11112 10560 11437 10588
rect 11112 10548 11118 10560
rect 11425 10557 11437 10560
rect 11471 10588 11483 10591
rect 11514 10588 11520 10600
rect 11471 10560 11520 10588
rect 11471 10557 11483 10560
rect 11425 10551 11483 10557
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 16684 10597 16712 10628
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 12032 10560 13093 10588
rect 12032 10548 12038 10560
rect 13081 10557 13093 10560
rect 13127 10588 13139 10591
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 13127 10560 13369 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 16669 10591 16727 10597
rect 13357 10551 13415 10557
rect 13464 10560 16528 10588
rect 9674 10529 9680 10532
rect 9646 10523 9680 10529
rect 9646 10520 9658 10523
rect 7800 10492 8708 10520
rect 9232 10492 9658 10520
rect 7800 10480 7806 10492
rect 7834 10452 7840 10464
rect 6656 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10452 7898 10464
rect 8570 10452 8576 10464
rect 7892 10424 8576 10452
rect 7892 10412 7898 10424
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 8680 10452 8708 10492
rect 9646 10489 9658 10492
rect 9732 10520 9738 10532
rect 11149 10523 11207 10529
rect 9732 10492 9794 10520
rect 9646 10483 9680 10489
rect 9674 10480 9680 10483
rect 9732 10480 9738 10492
rect 11149 10489 11161 10523
rect 11195 10520 11207 10523
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 11195 10492 11253 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 11241 10489 11253 10492
rect 11287 10520 11299 10523
rect 11606 10520 11612 10532
rect 11287 10492 11612 10520
rect 11287 10489 11299 10492
rect 11241 10483 11299 10489
rect 11606 10480 11612 10492
rect 11664 10480 11670 10532
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 12814 10523 12872 10529
rect 12814 10520 12826 10523
rect 12676 10492 12826 10520
rect 12676 10480 12682 10492
rect 12814 10489 12826 10492
rect 12860 10489 12872 10523
rect 13464 10520 13492 10560
rect 12814 10483 12872 10489
rect 13096 10492 13492 10520
rect 13096 10452 13124 10492
rect 13538 10480 13544 10532
rect 13596 10529 13602 10532
rect 16500 10529 16528 10560
rect 16669 10557 16681 10591
rect 16715 10557 16727 10591
rect 16669 10551 16727 10557
rect 13596 10523 13660 10529
rect 13596 10489 13614 10523
rect 13648 10489 13660 10523
rect 13596 10483 13660 10489
rect 15953 10523 16011 10529
rect 15953 10489 15965 10523
rect 15999 10520 16011 10523
rect 16485 10523 16543 10529
rect 15999 10489 16022 10520
rect 15953 10483 16022 10489
rect 16485 10489 16497 10523
rect 16531 10489 16543 10523
rect 16485 10483 16543 10489
rect 17212 10523 17270 10529
rect 17212 10489 17224 10523
rect 17258 10520 17270 10523
rect 17770 10520 17776 10532
rect 17258 10492 17776 10520
rect 17258 10489 17270 10492
rect 17212 10483 17270 10489
rect 13596 10480 13602 10483
rect 15994 10464 16022 10483
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 8680 10424 13124 10452
rect 13265 10455 13323 10461
rect 13265 10421 13277 10455
rect 13311 10452 13323 10455
rect 13446 10452 13452 10464
rect 13311 10424 13452 10452
rect 13311 10421 13323 10424
rect 13265 10415 13323 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14734 10452 14740 10464
rect 14695 10424 14740 10452
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 15994 10424 16028 10464
rect 16022 10412 16028 10424
rect 16080 10452 16086 10464
rect 17586 10452 17592 10464
rect 16080 10424 17592 10452
rect 16080 10412 16086 10424
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 18598 10452 18604 10464
rect 18555 10424 18604 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 3326 10248 3332 10260
rect 3287 10220 3332 10248
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3786 10208 3792 10260
rect 3844 10248 3850 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 3844 10220 4445 10248
rect 3844 10208 3850 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4433 10211 4491 10217
rect 4724 10220 4905 10248
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 4724 10180 4752 10220
rect 4893 10217 4905 10220
rect 4939 10248 4951 10251
rect 5994 10248 6000 10260
rect 4939 10220 6000 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6181 10251 6239 10257
rect 6181 10217 6193 10251
rect 6227 10248 6239 10251
rect 6270 10248 6276 10260
rect 6227 10220 6276 10248
rect 6227 10217 6239 10220
rect 6181 10211 6239 10217
rect 6270 10208 6276 10220
rect 6328 10248 6334 10260
rect 6457 10251 6515 10257
rect 6457 10248 6469 10251
rect 6328 10220 6469 10248
rect 6328 10208 6334 10220
rect 6457 10217 6469 10220
rect 6503 10248 6515 10251
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6503 10220 7021 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7374 10248 7380 10260
rect 7335 10220 7380 10248
rect 7009 10211 7067 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7653 10251 7711 10257
rect 7653 10217 7665 10251
rect 7699 10248 7711 10251
rect 7926 10248 7932 10260
rect 7699 10220 7932 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 8444 10220 9505 10248
rect 8444 10208 8450 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 10505 10251 10563 10257
rect 9640 10220 9685 10248
rect 9640 10208 9646 10220
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 10551 10220 10977 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10965 10217 10977 10220
rect 11011 10217 11023 10251
rect 10965 10211 11023 10217
rect 11793 10251 11851 10257
rect 11793 10217 11805 10251
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 2832 10152 4752 10180
rect 4801 10183 4859 10189
rect 2832 10140 2838 10152
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 5166 10180 5172 10192
rect 4847 10152 5172 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 6012 10180 6040 10208
rect 7466 10180 7472 10192
rect 5408 10152 5856 10180
rect 6012 10152 7472 10180
rect 5408 10140 5414 10152
rect 1664 10115 1722 10121
rect 1664 10081 1676 10115
rect 1710 10112 1722 10115
rect 2406 10112 2412 10124
rect 1710 10084 2412 10112
rect 1710 10081 1722 10084
rect 1664 10075 1722 10081
rect 2406 10072 2412 10084
rect 2464 10112 2470 10124
rect 4062 10112 4068 10124
rect 2464 10084 3556 10112
rect 4023 10084 4068 10112
rect 2464 10072 2470 10084
rect 3528 10053 3556 10084
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4338 10112 4344 10124
rect 4299 10084 4344 10112
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 5626 10112 5632 10124
rect 5587 10084 5632 10112
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10013 3571 10047
rect 5074 10044 5080 10056
rect 3513 10007 3571 10013
rect 4080 10016 4384 10044
rect 5035 10016 5080 10044
rect 1412 9908 1440 10007
rect 3436 9976 3464 10007
rect 4080 9976 4108 10016
rect 3436 9948 4108 9976
rect 4154 9936 4160 9988
rect 4212 9976 4218 9988
rect 4356 9976 4384 10016
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5718 10044 5724 10056
rect 5679 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5828 10053 5856 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 8021 10183 8079 10189
rect 8021 10149 8033 10183
rect 8067 10180 8079 10183
rect 8202 10180 8208 10192
rect 8067 10152 8208 10180
rect 8067 10149 8079 10152
rect 8021 10143 8079 10149
rect 8202 10140 8208 10152
rect 8260 10180 8266 10192
rect 8849 10183 8907 10189
rect 8849 10180 8861 10183
rect 8260 10152 8861 10180
rect 8260 10140 8266 10152
rect 8849 10149 8861 10152
rect 8895 10180 8907 10183
rect 10318 10180 10324 10192
rect 8895 10152 10324 10180
rect 8895 10149 8907 10152
rect 8849 10143 8907 10149
rect 9508 10124 9536 10152
rect 10318 10140 10324 10152
rect 10376 10140 10382 10192
rect 10413 10183 10471 10189
rect 10413 10149 10425 10183
rect 10459 10180 10471 10183
rect 11808 10180 11836 10211
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 12768 10220 13185 10248
rect 12768 10208 12774 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 13541 10251 13599 10257
rect 13541 10217 13553 10251
rect 13587 10248 13599 10251
rect 14366 10248 14372 10260
rect 13587 10220 14372 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14921 10251 14979 10257
rect 14921 10217 14933 10251
rect 14967 10248 14979 10251
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14967 10220 15301 10248
rect 14967 10217 14979 10220
rect 14921 10211 14979 10217
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 15289 10211 15347 10217
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 16117 10251 16175 10257
rect 16117 10248 16129 10251
rect 15703 10220 16129 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 16117 10217 16129 10220
rect 16163 10217 16175 10251
rect 16482 10248 16488 10260
rect 16443 10220 16488 10248
rect 16117 10211 16175 10217
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 17402 10248 17408 10260
rect 17363 10220 17408 10248
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 17862 10248 17868 10260
rect 17823 10220 17868 10248
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 10459 10152 11836 10180
rect 10459 10149 10471 10152
rect 10413 10143 10471 10149
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 11940 10152 12940 10180
rect 11940 10140 11946 10152
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7742 10112 7748 10124
rect 7156 10084 7748 10112
rect 7156 10072 7162 10084
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7892 10084 8125 10112
rect 7892 10072 7898 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 9490 10072 9496 10124
rect 9548 10072 9554 10124
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 11333 10115 11391 10121
rect 11333 10112 11345 10115
rect 10560 10084 11345 10112
rect 10560 10072 10566 10084
rect 11333 10081 11345 10084
rect 11379 10112 11391 10115
rect 12066 10112 12072 10124
rect 11379 10084 12072 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10112 12219 10115
rect 12710 10112 12716 10124
rect 12207 10084 12716 10112
rect 12207 10081 12219 10084
rect 12161 10075 12219 10081
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 12912 10121 12940 10152
rect 13446 10140 13452 10192
rect 13504 10180 13510 10192
rect 14829 10183 14887 10189
rect 13504 10152 14228 10180
rect 13504 10140 13510 10152
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 13262 10072 13268 10124
rect 13320 10112 13326 10124
rect 14200 10121 14228 10152
rect 14829 10149 14841 10183
rect 14875 10180 14887 10183
rect 16942 10180 16948 10192
rect 14875 10152 16948 10180
rect 14875 10149 14887 10152
rect 14829 10143 14887 10149
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 18598 10180 18604 10192
rect 17328 10152 18604 10180
rect 17328 10121 17356 10152
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13320 10084 13645 10112
rect 13320 10072 13326 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 14185 10115 14243 10121
rect 14185 10081 14197 10115
rect 14231 10112 14243 10115
rect 17313 10115 17371 10121
rect 14231 10084 16896 10112
rect 14231 10081 14243 10084
rect 14185 10075 14243 10081
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 6730 10044 6736 10056
rect 6643 10016 6736 10044
rect 5813 10007 5871 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 6914 10044 6920 10056
rect 6875 10016 6920 10044
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10013 8355 10047
rect 8662 10044 8668 10056
rect 8623 10016 8668 10044
rect 8297 10007 8355 10013
rect 5261 9979 5319 9985
rect 5261 9976 5273 9979
rect 4212 9948 4257 9976
rect 4356 9948 5273 9976
rect 4212 9936 4218 9948
rect 5261 9945 5273 9948
rect 5307 9945 5319 9979
rect 6748 9976 6776 10004
rect 5261 9939 5319 9945
rect 6012 9948 6592 9976
rect 6748 9948 8156 9976
rect 2314 9908 2320 9920
rect 1412 9880 2320 9908
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2958 9908 2964 9920
rect 2832 9880 2877 9908
rect 2919 9880 2964 9908
rect 2832 9868 2838 9880
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3292 9880 3893 9908
rect 3292 9868 3298 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 6012 9908 6040 9948
rect 5224 9880 6040 9908
rect 6365 9911 6423 9917
rect 5224 9868 5230 9880
rect 6365 9877 6377 9911
rect 6411 9908 6423 9911
rect 6454 9908 6460 9920
rect 6411 9880 6460 9908
rect 6411 9877 6423 9880
rect 6365 9871 6423 9877
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6564 9908 6592 9948
rect 7098 9908 7104 9920
rect 6564 9880 7104 9908
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 7558 9908 7564 9920
rect 7471 9880 7564 9908
rect 7558 9868 7564 9880
rect 7616 9908 7622 9920
rect 8018 9908 8024 9920
rect 7616 9880 8024 9908
rect 7616 9868 7622 9880
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8128 9908 8156 9948
rect 8202 9908 8208 9920
rect 8128 9880 8208 9908
rect 8202 9868 8208 9880
rect 8260 9908 8266 9920
rect 8312 9908 8340 10007
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 11238 10044 11244 10056
rect 10367 10016 11244 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 11422 10044 11428 10056
rect 11383 10016 11428 10044
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10013 11667 10047
rect 12250 10044 12256 10056
rect 12211 10016 12256 10044
rect 11609 10007 11667 10013
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 9766 9976 9772 9988
rect 8444 9948 9772 9976
rect 8444 9936 8450 9948
rect 9766 9936 9772 9948
rect 9824 9976 9830 9988
rect 10045 9979 10103 9985
rect 10045 9976 10057 9979
rect 9824 9948 10057 9976
rect 9824 9936 9830 9948
rect 10045 9945 10057 9948
rect 10091 9976 10103 9979
rect 10502 9976 10508 9988
rect 10091 9948 10508 9976
rect 10091 9945 10103 9948
rect 10045 9939 10103 9945
rect 10502 9936 10508 9948
rect 10560 9976 10566 9988
rect 10778 9976 10784 9988
rect 10560 9948 10784 9976
rect 10560 9936 10566 9948
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 10873 9979 10931 9985
rect 10873 9945 10885 9979
rect 10919 9976 10931 9979
rect 11146 9976 11152 9988
rect 10919 9948 11152 9976
rect 10919 9945 10931 9948
rect 10873 9939 10931 9945
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11624 9976 11652 10007
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12805 10047 12863 10053
rect 12483 10016 12517 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 13280 10044 13308 10072
rect 12851 10016 13308 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 12452 9976 12480 10007
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 15010 10044 15016 10056
rect 13780 10016 13825 10044
rect 14971 10016 15016 10044
rect 13780 10004 13786 10016
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15654 10004 15660 10056
rect 15712 10044 15718 10056
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15712 10016 15761 10044
rect 15712 10004 15718 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16022 10044 16028 10056
rect 15979 10016 16028 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16868 10044 16896 10084
rect 17313 10081 17325 10115
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 17773 10115 17831 10121
rect 17773 10112 17785 10115
rect 17644 10084 17785 10112
rect 17644 10072 17650 10084
rect 17773 10081 17785 10084
rect 17819 10081 17831 10115
rect 18506 10112 18512 10124
rect 18467 10084 18512 10112
rect 17773 10075 17831 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 17862 10044 17868 10056
rect 16868 10016 17868 10044
rect 16761 10007 16819 10013
rect 12618 9976 12624 9988
rect 11624 9948 12624 9976
rect 12618 9936 12624 9948
rect 12676 9976 12682 9988
rect 13740 9976 13768 10004
rect 16592 9976 16620 10007
rect 12676 9948 13768 9976
rect 14384 9948 16620 9976
rect 12676 9936 12682 9948
rect 8260 9880 8340 9908
rect 8260 9868 8266 9880
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 9125 9911 9183 9917
rect 9125 9908 9137 9911
rect 8904 9880 9137 9908
rect 8904 9868 8910 9880
rect 9125 9877 9137 9880
rect 9171 9877 9183 9911
rect 9125 9871 9183 9877
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 12986 9908 12992 9920
rect 11664 9880 12992 9908
rect 11664 9868 11670 9880
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13262 9908 13268 9920
rect 13127 9880 13268 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 13354 9868 13360 9920
rect 13412 9908 13418 9920
rect 14384 9908 14412 9948
rect 13412 9880 14412 9908
rect 14461 9911 14519 9917
rect 13412 9868 13418 9880
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 14642 9908 14648 9920
rect 14507 9880 14648 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 15010 9908 15016 9920
rect 14792 9880 15016 9908
rect 14792 9868 14798 9880
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 16592 9908 16620 9948
rect 16666 9936 16672 9988
rect 16724 9976 16730 9988
rect 16776 9976 16804 10007
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10044 18107 10047
rect 18414 10044 18420 10056
rect 18095 10016 18420 10044
rect 18095 10013 18107 10016
rect 18049 10007 18107 10013
rect 17770 9976 17776 9988
rect 16724 9948 17776 9976
rect 16724 9936 16730 9948
rect 17770 9936 17776 9948
rect 17828 9976 17834 9988
rect 18064 9976 18092 10007
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 17828 9948 18092 9976
rect 17828 9936 17834 9948
rect 17129 9911 17187 9917
rect 17129 9908 17141 9911
rect 16592 9880 17141 9908
rect 17129 9877 17141 9880
rect 17175 9877 17187 9911
rect 17129 9871 17187 9877
rect 17862 9868 17868 9920
rect 17920 9908 17926 9920
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 17920 9880 18337 9908
rect 17920 9868 17926 9880
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 3602 9704 3608 9716
rect 1964 9676 3608 9704
rect 1673 9639 1731 9645
rect 1673 9605 1685 9639
rect 1719 9636 1731 9639
rect 1964 9636 1992 9676
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 3786 9704 3792 9716
rect 3747 9676 3792 9704
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 8386 9704 8392 9716
rect 4396 9676 8392 9704
rect 4396 9664 4402 9676
rect 2774 9636 2780 9648
rect 1719 9608 1992 9636
rect 2056 9608 2780 9636
rect 1719 9605 1731 9608
rect 1673 9599 1731 9605
rect 2056 9577 2084 9608
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 3878 9636 3884 9648
rect 2915 9608 3884 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 3970 9596 3976 9648
rect 4028 9636 4034 9648
rect 5166 9636 5172 9648
rect 4028 9608 5172 9636
rect 4028 9596 4034 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 5261 9639 5319 9645
rect 5261 9605 5273 9639
rect 5307 9605 5319 9639
rect 5261 9599 5319 9605
rect 5353 9639 5411 9645
rect 5353 9605 5365 9639
rect 5399 9636 5411 9639
rect 5534 9636 5540 9648
rect 5399 9608 5540 9636
rect 5399 9605 5411 9608
rect 5353 9599 5411 9605
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9568 2191 9571
rect 2958 9568 2964 9580
rect 2179 9540 2964 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 4341 9571 4399 9577
rect 4341 9568 4353 9571
rect 3712 9540 4353 9568
rect 2222 9500 2228 9512
rect 2183 9472 2228 9500
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3142 9500 3148 9512
rect 3099 9472 3148 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3712 9500 3740 9540
rect 4341 9537 4353 9540
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4982 9568 4988 9580
rect 4755 9540 4988 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5276 9568 5304 9599
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5718 9636 5724 9648
rect 5644 9608 5724 9636
rect 5644 9568 5672 9608
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 6472 9645 6500 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 13446 9704 13452 9716
rect 8628 9676 13452 9704
rect 8628 9664 8634 9676
rect 6457 9639 6515 9645
rect 6457 9605 6469 9639
rect 6503 9605 6515 9639
rect 6457 9599 6515 9605
rect 6825 9639 6883 9645
rect 6825 9605 6837 9639
rect 6871 9636 6883 9639
rect 6914 9636 6920 9648
rect 6871 9608 6920 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 7650 9636 7656 9648
rect 7611 9608 7656 9636
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 8352 9608 8493 9636
rect 8352 9596 8358 9608
rect 8481 9605 8493 9608
rect 8527 9605 8539 9639
rect 8481 9599 8539 9605
rect 5276 9540 5672 9568
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 3970 9500 3976 9512
rect 3436 9472 3740 9500
rect 3931 9472 3976 9500
rect 1489 9435 1547 9441
rect 1489 9401 1501 9435
rect 1535 9432 1547 9435
rect 2866 9432 2872 9444
rect 1535 9404 2872 9432
rect 1535 9401 1547 9404
rect 1489 9395 1547 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3326 9432 3332 9444
rect 3239 9404 3332 9432
rect 3326 9392 3332 9404
rect 3384 9432 3390 9444
rect 3436 9432 3464 9472
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9500 4307 9503
rect 4614 9500 4620 9512
rect 4295 9472 4620 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6012 9500 6040 9531
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 7282 9568 7288 9580
rect 6144 9540 7288 9568
rect 6144 9528 6150 9540
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7834 9568 7840 9580
rect 7515 9540 7840 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8202 9568 8208 9580
rect 8163 9540 8208 9568
rect 8202 9528 8208 9540
rect 8260 9568 8266 9580
rect 9416 9577 9444 9676
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 13722 9704 13728 9716
rect 13683 9676 13728 9704
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 13872 9676 15608 9704
rect 13872 9664 13878 9676
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11241 9639 11299 9645
rect 11241 9636 11253 9639
rect 11112 9608 11253 9636
rect 11112 9596 11118 9608
rect 11241 9605 11253 9608
rect 11287 9605 11299 9639
rect 11241 9599 11299 9605
rect 11517 9639 11575 9645
rect 11517 9605 11529 9639
rect 11563 9636 11575 9639
rect 12066 9636 12072 9648
rect 11563 9608 12072 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 15580 9636 15608 9676
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 16025 9707 16083 9713
rect 16025 9704 16037 9707
rect 15712 9676 16037 9704
rect 15712 9664 15718 9676
rect 16025 9673 16037 9676
rect 16071 9673 16083 9707
rect 16025 9667 16083 9673
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 16448 9676 16620 9704
rect 16448 9664 16454 9676
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 15580 9608 15761 9636
rect 15749 9605 15761 9608
rect 15795 9636 15807 9639
rect 16592 9636 16620 9676
rect 16666 9664 16672 9716
rect 16724 9664 16730 9716
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 17586 9704 17592 9716
rect 17184 9676 17592 9704
rect 17184 9664 17190 9676
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 15795 9608 16620 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8260 9540 9045 9568
rect 8260 9528 8266 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 10962 9568 10968 9580
rect 10923 9540 10968 9568
rect 9401 9531 9459 9537
rect 10962 9528 10968 9540
rect 11020 9568 11026 9580
rect 16684 9577 16712 9664
rect 12345 9571 12403 9577
rect 12345 9568 12357 9571
rect 11020 9540 12357 9568
rect 11020 9528 11026 9540
rect 12345 9537 12357 9540
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 16669 9571 16727 9577
rect 16669 9537 16681 9571
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 6270 9500 6276 9512
rect 5868 9472 5913 9500
rect 6012 9472 6276 9500
rect 5868 9460 5874 9472
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 6638 9500 6644 9512
rect 6599 9472 6644 9500
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 8570 9500 8576 9512
rect 7208 9472 8576 9500
rect 3384 9404 3464 9432
rect 3384 9392 3390 9404
rect 3510 9392 3516 9444
rect 3568 9432 3574 9444
rect 7208 9441 7236 9472
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8720 9472 8861 9500
rect 8720 9460 8726 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9766 9500 9772 9512
rect 8987 9472 9772 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 10686 9460 10692 9512
rect 10744 9509 10750 9512
rect 10744 9500 10756 9509
rect 10744 9472 10789 9500
rect 10744 9463 10756 9472
rect 10744 9460 10750 9463
rect 11790 9460 11796 9512
rect 11848 9500 11854 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11848 9472 11897 9500
rect 11848 9460 11854 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 14185 9503 14243 9509
rect 11885 9463 11943 9469
rect 12406 9472 14136 9500
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 3568 9404 4108 9432
rect 3568 9392 3574 9404
rect 2590 9364 2596 9376
rect 2551 9336 2596 9364
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 3970 9364 3976 9376
rect 3651 9336 3976 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4080 9373 4108 9404
rect 5092 9404 7205 9432
rect 5092 9376 5120 9404
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 8018 9432 8024 9444
rect 7931 9404 8024 9432
rect 7193 9395 7251 9401
rect 8018 9392 8024 9404
rect 8076 9432 8082 9444
rect 12406 9432 12434 9472
rect 12618 9441 12624 9444
rect 12612 9432 12624 9441
rect 8076 9404 12434 9432
rect 12579 9404 12624 9432
rect 8076 9392 8082 9404
rect 12612 9395 12624 9404
rect 12618 9392 12624 9395
rect 12676 9392 12682 9444
rect 13814 9432 13820 9444
rect 13775 9404 13820 9432
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4764 9336 4813 9364
rect 4764 9324 4770 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 4801 9327 4859 9333
rect 4893 9367 4951 9373
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 5074 9364 5080 9376
rect 4939 9336 5080 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5592 9336 5733 9364
rect 5592 9324 5598 9336
rect 5721 9333 5733 9336
rect 5767 9364 5779 9367
rect 5902 9364 5908 9376
rect 5767 9336 5908 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6086 9324 6092 9376
rect 6144 9364 6150 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 6144 9336 6193 9364
rect 6144 9324 6150 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7926 9364 7932 9376
rect 7340 9336 7932 9364
rect 7340 9324 7346 9336
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8113 9367 8171 9373
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 8294 9364 8300 9376
rect 8159 9336 8300 9364
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 9585 9367 9643 9373
rect 9585 9333 9597 9367
rect 9631 9364 9643 9367
rect 9674 9364 9680 9376
rect 9631 9336 9680 9364
rect 9631 9333 9643 9336
rect 9585 9327 9643 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11238 9364 11244 9376
rect 11195 9336 11244 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11664 9336 11713 9364
rect 11664 9324 11670 9336
rect 11701 9333 11713 9336
rect 11747 9333 11759 9367
rect 11701 9327 11759 9333
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11940 9336 12081 9364
rect 11940 9324 11946 9336
rect 12069 9333 12081 9336
rect 12115 9333 12127 9367
rect 12069 9327 12127 9333
rect 12253 9367 12311 9373
rect 12253 9333 12265 9367
rect 12299 9364 12311 9367
rect 12342 9364 12348 9376
rect 12299 9336 12348 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13504 9336 14013 9364
rect 13504 9324 13510 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 14108 9364 14136 9472
rect 14185 9469 14197 9503
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14452 9503 14510 9509
rect 14452 9469 14464 9503
rect 14498 9500 14510 9503
rect 14734 9500 14740 9512
rect 14498 9472 14740 9500
rect 14498 9469 14510 9472
rect 14452 9463 14510 9469
rect 14200 9432 14228 9463
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 16482 9500 16488 9512
rect 15856 9472 16488 9500
rect 15194 9432 15200 9444
rect 14200 9404 15200 9432
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 15856 9441 15884 9472
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 15396 9404 15853 9432
rect 15396 9364 15424 9404
rect 15841 9401 15853 9404
rect 15887 9401 15899 9435
rect 15841 9395 15899 9401
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 16206 9432 16212 9444
rect 16080 9404 16212 9432
rect 16080 9392 16086 9404
rect 16206 9392 16212 9404
rect 16264 9432 16270 9444
rect 16960 9432 16988 9463
rect 16264 9404 16988 9432
rect 17212 9435 17270 9441
rect 16264 9392 16270 9404
rect 17212 9401 17224 9435
rect 17258 9432 17270 9435
rect 17402 9432 17408 9444
rect 17258 9404 17408 9432
rect 17258 9401 17270 9404
rect 17212 9395 17270 9401
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 15562 9364 15568 9376
rect 14108 9336 15424 9364
rect 15523 9336 15568 9364
rect 14001 9327 14059 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 16390 9364 16396 9376
rect 16351 9336 16396 9364
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 16485 9367 16543 9373
rect 16485 9333 16497 9367
rect 16531 9364 16543 9367
rect 17494 9364 17500 9376
rect 16531 9336 17500 9364
rect 16531 9333 16543 9336
rect 16485 9327 16543 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 17828 9336 18337 9364
rect 17828 9324 17834 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18506 9364 18512 9376
rect 18467 9336 18512 9364
rect 18325 9327 18383 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 2774 9160 2780 9172
rect 2746 9120 2780 9160
rect 2832 9120 2838 9172
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9129 3663 9163
rect 3605 9123 3663 9129
rect 2492 9095 2550 9101
rect 2492 9061 2504 9095
rect 2538 9092 2550 9095
rect 2746 9092 2774 9120
rect 3620 9092 3648 9123
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4706 9160 4712 9172
rect 3936 9132 4712 9160
rect 3936 9120 3942 9132
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 6178 9160 6184 9172
rect 5920 9132 6184 9160
rect 3694 9092 3700 9104
rect 2538 9064 2774 9092
rect 3607 9064 3700 9092
rect 2538 9061 2550 9064
rect 2492 9055 2550 9061
rect 3694 9052 3700 9064
rect 3752 9092 3758 9104
rect 4126 9095 4184 9101
rect 4126 9092 4138 9095
rect 3752 9064 4138 9092
rect 3752 9052 3758 9064
rect 4126 9061 4138 9064
rect 4172 9061 4184 9095
rect 4126 9055 4184 9061
rect 4338 9052 4344 9104
rect 4396 9092 4402 9104
rect 5920 9092 5948 9132
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 7282 9160 7288 9172
rect 6411 9132 7288 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 8202 9160 8208 9172
rect 8163 9132 8208 9160
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 8849 9163 8907 9169
rect 8849 9160 8861 9163
rect 8628 9132 8861 9160
rect 8628 9120 8634 9132
rect 8849 9129 8861 9132
rect 8895 9160 8907 9163
rect 9122 9160 9128 9172
rect 8895 9132 9128 9160
rect 8895 9129 8907 9132
rect 8849 9123 8907 9129
rect 9122 9120 9128 9132
rect 9180 9160 9186 9172
rect 9950 9160 9956 9172
rect 9180 9132 9956 9160
rect 9180 9120 9186 9132
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 10873 9163 10931 9169
rect 10873 9129 10885 9163
rect 10919 9160 10931 9163
rect 11238 9160 11244 9172
rect 10919 9132 11244 9160
rect 10919 9129 10931 9132
rect 10873 9123 10931 9129
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11422 9160 11428 9172
rect 11379 9132 11428 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 11701 9163 11759 9169
rect 11701 9160 11713 9163
rect 11572 9132 11713 9160
rect 11572 9120 11578 9132
rect 11701 9129 11713 9132
rect 11747 9160 11759 9163
rect 12066 9160 12072 9172
rect 11747 9132 12072 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 12250 9160 12256 9172
rect 12207 9132 12256 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12526 9160 12532 9172
rect 12487 9132 12532 9160
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12768 9132 13001 9160
rect 12768 9120 12774 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13354 9160 13360 9172
rect 13228 9132 13360 9160
rect 13228 9120 13234 9132
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 13780 9132 15424 9160
rect 13780 9120 13786 9132
rect 4396 9064 5948 9092
rect 5997 9095 6055 9101
rect 4396 9052 4402 9064
rect 5997 9061 6009 9095
rect 6043 9092 6055 9095
rect 8110 9092 8116 9104
rect 6043 9064 8116 9092
rect 6043 9061 6055 9064
rect 5997 9055 6055 9061
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 8478 9052 8484 9104
rect 8536 9092 8542 9104
rect 11146 9092 11152 9104
rect 8536 9064 11152 9092
rect 8536 9052 8542 9064
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 11256 9092 11284 9120
rect 11256 9064 11744 9092
rect 1486 9024 1492 9036
rect 1447 8996 1492 9024
rect 1486 8984 1492 8996
rect 1544 8984 1550 9036
rect 2130 9024 2136 9036
rect 2091 8996 2136 9024
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 2225 9027 2283 9033
rect 2225 8993 2237 9027
rect 2271 9024 2283 9027
rect 2314 9024 2320 9036
rect 2271 8996 2320 9024
rect 2271 8993 2283 8996
rect 2225 8987 2283 8993
rect 2314 8984 2320 8996
rect 2372 9024 2378 9036
rect 2774 9024 2780 9036
rect 2372 8996 2780 9024
rect 2372 8984 2378 8996
rect 2774 8984 2780 8996
rect 2832 9024 2838 9036
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 2832 8996 3893 9024
rect 2832 8984 2838 8996
rect 3881 8993 3893 8996
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 4614 9024 4620 9036
rect 4028 8996 4620 9024
rect 4028 8984 4034 8996
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 4764 8996 5457 9024
rect 4764 8984 4770 8996
rect 5445 8993 5457 8996
rect 5491 9024 5503 9027
rect 5626 9024 5632 9036
rect 5491 8996 5632 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 5626 8984 5632 8996
rect 5684 9024 5690 9036
rect 6086 9024 6092 9036
rect 5684 8996 6092 9024
rect 5684 8984 5690 8996
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6362 8984 6368 9036
rect 6420 9024 6426 9036
rect 6825 9027 6883 9033
rect 6825 9024 6837 9027
rect 6420 8996 6837 9024
rect 6420 8984 6426 8996
rect 6825 8993 6837 8996
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 7092 9027 7150 9033
rect 7092 8993 7104 9027
rect 7138 9024 7150 9027
rect 7834 9024 7840 9036
rect 7138 8996 7840 9024
rect 7138 8993 7150 8996
rect 7092 8987 7150 8993
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 8352 8996 10793 9024
rect 8352 8984 8358 8996
rect 10781 8993 10793 8996
rect 10827 9024 10839 9027
rect 11606 9024 11612 9036
rect 10827 8996 11612 9024
rect 10827 8993 10839 8996
rect 10781 8987 10839 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11716 9024 11744 9064
rect 12342 9052 12348 9104
rect 12400 9092 12406 9104
rect 12621 9095 12679 9101
rect 12621 9092 12633 9095
rect 12400 9064 12633 9092
rect 12400 9052 12406 9064
rect 12621 9061 12633 9064
rect 12667 9092 12679 9095
rect 15396 9092 15424 9132
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 15712 9132 15761 9160
rect 15712 9120 15718 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 17494 9160 17500 9172
rect 17455 9132 17500 9160
rect 15749 9123 15807 9129
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 17862 9160 17868 9172
rect 17644 9132 17868 9160
rect 17644 9120 17650 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18325 9163 18383 9169
rect 18325 9160 18337 9163
rect 18012 9132 18337 9160
rect 18012 9120 18018 9132
rect 18325 9129 18337 9132
rect 18371 9129 18383 9163
rect 18325 9123 18383 9129
rect 16270 9095 16328 9101
rect 16270 9092 16282 9095
rect 12667 9064 15240 9092
rect 15396 9064 16282 9092
rect 12667 9061 12679 9064
rect 12621 9055 12679 9061
rect 11716 8996 12940 9024
rect 5810 8956 5816 8968
rect 5771 8928 5816 8956
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 6270 8956 6276 8968
rect 5951 8928 6276 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 6270 8916 6276 8928
rect 6328 8916 6334 8968
rect 6454 8956 6460 8968
rect 6415 8928 6460 8956
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 7926 8916 7932 8968
rect 7984 8956 7990 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 7984 8928 9413 8956
rect 7984 8916 7990 8928
rect 9401 8925 9413 8928
rect 9447 8956 9459 8959
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9447 8928 10057 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10226 8956 10232 8968
rect 10139 8928 10232 8956
rect 10045 8919 10103 8925
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8888 1823 8891
rect 1811 8860 2268 8888
rect 1811 8857 1823 8860
rect 1765 8851 1823 8857
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2240 8820 2268 8860
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 8665 8891 8723 8897
rect 8665 8888 8677 8891
rect 5500 8860 6868 8888
rect 5500 8848 5506 8860
rect 3326 8820 3332 8832
rect 2240 8792 3332 8820
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 5258 8820 5264 8832
rect 5219 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 6730 8820 6736 8832
rect 6691 8792 6736 8820
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 6840 8820 6868 8860
rect 8220 8860 8677 8888
rect 8220 8820 8248 8860
rect 8665 8857 8677 8860
rect 8711 8857 8723 8891
rect 10060 8888 10088 8919
rect 10226 8916 10232 8928
rect 10284 8956 10290 8968
rect 10965 8959 11023 8965
rect 10284 8928 10732 8956
rect 10284 8916 10290 8928
rect 10704 8900 10732 8928
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 10060 8860 10548 8888
rect 8665 8851 8723 8857
rect 6840 8792 8248 8820
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8478 8820 8484 8832
rect 8352 8792 8397 8820
rect 8439 8792 8484 8820
rect 8352 8780 8358 8792
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 9582 8820 9588 8832
rect 9543 8792 9588 8820
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 10410 8820 10416 8832
rect 10371 8792 10416 8820
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10520 8820 10548 8860
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 10980 8888 11008 8919
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11514 8956 11520 8968
rect 11112 8928 11520 8956
rect 11112 8916 11118 8928
rect 11514 8916 11520 8928
rect 11572 8956 11578 8968
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11572 8928 11805 8956
rect 11572 8916 11578 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12912 8956 12940 8996
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14826 9024 14832 9036
rect 13872 8996 14832 9024
rect 13872 8984 13878 8996
rect 14826 8984 14832 8996
rect 14884 8984 14890 9036
rect 13446 8956 13452 8968
rect 12912 8928 13452 8956
rect 12805 8919 12863 8925
rect 10744 8860 11008 8888
rect 11992 8888 12020 8919
rect 12526 8888 12532 8900
rect 11992 8860 12532 8888
rect 10744 8848 10750 8860
rect 12526 8848 12532 8860
rect 12584 8888 12590 8900
rect 12820 8888 12848 8919
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8925 13599 8959
rect 14918 8956 14924 8968
rect 14879 8928 14924 8956
rect 13541 8919 13599 8925
rect 13556 8888 13584 8919
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 15212 8956 15240 9064
rect 16270 9061 16282 9064
rect 16316 9092 16328 9095
rect 17218 9092 17224 9104
rect 16316 9064 17224 9092
rect 16316 9061 16328 9064
rect 16270 9055 16328 9061
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 9024 15439 9027
rect 15470 9024 15476 9036
rect 15427 8996 15476 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 16022 9024 16028 9036
rect 15983 8996 16028 9024
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 15068 8928 15113 8956
rect 15212 8928 15700 8956
rect 15068 8916 15074 8928
rect 12584 8860 13584 8888
rect 12584 8848 12590 8860
rect 13630 8848 13636 8900
rect 13688 8888 13694 8900
rect 14001 8891 14059 8897
rect 14001 8888 14013 8891
rect 13688 8860 14013 8888
rect 13688 8848 13694 8860
rect 14001 8857 14013 8860
rect 14047 8888 14059 8891
rect 14550 8888 14556 8900
rect 14047 8860 14556 8888
rect 14047 8857 14059 8860
rect 14001 8851 14059 8857
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 12342 8820 12348 8832
rect 10520 8792 12348 8820
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 14090 8820 14096 8832
rect 14051 8792 14096 8820
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 15672 8829 15700 8928
rect 17052 8928 17969 8956
rect 17052 8888 17080 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 18049 8959 18107 8965
rect 18049 8925 18061 8959
rect 18095 8925 18107 8959
rect 18049 8919 18107 8925
rect 17402 8888 17408 8900
rect 16960 8860 17080 8888
rect 17363 8860 17408 8888
rect 16960 8832 16988 8860
rect 17402 8848 17408 8860
rect 17460 8888 17466 8900
rect 18064 8888 18092 8919
rect 17460 8860 18092 8888
rect 17460 8848 17466 8860
rect 14461 8823 14519 8829
rect 14461 8820 14473 8823
rect 14424 8792 14473 8820
rect 14424 8780 14430 8792
rect 14461 8789 14473 8792
rect 14507 8789 14519 8823
rect 14461 8783 14519 8789
rect 15657 8823 15715 8829
rect 15657 8789 15669 8823
rect 15703 8820 15715 8823
rect 16942 8820 16948 8832
rect 15703 8792 16948 8820
rect 15703 8789 15715 8792
rect 15657 8783 15715 8789
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 3050 8616 3056 8628
rect 2188 8588 3056 8616
rect 2188 8576 2194 8588
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6270 8616 6276 8628
rect 6231 8588 6276 8616
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 7834 8616 7840 8628
rect 7795 8588 7840 8616
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 8076 8588 10977 8616
rect 8076 8576 8082 8588
rect 10965 8585 10977 8588
rect 11011 8616 11023 8619
rect 11790 8616 11796 8628
rect 11011 8588 11796 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 17037 8619 17095 8625
rect 12406 8588 16528 8616
rect 3142 8508 3148 8560
rect 3200 8548 3206 8560
rect 3237 8551 3295 8557
rect 3237 8548 3249 8551
rect 3200 8520 3249 8548
rect 3200 8508 3206 8520
rect 3237 8517 3249 8520
rect 3283 8517 3295 8551
rect 3237 8511 3295 8517
rect 3326 8508 3332 8560
rect 3384 8548 3390 8560
rect 4249 8551 4307 8557
rect 3384 8520 3832 8548
rect 3384 8508 3390 8520
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3510 8480 3516 8492
rect 2832 8452 2877 8480
rect 3068 8452 3516 8480
rect 2832 8440 2838 8452
rect 3068 8421 3096 8452
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 3804 8489 3832 8520
rect 4249 8517 4261 8551
rect 4295 8548 4307 8551
rect 4295 8520 4844 8548
rect 4295 8517 4307 8520
rect 4249 8511 4307 8517
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 3878 8480 3884 8492
rect 3835 8452 3884 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 4614 8480 4620 8492
rect 4488 8452 4620 8480
rect 4488 8440 4494 8452
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4816 8489 4844 8520
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 5040 8520 5181 8548
rect 5040 8508 5046 8520
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 5442 8508 5448 8560
rect 5500 8548 5506 8560
rect 5626 8548 5632 8560
rect 5500 8520 5632 8548
rect 5500 8508 5506 8520
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 5736 8548 5764 8576
rect 9674 8548 9680 8560
rect 5736 8520 6500 8548
rect 9587 8520 9680 8548
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 5258 8480 5264 8492
rect 4939 8452 5264 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 2521 8415 2579 8421
rect 2521 8381 2533 8415
rect 2567 8412 2579 8415
rect 3053 8415 3111 8421
rect 2567 8384 3004 8412
rect 2567 8381 2579 8384
rect 2521 8375 2579 8381
rect 2866 8344 2872 8356
rect 2827 8316 2872 8344
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 2976 8344 3004 8384
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 4338 8412 4344 8424
rect 3467 8384 4344 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 4908 8412 4936 8443
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 5902 8480 5908 8492
rect 5767 8452 5908 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 6472 8480 6500 8520
rect 9600 8480 9628 8520
rect 9674 8508 9680 8520
rect 9732 8548 9738 8560
rect 12406 8548 12434 8588
rect 14277 8551 14335 8557
rect 14277 8548 14289 8551
rect 9732 8520 12434 8548
rect 13924 8520 14289 8548
rect 9732 8508 9738 8520
rect 6472 8452 6592 8480
rect 5350 8412 5356 8424
rect 4448 8384 4936 8412
rect 5311 8384 5356 8412
rect 4448 8356 4476 8384
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 6420 8384 6469 8412
rect 6420 8372 6426 8384
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6564 8412 6592 8452
rect 9508 8452 9628 8480
rect 9329 8415 9387 8421
rect 6564 8384 9260 8412
rect 6457 8375 6515 8381
rect 4430 8344 4436 8356
rect 2976 8316 4436 8344
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 4706 8344 4712 8356
rect 4667 8316 4712 8344
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 5684 8316 5917 8344
rect 5684 8304 5690 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 5905 8307 5963 8313
rect 6270 8304 6276 8356
rect 6328 8344 6334 8356
rect 6702 8347 6760 8353
rect 6702 8344 6714 8347
rect 6328 8316 6714 8344
rect 6328 8304 6334 8316
rect 6702 8313 6714 8316
rect 6748 8313 6760 8347
rect 6702 8307 6760 8313
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8344 8171 8347
rect 8478 8344 8484 8356
rect 8159 8316 8484 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 9232 8344 9260 8384
rect 9329 8381 9341 8415
rect 9375 8412 9387 8415
rect 9508 8412 9536 8452
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 11020 8452 12449 8480
rect 11020 8440 11026 8452
rect 12437 8449 12449 8452
rect 12483 8480 12495 8483
rect 12618 8480 12624 8492
rect 12483 8452 12624 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 13722 8480 13728 8492
rect 12851 8452 13728 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 13924 8489 13952 8520
rect 14277 8517 14289 8520
rect 14323 8517 14335 8551
rect 14277 8511 14335 8517
rect 14366 8508 14372 8560
rect 14424 8548 14430 8560
rect 15105 8551 15163 8557
rect 15105 8548 15117 8551
rect 14424 8520 14780 8548
rect 14424 8508 14430 8520
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14458 8480 14464 8492
rect 14139 8452 14464 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14752 8489 14780 8520
rect 14844 8520 15117 8548
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 9375 8384 9536 8412
rect 9585 8415 9643 8421
rect 9375 8381 9387 8384
rect 9329 8375 9387 8381
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9766 8412 9772 8424
rect 9631 8384 9772 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 13538 8412 13544 8424
rect 12943 8384 13544 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8412 13875 8415
rect 14844 8412 14872 8520
rect 15105 8517 15117 8520
rect 15151 8517 15163 8551
rect 15105 8511 15163 8517
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 16390 8548 16396 8560
rect 15979 8520 16396 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8480 14979 8483
rect 15562 8480 15568 8492
rect 14967 8452 15568 8480
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 15562 8440 15568 8452
rect 15620 8480 15626 8492
rect 15657 8483 15715 8489
rect 15657 8480 15669 8483
rect 15620 8452 15669 8480
rect 15620 8440 15626 8452
rect 15657 8449 15669 8452
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 16500 8489 16528 8588
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 18414 8616 18420 8628
rect 17083 8588 18420 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 17313 8551 17371 8557
rect 17313 8517 17325 8551
rect 17359 8548 17371 8551
rect 17359 8520 17816 8548
rect 17359 8517 17371 8520
rect 17313 8511 17371 8517
rect 16485 8483 16543 8489
rect 15804 8452 16344 8480
rect 15804 8440 15810 8452
rect 15470 8412 15476 8424
rect 13863 8384 14872 8412
rect 15431 8384 15476 8412
rect 13863 8381 13875 8384
rect 13817 8375 13875 8381
rect 15470 8372 15476 8384
rect 15528 8412 15534 8424
rect 16206 8412 16212 8424
rect 15528 8384 16212 8412
rect 15528 8372 15534 8384
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 16316 8421 16344 8452
rect 16485 8449 16497 8483
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8412 16359 8415
rect 16942 8412 16948 8424
rect 16347 8384 16948 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17788 8421 17816 8520
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 17773 8415 17831 8421
rect 17773 8381 17785 8415
rect 17819 8381 17831 8415
rect 17773 8375 17831 8381
rect 9677 8347 9735 8353
rect 9232 8316 9536 8344
rect 1397 8279 1455 8285
rect 1397 8245 1409 8279
rect 1443 8276 1455 8279
rect 1670 8276 1676 8288
rect 1443 8248 1676 8276
rect 1443 8245 1455 8248
rect 1397 8239 1455 8245
rect 1670 8236 1676 8248
rect 1728 8236 1734 8288
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 3881 8279 3939 8285
rect 3881 8276 3893 8279
rect 3568 8248 3893 8276
rect 3568 8236 3574 8248
rect 3881 8245 3893 8248
rect 3927 8245 3939 8279
rect 3881 8239 3939 8245
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4341 8279 4399 8285
rect 4341 8276 4353 8279
rect 4212 8248 4353 8276
rect 4212 8236 4218 8248
rect 4341 8245 4353 8248
rect 4387 8245 4399 8279
rect 4341 8239 4399 8245
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 5718 8276 5724 8288
rect 5316 8248 5724 8276
rect 5316 8236 5322 8248
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 5813 8279 5871 8285
rect 5813 8245 5825 8279
rect 5859 8276 5871 8279
rect 6454 8276 6460 8288
rect 5859 8248 6460 8276
rect 5859 8245 5871 8248
rect 5813 8239 5871 8245
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 8205 8279 8263 8285
rect 8205 8245 8217 8279
rect 8251 8276 8263 8279
rect 8662 8276 8668 8288
rect 8251 8248 8668 8276
rect 8251 8245 8263 8248
rect 8205 8239 8263 8245
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9398 8276 9404 8288
rect 9088 8248 9404 8276
rect 9088 8236 9094 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9508 8276 9536 8316
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 10318 8344 10324 8356
rect 9723 8316 10324 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 10318 8304 10324 8316
rect 10376 8304 10382 8356
rect 11514 8304 11520 8356
rect 11572 8344 11578 8356
rect 12066 8344 12072 8356
rect 11572 8316 12072 8344
rect 11572 8304 11578 8316
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 12161 8347 12219 8353
rect 12161 8313 12173 8347
rect 12207 8344 12219 8347
rect 12710 8344 12716 8356
rect 12207 8316 12716 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 16393 8347 16451 8353
rect 16393 8344 16405 8347
rect 14200 8316 16405 8344
rect 11238 8276 11244 8288
rect 9508 8248 11244 8276
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 11790 8276 11796 8288
rect 11751 8248 11796 8276
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12989 8279 13047 8285
rect 12308 8248 12353 8276
rect 12308 8236 12314 8248
rect 12989 8245 13001 8279
rect 13035 8276 13047 8279
rect 13170 8276 13176 8288
rect 13035 8248 13176 8276
rect 13035 8245 13047 8248
rect 12989 8239 13047 8245
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 13354 8276 13360 8288
rect 13315 8248 13360 8276
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13449 8279 13507 8285
rect 13449 8245 13461 8279
rect 13495 8276 13507 8279
rect 13538 8276 13544 8288
rect 13495 8248 13544 8276
rect 13495 8245 13507 8248
rect 13449 8239 13507 8245
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 14200 8276 14228 8316
rect 16393 8313 16405 8316
rect 16439 8313 16451 8347
rect 16393 8307 16451 8313
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 17310 8344 17316 8356
rect 16540 8316 17316 8344
rect 16540 8304 16546 8316
rect 17310 8304 17316 8316
rect 17368 8344 17374 8356
rect 17420 8344 17448 8375
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17920 8384 18061 8412
rect 17920 8372 17926 8384
rect 18049 8381 18061 8384
rect 18095 8412 18107 8415
rect 18138 8412 18144 8424
rect 18095 8384 18144 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 18414 8412 18420 8424
rect 18375 8384 18420 8412
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 17954 8344 17960 8356
rect 17368 8316 17448 8344
rect 17915 8316 17960 8344
rect 17368 8304 17374 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 13688 8248 14228 8276
rect 13688 8236 13694 8248
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 14645 8279 14703 8285
rect 14645 8276 14657 8279
rect 14608 8248 14657 8276
rect 14608 8236 14614 8248
rect 14645 8245 14657 8248
rect 14691 8245 14703 8279
rect 14645 8239 14703 8245
rect 15565 8279 15623 8285
rect 15565 8245 15577 8279
rect 15611 8276 15623 8279
rect 16666 8276 16672 8288
rect 15611 8248 16672 8276
rect 15611 8245 15623 8248
rect 15565 8239 15623 8245
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 17586 8276 17592 8288
rect 17547 8248 17592 8276
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 2087 8044 2605 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 3007 8044 3893 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3881 8041 3893 8044
rect 3927 8041 3939 8075
rect 3881 8035 3939 8041
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 5718 8072 5724 8084
rect 4387 8044 5724 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6270 8072 6276 8084
rect 5868 8044 6276 8072
rect 5868 8032 5874 8044
rect 6270 8032 6276 8044
rect 6328 8032 6334 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8041 6423 8075
rect 6365 8035 6423 8041
rect 1670 7964 1676 8016
rect 1728 8004 1734 8016
rect 3418 8004 3424 8016
rect 1728 7976 3188 8004
rect 3379 7976 3424 8004
rect 1728 7964 1734 7976
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2958 7936 2964 7948
rect 2179 7908 2964 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 1596 7800 1624 7899
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 2314 7868 2320 7880
rect 1995 7840 2320 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 3160 7877 3188 7976
rect 3418 7964 3424 7976
rect 3476 7964 3482 8016
rect 3605 8007 3663 8013
rect 3605 7973 3617 8007
rect 3651 8004 3663 8007
rect 6380 8004 6408 8035
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6696 8044 6837 8072
rect 6696 8032 6702 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 8018 8072 8024 8084
rect 6825 8035 6883 8041
rect 7024 8044 8024 8072
rect 3651 7976 6408 8004
rect 3651 7973 3663 7976
rect 3605 7967 3663 7973
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 4614 7936 4620 7948
rect 4295 7908 4620 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 5160 7939 5218 7945
rect 5160 7905 5172 7939
rect 5206 7936 5218 7939
rect 5902 7936 5908 7948
rect 5206 7908 5908 7936
rect 5206 7905 5218 7908
rect 5160 7899 5218 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 7024 7945 7052 8044
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8478 8072 8484 8084
rect 8343 8044 8484 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 8711 8044 9505 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 10735 8044 12480 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 8386 8004 8392 8016
rect 7208 7976 8392 8004
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 7009 7939 7067 7945
rect 6595 7908 6960 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 4430 7868 4436 7880
rect 4391 7840 4436 7868
rect 3145 7831 3203 7837
rect 3068 7800 3096 7831
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4764 7840 4905 7868
rect 4764 7828 4770 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 4893 7831 4951 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 4154 7800 4160 7812
rect 1596 7772 2774 7800
rect 3068 7772 4160 7800
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 2746 7732 2774 7772
rect 4154 7760 4160 7772
rect 4212 7760 4218 7812
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 6932 7800 6960 7908
rect 7009 7905 7021 7939
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7208 7877 7236 7976
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 9306 8004 9312 8016
rect 8496 7976 9312 8004
rect 7466 7936 7472 7948
rect 7427 7908 7472 7936
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 8036 7908 8217 7936
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 7156 7840 7205 7868
rect 7156 7828 7162 7840
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7374 7868 7380 7880
rect 7335 7840 7380 7868
rect 7193 7831 7251 7837
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 8036 7868 8064 7908
rect 8205 7905 8217 7908
rect 8251 7936 8263 7939
rect 8496 7936 8524 7976
rect 9306 7964 9312 7976
rect 9364 7964 9370 8016
rect 9398 7964 9404 8016
rect 9456 8004 9462 8016
rect 10229 8007 10287 8013
rect 10229 8004 10241 8007
rect 9456 7976 10241 8004
rect 9456 7964 9462 7976
rect 10229 7973 10241 7976
rect 10275 7973 10287 8007
rect 10229 7967 10287 7973
rect 11514 7964 11520 8016
rect 11572 8013 11578 8016
rect 11572 8007 11636 8013
rect 11572 7973 11590 8007
rect 11624 7973 11636 8007
rect 12452 8004 12480 8044
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12713 8075 12771 8081
rect 12713 8072 12725 8075
rect 12584 8044 12725 8072
rect 12584 8032 12590 8044
rect 12713 8041 12725 8044
rect 12759 8041 12771 8075
rect 12713 8035 12771 8041
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 13228 8044 13461 8072
rect 13228 8032 13234 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 16758 8072 16764 8084
rect 16540 8044 16764 8072
rect 16540 8032 16546 8044
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 17218 8072 17224 8084
rect 17179 8044 17224 8072
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 17589 8075 17647 8081
rect 17589 8041 17601 8075
rect 17635 8072 17647 8075
rect 17635 8044 17816 8072
rect 17635 8041 17647 8044
rect 17589 8035 17647 8041
rect 13538 8004 13544 8016
rect 12452 7976 13544 8004
rect 11572 7967 11636 7973
rect 11572 7964 11578 7967
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 14458 7964 14464 8016
rect 14516 8004 14522 8016
rect 17788 8013 17816 8044
rect 16086 8007 16144 8013
rect 16086 8004 16098 8007
rect 14516 7976 16098 8004
rect 14516 7964 14522 7976
rect 16086 7973 16098 7976
rect 16132 7973 16144 8007
rect 16086 7967 16144 7973
rect 17773 8007 17831 8013
rect 17773 7973 17785 8007
rect 17819 7973 17831 8007
rect 17773 7967 17831 7973
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 18417 8007 18475 8013
rect 18417 8004 18429 8007
rect 17920 7976 18429 8004
rect 17920 7964 17926 7976
rect 18417 7973 18429 7976
rect 18463 8004 18475 8007
rect 18598 8004 18604 8016
rect 18463 7976 18604 8004
rect 18463 7973 18475 7976
rect 18417 7967 18475 7973
rect 18598 7964 18604 7976
rect 18656 7964 18662 8016
rect 8251 7908 8524 7936
rect 8757 7939 8815 7945
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 10321 7939 10379 7945
rect 8803 7908 9720 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 7484 7840 8064 7868
rect 8113 7871 8171 7877
rect 7484 7800 7512 7840
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8386 7868 8392 7880
rect 8159 7840 8392 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 9692 7877 9720 7908
rect 10321 7905 10333 7939
rect 10367 7936 10379 7939
rect 11054 7936 11060 7948
rect 10367 7908 11060 7936
rect 10367 7905 10379 7908
rect 10321 7899 10379 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 15194 7936 15200 7948
rect 13863 7908 15200 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 15470 7896 15476 7948
rect 15528 7945 15534 7948
rect 15528 7936 15540 7945
rect 15528 7908 15573 7936
rect 15528 7899 15540 7908
rect 15528 7896 15534 7899
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 15712 7908 15761 7936
rect 15712 7896 15718 7908
rect 15749 7905 15761 7908
rect 15795 7936 15807 7939
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15795 7908 15853 7936
rect 15795 7905 15807 7908
rect 15749 7899 15807 7905
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 17276 7908 17417 7936
rect 17276 7896 17282 7908
rect 17405 7905 17417 7908
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9232 7840 9597 7868
rect 5960 7772 6776 7800
rect 6932 7772 7512 7800
rect 7837 7803 7895 7809
rect 5960 7760 5966 7772
rect 3786 7732 3792 7744
rect 2746 7704 3792 7732
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 4614 7732 4620 7744
rect 4304 7704 4620 7732
rect 4304 7692 4310 7704
rect 4614 7692 4620 7704
rect 4672 7732 4678 7744
rect 4709 7735 4767 7741
rect 4709 7732 4721 7735
rect 4672 7704 4721 7732
rect 4672 7692 4678 7704
rect 4709 7701 4721 7704
rect 4755 7701 4767 7735
rect 6748 7732 6776 7772
rect 7837 7769 7849 7803
rect 7883 7800 7895 7803
rect 9232 7800 9260 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 10134 7868 10140 7880
rect 10095 7840 10140 7868
rect 9677 7831 9735 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10870 7868 10876 7880
rect 10831 7840 10876 7868
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7868 13139 7871
rect 13538 7868 13544 7880
rect 13127 7840 13544 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 7883 7772 9260 7800
rect 7883 7769 7895 7772
rect 7837 7763 7895 7769
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 11146 7800 11152 7812
rect 9824 7772 11152 7800
rect 9824 7760 9830 7772
rect 11146 7760 11152 7772
rect 11204 7800 11210 7812
rect 11348 7800 11376 7831
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13906 7868 13912 7880
rect 13867 7840 13912 7868
rect 13906 7828 13912 7840
rect 13964 7828 13970 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 11204 7772 11376 7800
rect 11204 7760 11210 7772
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 14108 7800 14136 7831
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 12676 7772 13860 7800
rect 14108 7772 14381 7800
rect 12676 7760 12682 7772
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 6748 7704 8769 7732
rect 4709 7695 4767 7701
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 8757 7695 8815 7701
rect 8941 7735 8999 7741
rect 8941 7701 8953 7735
rect 8987 7732 8999 7735
rect 9030 7732 9036 7744
rect 8987 7704 9036 7732
rect 8987 7701 8999 7704
rect 8941 7695 8999 7701
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 11238 7732 11244 7744
rect 9180 7704 9225 7732
rect 11199 7704 11244 7732
rect 9180 7692 9186 7704
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 13265 7735 13323 7741
rect 13265 7701 13277 7735
rect 13311 7732 13323 7735
rect 13446 7732 13452 7744
rect 13311 7704 13452 7732
rect 13311 7701 13323 7704
rect 13265 7695 13323 7701
rect 13446 7692 13452 7704
rect 13504 7732 13510 7744
rect 13722 7732 13728 7744
rect 13504 7704 13728 7732
rect 13504 7692 13510 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 13832 7732 13860 7772
rect 14369 7769 14381 7772
rect 14415 7800 14427 7803
rect 14458 7800 14464 7812
rect 14415 7772 14464 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 17954 7800 17960 7812
rect 17915 7772 17960 7800
rect 17954 7760 17960 7772
rect 18012 7760 18018 7812
rect 15010 7732 15016 7744
rect 13832 7704 15016 7732
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 18138 7732 18144 7744
rect 18099 7704 18144 7732
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 1394 7528 1400 7540
rect 1355 7500 1400 7528
rect 1394 7488 1400 7500
rect 1452 7488 1458 7540
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 2961 7531 3019 7537
rect 2961 7528 2973 7531
rect 2372 7500 2973 7528
rect 2372 7488 2378 7500
rect 2961 7497 2973 7500
rect 3007 7497 3019 7531
rect 3510 7528 3516 7540
rect 3471 7500 3516 7528
rect 2961 7491 3019 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5902 7528 5908 7540
rect 4939 7500 5908 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 6454 7528 6460 7540
rect 6415 7500 6460 7528
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 7466 7528 7472 7540
rect 6788 7500 7472 7528
rect 6788 7488 6794 7500
rect 7466 7488 7472 7500
rect 7524 7528 7530 7540
rect 8754 7528 8760 7540
rect 7524 7500 8760 7528
rect 7524 7488 7530 7500
rect 8754 7488 8760 7500
rect 8812 7528 8818 7540
rect 8812 7500 12112 7528
rect 8812 7488 8818 7500
rect 3050 7460 3056 7472
rect 3011 7432 3056 7460
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 4982 7460 4988 7472
rect 4163 7432 4988 7460
rect 2682 7352 2688 7404
rect 2740 7392 2746 7404
rect 4163 7392 4191 7432
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 8478 7460 8484 7472
rect 6880 7432 8340 7460
rect 8439 7432 8484 7460
rect 6880 7420 6886 7432
rect 2740 7364 4191 7392
rect 4249 7395 4307 7401
rect 2740 7352 2746 7364
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4430 7392 4436 7404
rect 4295 7364 4436 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 6730 7392 6736 7404
rect 6196 7364 6736 7392
rect 1578 7324 1584 7336
rect 1539 7296 1584 7324
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 1837 7327 1895 7333
rect 1837 7324 1849 7327
rect 1728 7296 1849 7324
rect 1728 7284 1734 7296
rect 1837 7293 1849 7296
rect 1883 7324 1895 7327
rect 3510 7324 3516 7336
rect 1883 7296 3516 7324
rect 1883 7293 1895 7296
rect 1837 7287 1895 7293
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 3786 7324 3792 7336
rect 3660 7296 3792 7324
rect 3660 7284 3666 7296
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4062 7324 4068 7336
rect 4023 7296 4068 7324
rect 4062 7284 4068 7296
rect 4120 7324 4126 7336
rect 4522 7324 4528 7336
rect 4120 7296 4528 7324
rect 4120 7284 4126 7296
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 6017 7327 6075 7333
rect 6017 7293 6029 7327
rect 6063 7324 6075 7327
rect 6196 7324 6224 7364
rect 6730 7352 6736 7364
rect 6788 7392 6794 7404
rect 7098 7392 7104 7404
rect 6788 7364 7104 7392
rect 6788 7352 6794 7364
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 7834 7392 7840 7404
rect 7791 7364 7840 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 7975 7364 8248 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 6063 7296 6224 7324
rect 6273 7327 6331 7333
rect 6063 7293 6075 7296
rect 6017 7287 6075 7293
rect 6273 7293 6285 7327
rect 6319 7324 6331 7327
rect 6362 7324 6368 7336
rect 6319 7296 6368 7324
rect 6319 7293 6331 7296
rect 6273 7287 6331 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6638 7284 6644 7336
rect 6696 7324 6702 7336
rect 8105 7327 8163 7333
rect 8105 7324 8117 7327
rect 6696 7296 8117 7324
rect 6696 7284 6702 7296
rect 8105 7293 8117 7296
rect 8151 7293 8163 7327
rect 8105 7287 8163 7293
rect 2498 7216 2504 7268
rect 2556 7256 2562 7268
rect 3234 7256 3240 7268
rect 2556 7228 3096 7256
rect 3195 7228 3240 7256
rect 2556 7216 2562 7228
rect 3068 7188 3096 7228
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 7558 7256 7564 7268
rect 3344 7228 7564 7256
rect 3344 7188 3372 7228
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 8220 7256 8248 7364
rect 7708 7228 7753 7256
rect 8128 7228 8248 7256
rect 8312 7256 8340 7432
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9824 7364 10149 7392
rect 9824 7352 9830 7364
rect 10137 7361 10149 7364
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11664 7364 11897 7392
rect 11664 7352 11670 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 12084 7392 12112 7500
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 12308 7500 12357 7528
rect 12308 7488 12314 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 13173 7531 13231 7537
rect 13173 7528 13185 7531
rect 12768 7500 13185 7528
rect 12768 7488 12774 7500
rect 13173 7497 13185 7500
rect 13219 7497 13231 7531
rect 13173 7491 13231 7497
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 14553 7531 14611 7537
rect 14553 7528 14565 7531
rect 13964 7500 14565 7528
rect 13964 7488 13970 7500
rect 14553 7497 14565 7500
rect 14599 7497 14611 7531
rect 14553 7491 14611 7497
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15381 7531 15439 7537
rect 15381 7528 15393 7531
rect 15252 7500 15393 7528
rect 15252 7488 15258 7500
rect 15381 7497 15393 7500
rect 15427 7497 15439 7531
rect 15381 7491 15439 7497
rect 16761 7531 16819 7537
rect 16761 7497 16773 7531
rect 16807 7528 16819 7531
rect 17126 7528 17132 7540
rect 16807 7500 17132 7528
rect 16807 7497 16819 7500
rect 16761 7491 16819 7497
rect 17126 7488 17132 7500
rect 17184 7488 17190 7540
rect 17310 7528 17316 7540
rect 17271 7500 17316 7528
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 17497 7531 17555 7537
rect 17497 7497 17509 7531
rect 17543 7528 17555 7531
rect 17862 7528 17868 7540
rect 17543 7500 17868 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 12161 7463 12219 7469
rect 12161 7429 12173 7463
rect 12207 7460 12219 7463
rect 12526 7460 12532 7472
rect 12207 7432 12532 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 14369 7463 14427 7469
rect 14369 7460 14381 7463
rect 12636 7432 14381 7460
rect 12636 7392 12664 7432
rect 14369 7429 14381 7432
rect 14415 7429 14427 7463
rect 14369 7423 14427 7429
rect 12084 7364 12664 7392
rect 11885 7355 11943 7361
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12768 7364 13001 7392
rect 12768 7352 12774 7364
rect 12989 7361 13001 7364
rect 13035 7392 13047 7395
rect 13630 7392 13636 7404
rect 13035 7364 13636 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13630 7352 13636 7364
rect 13688 7392 13694 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13688 7364 13737 7392
rect 13688 7352 13694 7364
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 8570 7324 8576 7336
rect 8531 7296 8576 7324
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 8829 7327 8887 7333
rect 8829 7324 8841 7327
rect 8720 7296 8841 7324
rect 8720 7284 8726 7296
rect 8829 7293 8841 7296
rect 8875 7293 8887 7327
rect 8829 7287 8887 7293
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 9364 7296 12817 7324
rect 9364 7284 9370 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 13538 7324 13544 7336
rect 13499 7296 13544 7324
rect 12805 7287 12863 7293
rect 8312 7228 10180 7256
rect 7708 7216 7714 7228
rect 8128 7200 8156 7228
rect 3602 7188 3608 7200
rect 3068 7160 3372 7188
rect 3563 7160 3608 7188
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 3973 7191 4031 7197
rect 3973 7157 3985 7191
rect 4019 7188 4031 7191
rect 4154 7188 4160 7200
rect 4019 7160 4160 7188
rect 4019 7157 4031 7160
rect 3973 7151 4031 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4304 7160 4445 7188
rect 4304 7148 4310 7160
rect 4433 7157 4445 7160
rect 4479 7157 4491 7191
rect 4798 7188 4804 7200
rect 4759 7160 4804 7188
rect 4433 7151 4491 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6144 7160 6837 7188
rect 6144 7148 6150 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 6917 7191 6975 7197
rect 6917 7157 6929 7191
rect 6963 7188 6975 7191
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 6963 7160 7297 7188
rect 6963 7157 6975 7160
rect 6917 7151 6975 7157
rect 7285 7157 7297 7160
rect 7331 7157 7343 7191
rect 7285 7151 7343 7157
rect 8110 7148 8116 7200
rect 8168 7148 8174 7200
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9548 7160 9965 7188
rect 9548 7148 9554 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 10152 7188 10180 7228
rect 10226 7216 10232 7268
rect 10284 7256 10290 7268
rect 10404 7259 10462 7265
rect 10404 7256 10416 7259
rect 10284 7228 10416 7256
rect 10284 7216 10290 7228
rect 10404 7225 10416 7228
rect 10450 7256 10462 7259
rect 10962 7256 10968 7268
rect 10450 7228 10968 7256
rect 10450 7225 10462 7228
rect 10404 7219 10462 7225
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 11296 7228 11836 7256
rect 11296 7216 11302 7228
rect 11330 7188 11336 7200
rect 10152 7160 11336 7188
rect 9953 7151 10011 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11514 7188 11520 7200
rect 11475 7160 11520 7188
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 11808 7197 11836 7228
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12713 7259 12771 7265
rect 12713 7256 12725 7259
rect 12676 7228 12725 7256
rect 12676 7216 12682 7228
rect 12713 7225 12725 7228
rect 12759 7225 12771 7259
rect 12820 7256 12848 7287
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14384 7324 14412 7423
rect 14458 7420 14464 7472
rect 14516 7460 14522 7472
rect 16485 7463 16543 7469
rect 16485 7460 16497 7463
rect 14516 7432 16497 7460
rect 14516 7420 14522 7432
rect 16485 7429 16497 7432
rect 16531 7460 16543 7463
rect 16666 7460 16672 7472
rect 16531 7432 16672 7460
rect 16531 7429 16543 7432
rect 16485 7423 16543 7429
rect 16666 7420 16672 7432
rect 16724 7460 16730 7472
rect 18138 7460 18144 7472
rect 16724 7432 18144 7460
rect 16724 7420 16730 7432
rect 18138 7420 18144 7432
rect 18196 7420 18202 7472
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15470 7392 15476 7404
rect 15243 7364 15476 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15470 7352 15476 7364
rect 15528 7392 15534 7404
rect 15933 7395 15991 7401
rect 15933 7392 15945 7395
rect 15528 7364 15945 7392
rect 15528 7352 15534 7364
rect 15933 7361 15945 7364
rect 15979 7361 15991 7395
rect 15933 7355 15991 7361
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 16632 7364 17141 7392
rect 16632 7352 16638 7364
rect 17129 7361 17141 7364
rect 17175 7392 17187 7395
rect 18506 7392 18512 7404
rect 17175 7364 17632 7392
rect 18467 7364 18512 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 13872 7296 14320 7324
rect 14384 7296 14933 7324
rect 13872 7284 13878 7296
rect 14185 7259 14243 7265
rect 14185 7256 14197 7259
rect 12820 7228 14197 7256
rect 12713 7219 12771 7225
rect 14185 7225 14197 7228
rect 14231 7225 14243 7259
rect 14292 7256 14320 7296
rect 14921 7293 14933 7296
rect 14967 7324 14979 7327
rect 17218 7324 17224 7336
rect 14967 7296 17224 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 17604 7333 17632 7364
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 17589 7327 17647 7333
rect 17589 7293 17601 7327
rect 17635 7293 17647 7327
rect 17862 7324 17868 7336
rect 17823 7296 17868 7324
rect 17589 7287 17647 7293
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 15013 7259 15071 7265
rect 15013 7256 15025 7259
rect 14292 7228 15025 7256
rect 14185 7219 14243 7225
rect 15013 7225 15025 7228
rect 15059 7256 15071 7259
rect 16209 7259 16267 7265
rect 16209 7256 16221 7259
rect 15059 7228 16221 7256
rect 15059 7225 15071 7228
rect 15013 7219 15071 7225
rect 16209 7225 16221 7228
rect 16255 7225 16267 7259
rect 16482 7256 16488 7268
rect 16209 7219 16267 7225
rect 16316 7228 16488 7256
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 13170 7188 13176 7200
rect 11839 7160 13176 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 13538 7188 13544 7200
rect 13320 7160 13544 7188
rect 13320 7148 13326 7160
rect 13538 7148 13544 7160
rect 13596 7188 13602 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13596 7160 13645 7188
rect 13596 7148 13602 7160
rect 13633 7157 13645 7160
rect 13679 7157 13691 7191
rect 14090 7188 14096 7200
rect 14051 7160 14096 7188
rect 13633 7151 13691 7157
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 15746 7188 15752 7200
rect 15707 7160 15752 7188
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16316 7188 16344 7228
rect 16482 7216 16488 7228
rect 16540 7216 16546 7268
rect 18325 7259 18383 7265
rect 18325 7256 18337 7259
rect 17788 7228 18337 7256
rect 17788 7197 17816 7228
rect 18325 7225 18337 7228
rect 18371 7225 18383 7259
rect 18325 7219 18383 7225
rect 15887 7160 16344 7188
rect 17773 7191 17831 7197
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 17773 7157 17785 7191
rect 17819 7157 17831 7191
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 17773 7151 17831 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 1636 6956 1891 6984
rect 1636 6944 1642 6956
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6817 1639 6851
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1581 6811 1639 6817
rect 1596 6780 1624 6811
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 1863 6848 1891 6956
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 2133 6987 2191 6993
rect 2133 6984 2145 6987
rect 2096 6956 2145 6984
rect 2096 6944 2102 6956
rect 2133 6953 2145 6956
rect 2179 6953 2191 6987
rect 2682 6984 2688 6996
rect 2133 6947 2191 6953
rect 2339 6956 2688 6984
rect 1949 6919 2007 6925
rect 1949 6885 1961 6919
rect 1995 6916 2007 6919
rect 2339 6916 2367 6956
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 4246 6984 4252 6996
rect 4207 6956 4252 6984
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 5997 6987 6055 6993
rect 5997 6984 6009 6987
rect 4856 6956 6009 6984
rect 4856 6944 4862 6956
rect 5997 6953 6009 6956
rect 6043 6953 6055 6987
rect 5997 6947 6055 6953
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8849 6987 8907 6993
rect 8849 6984 8861 6987
rect 8444 6956 8861 6984
rect 8444 6944 8450 6956
rect 8849 6953 8861 6956
rect 8895 6953 8907 6987
rect 8849 6947 8907 6953
rect 9493 6987 9551 6993
rect 9493 6953 9505 6987
rect 9539 6984 9551 6987
rect 10410 6984 10416 6996
rect 9539 6956 10416 6984
rect 9539 6953 9551 6956
rect 9493 6947 9551 6953
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 12250 6984 12256 6996
rect 10888 6956 12256 6984
rect 1995 6888 2367 6916
rect 1995 6885 2007 6888
rect 1949 6879 2007 6885
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 2562 6919 2620 6925
rect 2562 6916 2574 6919
rect 2464 6888 2574 6916
rect 2464 6876 2470 6888
rect 2562 6885 2574 6888
rect 2608 6885 2620 6919
rect 4338 6916 4344 6928
rect 4251 6888 4344 6916
rect 2562 6879 2620 6885
rect 4338 6876 4344 6888
rect 4396 6916 4402 6928
rect 4982 6916 4988 6928
rect 4396 6888 4988 6916
rect 4396 6876 4402 6888
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 5169 6919 5227 6925
rect 5169 6885 5181 6919
rect 5215 6916 5227 6919
rect 5442 6916 5448 6928
rect 5215 6888 5448 6916
rect 5215 6885 5227 6888
rect 5169 6879 5227 6885
rect 5442 6876 5448 6888
rect 5500 6916 5506 6928
rect 6454 6916 6460 6928
rect 5500 6888 6460 6916
rect 5500 6876 5506 6888
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 6546 6876 6552 6928
rect 6604 6916 6610 6928
rect 6825 6919 6883 6925
rect 6825 6916 6837 6919
rect 6604 6888 6837 6916
rect 6604 6876 6610 6888
rect 6825 6885 6837 6888
rect 6871 6885 6883 6919
rect 6825 6879 6883 6885
rect 7736 6919 7794 6925
rect 7736 6885 7748 6919
rect 7782 6916 7794 6919
rect 8110 6916 8116 6928
rect 7782 6888 8116 6916
rect 7782 6885 7794 6888
rect 7736 6879 7794 6885
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 10888 6916 10916 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 13538 6944 13544 6996
rect 13596 6984 13602 6996
rect 15381 6987 15439 6993
rect 13596 6956 15056 6984
rect 13596 6944 13602 6956
rect 8536 6888 10916 6916
rect 8536 6876 8542 6888
rect 10962 6876 10968 6928
rect 11020 6876 11026 6928
rect 11422 6916 11428 6928
rect 11383 6888 11428 6916
rect 11422 6876 11428 6888
rect 11480 6876 11486 6928
rect 11698 6916 11704 6928
rect 11659 6888 11704 6916
rect 11698 6876 11704 6888
rect 11756 6916 11762 6928
rect 12161 6919 12219 6925
rect 12161 6916 12173 6919
rect 11756 6888 12173 6916
rect 11756 6876 11762 6888
rect 12161 6885 12173 6888
rect 12207 6916 12219 6919
rect 12618 6916 12624 6928
rect 12207 6888 12624 6916
rect 12207 6885 12219 6888
rect 12161 6879 12219 6885
rect 12618 6876 12624 6888
rect 12676 6876 12682 6928
rect 14737 6919 14795 6925
rect 14737 6916 14749 6919
rect 12820 6888 13124 6916
rect 2038 6848 2044 6860
rect 1863 6820 2044 6848
rect 2038 6808 2044 6820
rect 2096 6848 2102 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 2096 6820 2329 6848
rect 2096 6808 2102 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 3142 6848 3148 6860
rect 2317 6811 2375 6817
rect 2424 6820 3148 6848
rect 2424 6780 2452 6820
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 4430 6808 4436 6860
rect 4488 6848 4494 6860
rect 5074 6848 5080 6860
rect 4488 6820 4568 6848
rect 5035 6820 5080 6848
rect 4488 6808 4494 6820
rect 4540 6789 4568 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 5776 6820 6101 6848
rect 5776 6808 5782 6820
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 6730 6848 6736 6860
rect 6089 6811 6147 6817
rect 6288 6820 6736 6848
rect 6288 6789 6316 6820
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 7024 6820 7481 6848
rect 1596 6752 2452 6780
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 3384 6684 3893 6712
rect 3384 6672 3390 6684
rect 3881 6681 3893 6684
rect 3927 6681 3939 6715
rect 5276 6712 5304 6743
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6917 6783 6975 6789
rect 6917 6780 6929 6783
rect 6696 6752 6929 6780
rect 6696 6740 6702 6752
rect 6917 6749 6929 6752
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 5626 6712 5632 6724
rect 3881 6675 3939 6681
rect 4264 6684 5304 6712
rect 5587 6684 5632 6712
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 3697 6647 3755 6653
rect 3697 6613 3709 6647
rect 3743 6644 3755 6647
rect 4264 6644 4292 6684
rect 5184 6656 5212 6684
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 6822 6672 6828 6724
rect 6880 6712 6886 6724
rect 7024 6712 7052 6820
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 8018 6848 8024 6860
rect 7469 6811 7527 6817
rect 7576 6820 8024 6848
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 7576 6780 7604 6820
rect 8018 6808 8024 6820
rect 8076 6808 8082 6860
rect 9674 6848 9680 6860
rect 9324 6820 9680 6848
rect 9324 6789 9352 6820
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 10980 6848 11008 6876
rect 9876 6820 11008 6848
rect 11077 6851 11135 6857
rect 7423 6752 7604 6780
rect 9309 6783 9367 6789
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9582 6780 9588 6792
rect 9447 6752 9588 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 6880 6684 7052 6712
rect 6880 6672 6886 6684
rect 3743 6616 4292 6644
rect 3743 6613 3755 6616
rect 3697 6607 3755 6613
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4396 6616 4721 6644
rect 4396 6604 4402 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 5166 6604 5172 6656
rect 5224 6604 5230 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6457 6647 6515 6653
rect 6457 6644 6469 6647
rect 5868 6616 6469 6644
rect 5868 6604 5874 6616
rect 6457 6613 6469 6616
rect 6503 6613 6515 6647
rect 7116 6644 7144 6743
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9876 6712 9904 6820
rect 11077 6817 11089 6851
rect 11123 6848 11135 6851
rect 11123 6820 11928 6848
rect 11123 6817 11135 6820
rect 11077 6811 11135 6817
rect 11900 6789 11928 6820
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 8812 6684 9904 6712
rect 9953 6715 10011 6721
rect 8812 6672 8818 6684
rect 9953 6681 9965 6715
rect 9999 6712 10011 6715
rect 10226 6712 10232 6724
rect 9999 6684 10232 6712
rect 9999 6681 10011 6684
rect 9953 6675 10011 6681
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 8478 6644 8484 6656
rect 7116 6616 8484 6644
rect 6457 6607 6515 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 9861 6647 9919 6653
rect 9861 6644 9873 6647
rect 9640 6616 9873 6644
rect 9640 6604 9646 6616
rect 9861 6613 9873 6616
rect 9907 6613 9919 6647
rect 9861 6607 9919 6613
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11348 6644 11376 6743
rect 11900 6712 11928 6743
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 12032 6752 12081 6780
rect 12032 6740 12038 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12710 6780 12716 6792
rect 12069 6743 12127 6749
rect 12176 6752 12716 6780
rect 12176 6712 12204 6752
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 11900 6684 12204 6712
rect 12529 6715 12587 6721
rect 12529 6681 12541 6715
rect 12575 6712 12587 6715
rect 12820 6712 12848 6888
rect 12986 6848 12992 6860
rect 12947 6820 12992 6848
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 13096 6848 13124 6888
rect 13740 6888 14749 6916
rect 13740 6848 13768 6888
rect 14737 6885 14749 6888
rect 14783 6885 14795 6919
rect 14737 6879 14795 6885
rect 13096 6820 13768 6848
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14182 6848 14188 6860
rect 13872 6820 13917 6848
rect 14016 6820 14188 6848
rect 13872 6808 13878 6820
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13909 6783 13967 6789
rect 12943 6752 13492 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 13464 6721 13492 6752
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 14016 6780 14044 6820
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 15028 6848 15056 6956
rect 15381 6953 15393 6987
rect 15427 6984 15439 6987
rect 15746 6984 15752 6996
rect 15427 6956 15752 6984
rect 15427 6953 15439 6956
rect 15381 6947 15439 6953
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 17218 6984 17224 6996
rect 17179 6956 17224 6984
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 17494 6984 17500 6996
rect 17455 6956 17500 6984
rect 17494 6944 17500 6956
rect 17552 6944 17558 6996
rect 17773 6987 17831 6993
rect 17773 6953 17785 6987
rect 17819 6984 17831 6987
rect 17862 6984 17868 6996
rect 17819 6956 17868 6984
rect 17819 6953 17831 6956
rect 17773 6947 17831 6953
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 17957 6919 18015 6925
rect 17957 6885 17969 6919
rect 18003 6916 18015 6919
rect 18046 6916 18052 6928
rect 18003 6888 18052 6916
rect 18003 6885 18015 6888
rect 17957 6879 18015 6885
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 15657 6851 15715 6857
rect 15657 6848 15669 6851
rect 15028 6820 15669 6848
rect 15657 6817 15669 6820
rect 15703 6817 15715 6851
rect 18138 6848 18144 6860
rect 18099 6820 18144 6848
rect 15657 6811 15715 6817
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 18322 6848 18328 6860
rect 18283 6820 18328 6848
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 13955 6752 14044 6780
rect 14093 6783 14151 6789
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 14093 6749 14105 6783
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6749 14887 6783
rect 15010 6780 15016 6792
rect 14971 6752 15016 6780
rect 14829 6743 14887 6749
rect 12575 6684 12848 6712
rect 13449 6715 13507 6721
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 13449 6681 13461 6715
rect 13495 6681 13507 6715
rect 13449 6675 13507 6681
rect 13538 6672 13544 6724
rect 13596 6712 13602 6724
rect 14108 6712 14136 6743
rect 14844 6712 14872 6743
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 13596 6684 14136 6712
rect 14200 6684 14872 6712
rect 13596 6672 13602 6684
rect 11204 6616 11376 6644
rect 13357 6647 13415 6653
rect 11204 6604 11210 6616
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 14200 6644 14228 6684
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 15562 6712 15568 6724
rect 15160 6684 15568 6712
rect 15160 6672 15166 6684
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 15930 6712 15936 6724
rect 15843 6684 15936 6712
rect 15930 6672 15936 6684
rect 15988 6712 15994 6724
rect 16482 6712 16488 6724
rect 15988 6684 16488 6712
rect 15988 6672 15994 6684
rect 16482 6672 16488 6684
rect 16540 6712 16546 6724
rect 17954 6712 17960 6724
rect 16540 6684 17960 6712
rect 16540 6672 16546 6684
rect 17954 6672 17960 6684
rect 18012 6672 18018 6724
rect 18506 6712 18512 6724
rect 18467 6684 18512 6712
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 14366 6644 14372 6656
rect 13403 6616 14228 6644
rect 14327 6616 14372 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 14884 6616 15485 6644
rect 14884 6604 14890 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 16945 6647 17003 6653
rect 16945 6644 16957 6647
rect 16172 6616 16957 6644
rect 16172 6604 16178 6616
rect 16945 6613 16957 6616
rect 16991 6613 17003 6647
rect 16945 6607 17003 6613
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 2593 6443 2651 6449
rect 2593 6409 2605 6443
rect 2639 6440 2651 6443
rect 2958 6440 2964 6452
rect 2639 6412 2820 6440
rect 2919 6412 2964 6440
rect 2639 6409 2651 6412
rect 2593 6403 2651 6409
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6341 2743 6375
rect 2792 6372 2820 6412
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 6380 6412 7941 6440
rect 2866 6372 2872 6384
rect 2792 6344 2872 6372
rect 2685 6335 2743 6341
rect 2700 6304 2728 6335
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 3344 6344 4476 6372
rect 3344 6304 3372 6344
rect 3510 6304 3516 6316
rect 1596 6276 2728 6304
rect 2884 6276 3372 6304
rect 3471 6276 3516 6304
rect 1596 6245 1624 6276
rect 1581 6239 1639 6245
rect 1581 6205 1593 6239
rect 1627 6205 1639 6239
rect 2130 6236 2136 6248
rect 2091 6208 2136 6236
rect 1581 6199 1639 6205
rect 2130 6196 2136 6208
rect 2188 6196 2194 6248
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2682 6236 2688 6248
rect 2455 6208 2688 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 2884 6245 2912 6276
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6205 2927 6239
rect 3326 6236 3332 6248
rect 3287 6208 3332 6236
rect 2869 6199 2927 6205
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3602 6236 3608 6248
rect 3467 6208 3608 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4154 6236 4160 6248
rect 4019 6208 4160 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4448 6236 4476 6344
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6273 5687 6307
rect 5810 6304 5816 6316
rect 5771 6276 5816 6304
rect 5629 6267 5687 6273
rect 4798 6236 4804 6248
rect 4448 6208 4804 6236
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5166 6196 5172 6248
rect 5224 6245 5230 6248
rect 5224 6236 5236 6245
rect 5442 6236 5448 6248
rect 5224 6208 5269 6236
rect 5403 6208 5448 6236
rect 5224 6199 5236 6208
rect 5224 6196 5230 6199
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6168 2007 6171
rect 1995 6140 3832 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 1854 6100 1860 6112
rect 1815 6072 1860 6100
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2406 6100 2412 6112
rect 2363 6072 2412 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 3804 6109 3832 6140
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 5460 6168 5488 6196
rect 4764 6140 5488 6168
rect 4764 6128 4770 6140
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 5644 6168 5672 6267
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6236 5963 6239
rect 6380 6236 6408 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 8444 6412 10088 6440
rect 8444 6400 8450 6412
rect 7837 6375 7895 6381
rect 7837 6341 7849 6375
rect 7883 6372 7895 6375
rect 8110 6372 8116 6384
rect 7883 6344 8116 6372
rect 7883 6341 7895 6344
rect 7837 6335 7895 6341
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 8478 6304 8484 6316
rect 8439 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 5951 6208 6408 6236
rect 6457 6239 6515 6245
rect 5951 6205 5963 6208
rect 5905 6199 5963 6205
rect 6457 6205 6469 6239
rect 6503 6236 6515 6239
rect 6503 6208 6868 6236
rect 6503 6205 6515 6208
rect 6457 6199 6515 6205
rect 6840 6180 6868 6208
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 8352 6208 8769 6236
rect 8352 6196 8358 6208
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6236 9091 6239
rect 9079 6208 9260 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 6702 6171 6760 6177
rect 6702 6168 6714 6171
rect 5592 6140 6714 6168
rect 5592 6128 5598 6140
rect 6702 6137 6714 6140
rect 6748 6137 6760 6171
rect 6702 6131 6760 6137
rect 6822 6128 6828 6180
rect 6880 6128 6886 6180
rect 9122 6168 9128 6180
rect 8312 6140 9128 6168
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6069 3847 6103
rect 3789 6063 3847 6069
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 4028 6072 4077 6100
rect 4028 6060 4034 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 6236 6072 6285 6100
rect 6236 6060 6242 6072
rect 6273 6069 6285 6072
rect 6319 6069 6331 6103
rect 6273 6063 6331 6069
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 7926 6100 7932 6112
rect 6512 6072 7932 6100
rect 6512 6060 6518 6072
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8312 6109 8340 6140
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6069 8355 6103
rect 8297 6063 8355 6069
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 8444 6072 8489 6100
rect 8444 6060 8450 6072
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8628 6072 8953 6100
rect 8628 6060 8634 6072
rect 8941 6069 8953 6072
rect 8987 6100 8999 6103
rect 9232 6100 9260 6208
rect 9300 6171 9358 6177
rect 9300 6137 9312 6171
rect 9346 6168 9358 6171
rect 9490 6168 9496 6180
rect 9346 6140 9496 6168
rect 9346 6137 9358 6140
rect 9300 6131 9358 6137
rect 9490 6128 9496 6140
rect 9548 6128 9554 6180
rect 10060 6168 10088 6412
rect 10152 6412 10517 6440
rect 10152 6384 10180 6412
rect 10505 6409 10517 6412
rect 10551 6440 10563 6443
rect 11054 6440 11060 6452
rect 10551 6412 11060 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11204 6412 11529 6440
rect 11204 6400 11210 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11974 6440 11980 6452
rect 11935 6412 11980 6440
rect 11517 6403 11575 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12805 6443 12863 6449
rect 12805 6409 12817 6443
rect 12851 6440 12863 6443
rect 12986 6440 12992 6452
rect 12851 6412 12992 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13630 6440 13636 6452
rect 13591 6412 13636 6440
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 13740 6412 15148 6440
rect 10134 6332 10140 6384
rect 10192 6332 10198 6384
rect 10413 6375 10471 6381
rect 10413 6341 10425 6375
rect 10459 6372 10471 6375
rect 10594 6372 10600 6384
rect 10459 6344 10600 6372
rect 10459 6341 10471 6344
rect 10413 6335 10471 6341
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 11701 6375 11759 6381
rect 11701 6372 11713 6375
rect 10704 6344 11713 6372
rect 10704 6245 10732 6344
rect 11701 6341 11713 6344
rect 11747 6372 11759 6375
rect 13740 6372 13768 6412
rect 11747 6344 13768 6372
rect 11747 6341 11759 6344
rect 11701 6335 11759 6341
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11514 6304 11520 6316
rect 11011 6276 11520 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12032 6276 12449 6304
rect 12032 6264 12038 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 13357 6307 13415 6313
rect 13357 6304 13369 6307
rect 12667 6276 13369 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 13357 6273 13369 6276
rect 13403 6304 13415 6307
rect 13538 6304 13544 6316
rect 13403 6276 13544 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6205 10747 6239
rect 11054 6236 11060 6248
rect 11015 6208 11060 6236
rect 10689 6199 10747 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11149 6239 11207 6245
rect 11149 6205 11161 6239
rect 11195 6236 11207 6239
rect 11790 6236 11796 6248
rect 11195 6208 11796 6236
rect 11195 6205 11207 6208
rect 11149 6199 11207 6205
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 11940 6208 11985 6236
rect 11940 6196 11946 6208
rect 12158 6196 12164 6248
rect 12216 6236 12222 6248
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12216 6208 13277 6236
rect 12216 6196 12222 6208
rect 10060 6140 12388 6168
rect 12360 6112 12388 6140
rect 8987 6072 9260 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10962 6100 10968 6112
rect 9916 6072 10968 6100
rect 9916 6060 9922 6072
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 12342 6100 12348 6112
rect 12303 6072 12348 6100
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 13004 6100 13032 6208
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13556 6236 13584 6264
rect 14746 6239 14804 6245
rect 14746 6236 14758 6239
rect 13556 6208 14758 6236
rect 13265 6199 13323 6205
rect 14746 6205 14758 6208
rect 14792 6205 14804 6239
rect 14746 6199 14804 6205
rect 14918 6196 14924 6248
rect 14976 6236 14982 6248
rect 15120 6245 15148 6412
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17000 6412 17417 6440
rect 17000 6400 17006 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17405 6403 17463 6409
rect 17773 6443 17831 6449
rect 17773 6409 17785 6443
rect 17819 6440 17831 6443
rect 18322 6440 18328 6452
rect 17819 6412 18328 6440
rect 17819 6409 17831 6412
rect 17773 6403 17831 6409
rect 17420 6304 17448 6403
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 17420 6276 17908 6304
rect 15013 6239 15071 6245
rect 15013 6236 15025 6239
rect 14976 6208 15025 6236
rect 14976 6196 14982 6208
rect 15013 6205 15025 6208
rect 15059 6205 15071 6239
rect 15013 6199 15071 6205
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6205 15163 6239
rect 15105 6199 15163 6205
rect 15194 6196 15200 6248
rect 15252 6236 15258 6248
rect 17880 6245 17908 6276
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 15252 6208 17233 6236
rect 15252 6196 15258 6208
rect 17221 6205 17233 6208
rect 17267 6236 17279 6239
rect 17589 6239 17647 6245
rect 17589 6236 17601 6239
rect 17267 6208 17601 6236
rect 17267 6205 17279 6208
rect 17221 6199 17279 6205
rect 17589 6205 17601 6208
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6205 17923 6239
rect 18414 6236 18420 6248
rect 17865 6199 17923 6205
rect 17972 6208 18420 6236
rect 13170 6168 13176 6180
rect 13083 6140 13176 6168
rect 13170 6128 13176 6140
rect 13228 6168 13234 6180
rect 14458 6168 14464 6180
rect 13228 6140 14464 6168
rect 13228 6128 13234 6140
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 14826 6128 14832 6180
rect 14884 6168 14890 6180
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 14884 6140 15577 6168
rect 14884 6128 14890 6140
rect 15565 6137 15577 6140
rect 15611 6137 15623 6171
rect 17972 6168 18000 6208
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 15565 6131 15623 6137
rect 15672 6140 18000 6168
rect 18325 6171 18383 6177
rect 14550 6100 14556 6112
rect 13004 6072 14556 6100
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 14918 6100 14924 6112
rect 14792 6072 14924 6100
rect 14792 6060 14798 6072
rect 14918 6060 14924 6072
rect 14976 6100 14982 6112
rect 15289 6103 15347 6109
rect 15289 6100 15301 6103
rect 14976 6072 15301 6100
rect 14976 6060 14982 6072
rect 15289 6069 15301 6072
rect 15335 6069 15347 6103
rect 15289 6063 15347 6069
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15672 6100 15700 6140
rect 18325 6137 18337 6171
rect 18371 6137 18383 6171
rect 18506 6168 18512 6180
rect 18467 6140 18512 6168
rect 18325 6131 18383 6137
rect 18046 6100 18052 6112
rect 15528 6072 15700 6100
rect 18007 6072 18052 6100
rect 15528 6060 15534 6072
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18340 6100 18368 6131
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 18414 6100 18420 6112
rect 18340 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 3697 5899 3755 5905
rect 3697 5865 3709 5899
rect 3743 5896 3755 5899
rect 3786 5896 3792 5908
rect 3743 5868 3792 5896
rect 3743 5865 3755 5868
rect 3697 5859 3755 5865
rect 3786 5856 3792 5868
rect 3844 5896 3850 5908
rect 4062 5896 4068 5908
rect 3844 5868 4068 5896
rect 3844 5856 3850 5868
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4338 5896 4344 5908
rect 4299 5868 4344 5896
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 4706 5896 4712 5908
rect 4667 5868 4712 5896
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4948 5868 5089 5896
rect 4948 5856 4954 5868
rect 5077 5865 5089 5868
rect 5123 5896 5135 5899
rect 5258 5896 5264 5908
rect 5123 5868 5264 5896
rect 5123 5865 5135 5868
rect 5077 5859 5135 5865
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6840 5868 7205 5896
rect 1848 5831 1906 5837
rect 1848 5797 1860 5831
rect 1894 5828 1906 5831
rect 3970 5828 3976 5840
rect 1894 5800 3976 5828
rect 1894 5797 1906 5800
rect 1848 5791 1906 5797
rect 3970 5788 3976 5800
rect 4028 5828 4034 5840
rect 6672 5831 6730 5837
rect 4028 5800 4568 5828
rect 4028 5788 4034 5800
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 3053 5763 3111 5769
rect 1535 5732 3004 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 2976 5692 3004 5732
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3234 5760 3240 5772
rect 3099 5732 3240 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3694 5760 3700 5772
rect 3559 5732 3700 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 4141 5732 4261 5760
rect 4141 5692 4169 5732
rect 4249 5729 4261 5732
rect 4295 5760 4307 5763
rect 4338 5760 4344 5772
rect 4295 5732 4344 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 4540 5704 4568 5800
rect 6672 5797 6684 5831
rect 6718 5828 6730 5831
rect 6840 5828 6868 5868
rect 7193 5865 7205 5868
rect 7239 5896 7251 5899
rect 8478 5896 8484 5908
rect 7239 5868 8484 5896
rect 7239 5865 7251 5868
rect 7193 5859 7251 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 9401 5899 9459 5905
rect 9401 5896 9413 5899
rect 8588 5868 9413 5896
rect 6718 5800 6868 5828
rect 6718 5797 6730 5800
rect 6672 5791 6730 5797
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8588 5828 8616 5868
rect 9401 5865 9413 5868
rect 9447 5896 9459 5899
rect 9766 5896 9772 5908
rect 9447 5868 9772 5896
rect 9447 5865 9459 5868
rect 9401 5859 9459 5865
rect 9766 5856 9772 5868
rect 9824 5896 9830 5908
rect 11425 5899 11483 5905
rect 11425 5896 11437 5899
rect 9824 5868 11437 5896
rect 9824 5856 9830 5868
rect 11425 5865 11437 5868
rect 11471 5896 11483 5899
rect 13538 5896 13544 5908
rect 11471 5868 12296 5896
rect 13499 5868 13544 5896
rect 11471 5865 11483 5868
rect 11425 5859 11483 5865
rect 8168 5800 8616 5828
rect 8941 5831 8999 5837
rect 8168 5788 8174 5800
rect 8941 5797 8953 5831
rect 8987 5828 8999 5831
rect 9674 5828 9680 5840
rect 8987 5800 9680 5828
rect 8987 5797 8999 5800
rect 8941 5791 8999 5797
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 11146 5828 11152 5840
rect 10192 5800 11152 5828
rect 10192 5788 10198 5800
rect 11146 5788 11152 5800
rect 11204 5828 11210 5840
rect 11204 5800 12204 5828
rect 11204 5788 11210 5800
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 5169 5763 5227 5769
rect 5169 5760 5181 5763
rect 4948 5732 5181 5760
rect 4948 5720 4954 5732
rect 5169 5729 5181 5732
rect 5215 5760 5227 5763
rect 5626 5760 5632 5772
rect 5215 5732 5632 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 6880 5732 6929 5760
rect 6880 5720 6886 5732
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 6917 5723 6975 5729
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 7466 5760 7472 5772
rect 7147 5732 7472 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 2976 5664 4169 5692
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 4580 5664 5273 5692
rect 4580 5652 4586 5664
rect 5261 5661 5273 5664
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 3329 5627 3387 5633
rect 3329 5624 3341 5627
rect 3108 5596 3341 5624
rect 3108 5584 3114 5596
rect 3329 5593 3341 5596
rect 3375 5593 3387 5627
rect 3329 5587 3387 5593
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 5166 5624 5172 5636
rect 4396 5596 5172 5624
rect 4396 5584 4402 5596
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 6932 5624 6960 5723
rect 7466 5720 7472 5732
rect 7524 5760 7530 5772
rect 7834 5760 7840 5772
rect 7524 5732 7840 5760
rect 7524 5720 7530 5732
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8317 5763 8375 5769
rect 8317 5729 8329 5763
rect 8363 5760 8375 5763
rect 9030 5760 9036 5772
rect 8363 5732 9036 5760
rect 8363 5729 8375 5732
rect 8317 5723 8375 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 9456 5732 9505 5760
rect 9456 5720 9462 5732
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5760 10011 5763
rect 10152 5760 10180 5788
rect 9999 5732 10180 5760
rect 10220 5763 10278 5769
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 10220 5729 10232 5763
rect 10266 5760 10278 5763
rect 10594 5760 10600 5772
rect 10266 5732 10600 5760
rect 10266 5729 10278 5732
rect 10220 5723 10278 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 11330 5760 11336 5772
rect 11112 5732 11336 5760
rect 11112 5720 11118 5732
rect 11330 5720 11336 5732
rect 11388 5760 11394 5772
rect 11793 5763 11851 5769
rect 11793 5760 11805 5763
rect 11388 5732 11805 5760
rect 11388 5720 11394 5732
rect 11793 5729 11805 5732
rect 11839 5760 11851 5763
rect 11974 5760 11980 5772
rect 11839 5732 11980 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12176 5769 12204 5800
rect 12161 5763 12219 5769
rect 12161 5729 12173 5763
rect 12207 5729 12219 5763
rect 12268 5760 12296 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 14274 5896 14280 5908
rect 13872 5868 14280 5896
rect 13872 5856 13878 5868
rect 14274 5856 14280 5868
rect 14332 5896 14338 5908
rect 14826 5896 14832 5908
rect 14332 5868 14832 5896
rect 14332 5856 14338 5868
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 15252 5868 15669 5896
rect 15252 5856 15258 5868
rect 15657 5865 15669 5868
rect 15703 5896 15715 5899
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15703 5868 16129 5896
rect 15703 5865 15715 5868
rect 15657 5859 15715 5865
rect 16117 5865 16129 5868
rect 16163 5896 16175 5899
rect 17310 5896 17316 5908
rect 16163 5868 17316 5896
rect 16163 5865 16175 5868
rect 16117 5859 16175 5865
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 18414 5896 18420 5908
rect 17819 5868 18420 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 12428 5831 12486 5837
rect 12428 5797 12440 5831
rect 12474 5828 12486 5831
rect 12526 5828 12532 5840
rect 12474 5800 12532 5828
rect 12474 5797 12486 5800
rect 12428 5791 12486 5797
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 17405 5831 17463 5837
rect 17405 5828 17417 5831
rect 12676 5800 17417 5828
rect 12676 5788 12682 5800
rect 17405 5797 17417 5800
rect 17451 5828 17463 5831
rect 17451 5800 17908 5828
rect 17451 5797 17463 5800
rect 17405 5791 17463 5797
rect 13998 5760 14004 5772
rect 12268 5732 14004 5760
rect 12161 5723 12219 5729
rect 13998 5720 14004 5732
rect 14056 5720 14062 5772
rect 14090 5720 14096 5772
rect 14148 5760 14154 5772
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14148 5732 14749 5760
rect 14148 5720 14154 5732
rect 14737 5729 14749 5732
rect 14783 5760 14795 5763
rect 14826 5760 14832 5772
rect 14783 5732 14832 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 15562 5760 15568 5772
rect 15523 5732 15568 5760
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 16758 5720 16764 5772
rect 16816 5760 16822 5772
rect 17880 5769 17908 5800
rect 18046 5788 18052 5840
rect 18104 5828 18110 5840
rect 18325 5831 18383 5837
rect 18325 5828 18337 5831
rect 18104 5800 18337 5828
rect 18104 5788 18110 5800
rect 18325 5797 18337 5800
rect 18371 5797 18383 5831
rect 18325 5791 18383 5797
rect 17313 5763 17371 5769
rect 17313 5760 17325 5763
rect 16816 5732 17325 5760
rect 16816 5720 16822 5732
rect 17313 5729 17325 5732
rect 17359 5760 17371 5763
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 17359 5732 17601 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 17589 5729 17601 5732
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 9309 5695 9367 5701
rect 8628 5664 8721 5692
rect 8628 5652 8634 5664
rect 9309 5661 9321 5695
rect 9355 5692 9367 5695
rect 9858 5692 9864 5704
rect 9355 5664 9864 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 14458 5692 14464 5704
rect 13771 5664 14464 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5692 15071 5695
rect 15102 5692 15108 5704
rect 15059 5664 15108 5692
rect 15059 5661 15071 5664
rect 15013 5655 15071 5661
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15749 5695 15807 5701
rect 15749 5661 15761 5695
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 6932 5596 7696 5624
rect 2958 5556 2964 5568
rect 2919 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3234 5556 3240 5568
rect 3195 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3844 5528 3893 5556
rect 3844 5516 3850 5528
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 7668 5556 7696 5596
rect 8588 5556 8616 5652
rect 11609 5627 11667 5633
rect 11609 5624 11621 5627
rect 10888 5596 11621 5624
rect 7668 5528 8616 5556
rect 9861 5559 9919 5565
rect 3881 5519 3939 5525
rect 9861 5525 9873 5559
rect 9907 5556 9919 5559
rect 10318 5556 10324 5568
rect 9907 5528 10324 5556
rect 9907 5525 9919 5528
rect 9861 5519 9919 5525
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 10888 5556 10916 5596
rect 11609 5593 11621 5596
rect 11655 5593 11667 5627
rect 11609 5587 11667 5593
rect 11882 5584 11888 5636
rect 11940 5624 11946 5636
rect 11977 5627 12035 5633
rect 11977 5624 11989 5627
rect 11940 5596 11989 5624
rect 11940 5584 11946 5596
rect 11977 5593 11989 5596
rect 12023 5624 12035 5627
rect 12158 5624 12164 5636
rect 12023 5596 12164 5624
rect 12023 5593 12035 5596
rect 11977 5587 12035 5593
rect 12158 5584 12164 5596
rect 12216 5584 12222 5636
rect 14826 5624 14832 5636
rect 13556 5596 14832 5624
rect 11330 5556 11336 5568
rect 10744 5528 10916 5556
rect 11291 5528 11336 5556
rect 10744 5516 10750 5528
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 13556 5556 13584 5596
rect 14826 5584 14832 5596
rect 14884 5584 14890 5636
rect 15120 5624 15148 5652
rect 15764 5624 15792 5655
rect 18506 5624 18512 5636
rect 15120 5596 15792 5624
rect 18467 5596 18512 5624
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 11756 5528 13584 5556
rect 11756 5516 11762 5528
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 13814 5556 13820 5568
rect 13688 5528 13820 5556
rect 13688 5516 13694 5528
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14090 5556 14096 5568
rect 14051 5528 14096 5556
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 14366 5556 14372 5568
rect 14327 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14458 5516 14464 5568
rect 14516 5556 14522 5568
rect 15197 5559 15255 5565
rect 15197 5556 15209 5559
rect 14516 5528 15209 5556
rect 14516 5516 14522 5528
rect 15197 5525 15209 5528
rect 15243 5525 15255 5559
rect 18046 5556 18052 5568
rect 18007 5528 18052 5556
rect 15197 5519 15255 5525
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 1578 5312 1584 5364
rect 1636 5352 1642 5364
rect 2038 5352 2044 5364
rect 1636 5324 2044 5352
rect 1636 5312 1642 5324
rect 2038 5312 2044 5324
rect 2096 5352 2102 5364
rect 3694 5352 3700 5364
rect 2096 5324 3700 5352
rect 2096 5312 2102 5324
rect 2792 5225 2820 5324
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 5442 5352 5448 5364
rect 5224 5324 5448 5352
rect 5224 5312 5230 5324
rect 5442 5312 5448 5324
rect 5500 5352 5506 5364
rect 6546 5352 6552 5364
rect 5500 5324 6040 5352
rect 6507 5324 6552 5352
rect 5500 5312 5506 5324
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 5905 5287 5963 5293
rect 5905 5284 5917 5287
rect 3660 5256 5917 5284
rect 3660 5244 3666 5256
rect 5905 5253 5917 5256
rect 5951 5253 5963 5287
rect 6012 5284 6040 5324
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 6656 5324 8217 5352
rect 6656 5284 6684 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 8386 5312 8392 5364
rect 8444 5352 8450 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8444 5324 8493 5352
rect 8444 5312 8450 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 9122 5312 9128 5364
rect 9180 5352 9186 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 9180 5324 9321 5352
rect 9180 5312 9186 5324
rect 9309 5321 9321 5324
rect 9355 5321 9367 5355
rect 9309 5315 9367 5321
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10137 5355 10195 5361
rect 10137 5352 10149 5355
rect 9824 5324 10149 5352
rect 9824 5312 9830 5324
rect 10137 5321 10149 5324
rect 10183 5321 10195 5355
rect 16574 5352 16580 5364
rect 10137 5315 10195 5321
rect 10244 5324 16580 5352
rect 7650 5284 7656 5296
rect 6012 5256 6684 5284
rect 7208 5256 7656 5284
rect 5905 5247 5963 5253
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 3510 5216 3516 5228
rect 3016 5188 3516 5216
rect 3016 5176 3022 5188
rect 3510 5176 3516 5188
rect 3568 5216 3574 5228
rect 3697 5219 3755 5225
rect 3697 5216 3709 5219
rect 3568 5188 3709 5216
rect 3568 5176 3574 5188
rect 3697 5185 3709 5188
rect 3743 5185 3755 5219
rect 4430 5216 4436 5228
rect 4391 5188 4436 5216
rect 3697 5179 3755 5185
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 7208 5225 7236 5256
rect 7650 5244 7656 5256
rect 7708 5284 7714 5296
rect 7708 5256 9168 5284
rect 7708 5244 7714 5256
rect 9140 5228 9168 5256
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 10244 5284 10272 5324
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 9272 5256 10272 5284
rect 14093 5287 14151 5293
rect 9272 5244 9278 5256
rect 14093 5253 14105 5287
rect 14139 5253 14151 5287
rect 14093 5247 14151 5253
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4663 5188 5365 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 5353 5179 5411 5185
rect 5828 5188 6193 5216
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3142 5148 3148 5160
rect 3099 5120 3148 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 3786 5148 3792 5160
rect 3651 5120 3792 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4304 5120 4353 5148
rect 4304 5108 4310 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 4632 5148 4660 5179
rect 4580 5120 4660 5148
rect 4580 5108 4586 5120
rect 5258 5108 5264 5160
rect 5316 5148 5322 5160
rect 5828 5148 5856 5188
rect 6181 5185 6193 5188
rect 6227 5185 6239 5219
rect 6181 5179 6239 5185
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 8018 5216 8024 5228
rect 7979 5188 8024 5216
rect 7193 5179 7251 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8220 5188 8524 5216
rect 5316 5120 5856 5148
rect 5316 5108 5322 5120
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 5960 5120 6101 5148
rect 5960 5108 5966 5120
rect 6089 5117 6101 5120
rect 6135 5117 6147 5151
rect 6089 5111 6147 5117
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 8220 5148 8248 5188
rect 6963 5120 8248 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 8352 5120 8401 5148
rect 8352 5108 8358 5120
rect 8389 5117 8401 5120
rect 8435 5117 8447 5151
rect 8496 5148 8524 5188
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 8754 5216 8760 5228
rect 8628 5188 8760 5216
rect 8628 5176 8634 5188
rect 8754 5176 8760 5188
rect 8812 5216 8818 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8812 5188 8953 5216
rect 8812 5176 8818 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 8941 5179 8999 5185
rect 9122 5176 9128 5188
rect 9180 5216 9186 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9180 5188 9873 5216
rect 9180 5176 9186 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 9861 5179 9919 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 13814 5216 13820 5228
rect 13004 5188 13820 5216
rect 9214 5148 9220 5160
rect 8496 5120 9220 5148
rect 8389 5111 8447 5117
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9674 5148 9680 5160
rect 9635 5120 9680 5148
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5148 10839 5151
rect 10870 5148 10876 5160
rect 10827 5120 10876 5148
rect 10827 5117 10839 5120
rect 10781 5111 10839 5117
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 12825 5151 12883 5157
rect 12825 5117 12837 5151
rect 12871 5148 12883 5151
rect 13004 5148 13032 5188
rect 13814 5176 13820 5188
rect 13872 5216 13878 5228
rect 14108 5216 14136 5247
rect 16206 5244 16212 5296
rect 16264 5284 16270 5296
rect 17681 5287 17739 5293
rect 17681 5284 17693 5287
rect 16264 5256 17693 5284
rect 16264 5244 16270 5256
rect 17681 5253 17693 5256
rect 17727 5253 17739 5287
rect 17681 5247 17739 5253
rect 15562 5216 15568 5228
rect 13872 5188 14136 5216
rect 15523 5188 15568 5216
rect 13872 5176 13878 5188
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16482 5216 16488 5228
rect 15979 5188 16488 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 12871 5120 13032 5148
rect 13081 5151 13139 5157
rect 12871 5117 12883 5120
rect 12825 5111 12883 5117
rect 13081 5117 13093 5151
rect 13127 5148 13139 5151
rect 13725 5151 13783 5157
rect 13127 5120 13584 5148
rect 13127 5117 13139 5120
rect 13081 5111 13139 5117
rect 2532 5083 2590 5089
rect 2532 5049 2544 5083
rect 2578 5080 2590 5083
rect 2958 5080 2964 5092
rect 2578 5052 2964 5080
rect 2578 5049 2590 5052
rect 2532 5043 2590 5049
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 4706 5080 4712 5092
rect 3559 5052 4712 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5169 5083 5227 5089
rect 5169 5049 5181 5083
rect 5215 5080 5227 5083
rect 5629 5083 5687 5089
rect 5629 5080 5641 5083
rect 5215 5052 5641 5080
rect 5215 5049 5227 5052
rect 5169 5043 5227 5049
rect 5629 5049 5641 5052
rect 5675 5049 5687 5083
rect 9769 5083 9827 5089
rect 9769 5080 9781 5083
rect 5629 5043 5687 5049
rect 6104 5052 9781 5080
rect 1397 5015 1455 5021
rect 1397 4981 1409 5015
rect 1443 5012 1455 5015
rect 2222 5012 2228 5024
rect 1443 4984 2228 5012
rect 1443 4981 1455 4984
rect 1397 4975 1455 4981
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 2832 4984 2881 5012
rect 2832 4972 2838 4984
rect 2869 4981 2881 4984
rect 2915 4981 2927 5015
rect 3142 5012 3148 5024
rect 3103 4984 3148 5012
rect 2869 4975 2927 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 3973 5015 4031 5021
rect 3973 4981 3985 5015
rect 4019 5012 4031 5015
rect 4062 5012 4068 5024
rect 4019 4984 4068 5012
rect 4019 4981 4031 4984
rect 3973 4975 4031 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4798 5012 4804 5024
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5350 5012 5356 5024
rect 5307 4984 5356 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5350 4972 5356 4984
rect 5408 5012 5414 5024
rect 6104 5012 6132 5052
rect 9769 5049 9781 5052
rect 9815 5080 9827 5083
rect 11241 5083 11299 5089
rect 11241 5080 11253 5083
rect 9815 5052 11253 5080
rect 9815 5049 9827 5052
rect 9769 5043 9827 5049
rect 11241 5049 11253 5052
rect 11287 5080 11299 5083
rect 11425 5083 11483 5089
rect 11425 5080 11437 5083
rect 11287 5052 11437 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 11425 5049 11437 5052
rect 11471 5080 11483 5083
rect 13446 5080 13452 5092
rect 11471 5052 13452 5080
rect 11471 5049 11483 5052
rect 11425 5043 11483 5049
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 5408 4984 6132 5012
rect 7009 5015 7067 5021
rect 5408 4972 5414 4984
rect 7009 4981 7021 5015
rect 7055 5012 7067 5015
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 7055 4984 7389 5012
rect 7055 4981 7067 4984
rect 7009 4975 7067 4981
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 7742 5012 7748 5024
rect 7703 4984 7748 5012
rect 7377 4975 7435 4981
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8110 5012 8116 5024
rect 7892 4984 8116 5012
rect 7892 4972 7898 4984
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 8352 4984 8861 5012
rect 8352 4972 8358 4984
rect 8849 4981 8861 4984
rect 8895 5012 8907 5015
rect 9030 5012 9036 5024
rect 8895 4984 9036 5012
rect 8895 4981 8907 4984
rect 8849 4975 8907 4981
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 10410 5012 10416 5024
rect 10371 4984 10416 5012
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 10686 5012 10692 5024
rect 10560 4984 10692 5012
rect 10560 4972 10566 4984
rect 10686 4972 10692 4984
rect 10744 5012 10750 5024
rect 10873 5015 10931 5021
rect 10873 5012 10885 5015
rect 10744 4984 10885 5012
rect 10744 4972 10750 4984
rect 10873 4981 10885 4984
rect 10919 4981 10931 5015
rect 10873 4975 10931 4981
rect 11701 5015 11759 5021
rect 11701 4981 11713 5015
rect 11747 5012 11759 5015
rect 12342 5012 12348 5024
rect 11747 4984 12348 5012
rect 11747 4981 11759 4984
rect 11701 4975 11759 4981
rect 12342 4972 12348 4984
rect 12400 5012 12406 5024
rect 12526 5012 12532 5024
rect 12400 4984 12532 5012
rect 12400 4972 12406 4984
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 12676 4984 13277 5012
rect 12676 4972 12682 4984
rect 13265 4981 13277 4984
rect 13311 4981 13323 5015
rect 13556 5012 13584 5120
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 14366 5148 14372 5160
rect 13771 5120 14372 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 15028 5120 15485 5148
rect 13633 5083 13691 5089
rect 13633 5049 13645 5083
rect 13679 5080 13691 5083
rect 14458 5080 14464 5092
rect 13679 5052 14464 5080
rect 13679 5049 13691 5052
rect 13633 5043 13691 5049
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 14366 5012 14372 5024
rect 13556 4984 14372 5012
rect 13265 4975 13323 4981
rect 14366 4972 14372 4984
rect 14424 5012 14430 5024
rect 14734 5012 14740 5024
rect 14424 4984 14740 5012
rect 14424 4972 14430 4984
rect 14734 4972 14740 4984
rect 14792 5012 14798 5024
rect 15028 5012 15056 5120
rect 15473 5117 15485 5120
rect 15519 5117 15531 5151
rect 17696 5148 17724 5247
rect 18506 5216 18512 5228
rect 18467 5188 18512 5216
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 17865 5151 17923 5157
rect 17865 5148 17877 5151
rect 17696 5120 17877 5148
rect 15473 5111 15531 5117
rect 17865 5117 17877 5120
rect 17911 5117 17923 5151
rect 17865 5111 17923 5117
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18325 5151 18383 5157
rect 18325 5148 18337 5151
rect 18104 5120 18337 5148
rect 18104 5108 18110 5120
rect 18325 5117 18337 5120
rect 18371 5117 18383 5151
rect 18325 5111 18383 5117
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 15206 5083 15264 5089
rect 15206 5080 15218 5083
rect 15160 5052 15218 5080
rect 15160 5040 15166 5052
rect 15206 5049 15218 5052
rect 15252 5049 15264 5083
rect 15206 5043 15264 5049
rect 18046 5012 18052 5024
rect 14792 4984 15056 5012
rect 18007 4984 18052 5012
rect 14792 4972 14798 4984
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1854 4808 1860 4820
rect 1815 4780 1860 4808
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2501 4811 2559 4817
rect 2501 4777 2513 4811
rect 2547 4808 2559 4811
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2547 4780 2973 4808
rect 2547 4777 2559 4780
rect 2501 4771 2559 4777
rect 2961 4777 2973 4780
rect 3007 4777 3019 4811
rect 2961 4771 3019 4777
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 4062 4808 4068 4820
rect 3467 4780 4068 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 7101 4811 7159 4817
rect 4304 4780 6592 4808
rect 4304 4768 4310 4780
rect 1394 4740 1400 4752
rect 1355 4712 1400 4740
rect 1394 4700 1400 4712
rect 1452 4700 1458 4752
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 2409 4743 2467 4749
rect 1627 4712 2176 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 1946 4672 1952 4684
rect 1907 4644 1952 4672
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2148 4672 2176 4712
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 3142 4740 3148 4752
rect 2455 4712 3148 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 4798 4740 4804 4752
rect 3375 4712 4804 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 5074 4700 5080 4752
rect 5132 4740 5138 4752
rect 6564 4740 6592 4780
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 7147 4780 7481 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 7469 4777 7481 4780
rect 7515 4777 7527 4811
rect 7469 4771 7527 4777
rect 8110 4768 8116 4820
rect 8168 4808 8174 4820
rect 9217 4811 9275 4817
rect 8168 4780 8800 4808
rect 8168 4768 8174 4780
rect 6822 4740 6828 4752
rect 5132 4712 6500 4740
rect 6564 4712 6828 4740
rect 5132 4700 5138 4712
rect 3050 4672 3056 4684
rect 2148 4644 3056 4672
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3878 4672 3884 4684
rect 3839 4644 3884 4672
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 4148 4675 4206 4681
rect 4148 4641 4160 4675
rect 4194 4672 4206 4675
rect 5718 4672 5724 4684
rect 4194 4644 5304 4672
rect 5679 4644 5724 4672
rect 4194 4641 4206 4644
rect 4148 4635 4206 4641
rect 5276 4616 5304 4644
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6362 4632 6368 4684
rect 6420 4632 6426 4684
rect 6472 4672 6500 4712
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 7837 4743 7895 4749
rect 7837 4740 7849 4743
rect 6932 4712 7849 4740
rect 6932 4672 6960 4712
rect 7837 4709 7849 4712
rect 7883 4709 7895 4743
rect 8772 4740 8800 4780
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9398 4808 9404 4820
rect 9263 4780 9404 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9769 4811 9827 4817
rect 9769 4777 9781 4811
rect 9815 4808 9827 4811
rect 11974 4808 11980 4820
rect 9815 4780 11980 4808
rect 9815 4777 9827 4780
rect 9769 4771 9827 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 12250 4808 12256 4820
rect 12207 4780 12256 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12618 4808 12624 4820
rect 12579 4780 12624 4808
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12759 4780 13093 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 13449 4811 13507 4817
rect 13449 4777 13461 4811
rect 13495 4808 13507 4811
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 13495 4780 14381 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 14369 4777 14381 4780
rect 14415 4777 14427 4811
rect 14826 4808 14832 4820
rect 14739 4780 14832 4808
rect 14369 4771 14427 4777
rect 14826 4768 14832 4780
rect 14884 4808 14890 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 14884 4780 15301 4808
rect 14884 4768 14890 4780
rect 15289 4777 15301 4780
rect 15335 4808 15347 4811
rect 16114 4808 16120 4820
rect 15335 4780 16120 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 10686 4740 10692 4752
rect 8772 4712 10692 4740
rect 7837 4703 7895 4709
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 10904 4743 10962 4749
rect 10904 4709 10916 4743
rect 10950 4740 10962 4743
rect 11330 4740 11336 4752
rect 10950 4712 11336 4740
rect 10950 4709 10962 4712
rect 10904 4703 10962 4709
rect 11330 4700 11336 4712
rect 11388 4740 11394 4752
rect 11388 4712 11744 4740
rect 11388 4700 11394 4712
rect 6472 4644 6960 4672
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4672 7067 4675
rect 7374 4672 7380 4684
rect 7055 4644 7380 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 9214 4672 9220 4684
rect 8619 4644 9220 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4672 9367 4675
rect 9766 4672 9772 4684
rect 9355 4644 9772 4672
rect 9355 4641 9367 4644
rect 9309 4635 9367 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 11422 4672 11428 4684
rect 10152 4644 11428 4672
rect 2222 4604 2228 4616
rect 2183 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4564 2286 4616
rect 3510 4604 3516 4616
rect 3471 4576 3516 4604
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 5316 4576 5457 4604
rect 5316 4564 5322 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5592 4576 5641 4604
rect 5592 4564 5598 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 6380 4604 6408 4632
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6380 4576 6469 4604
rect 5629 4567 5687 4573
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 7650 4604 7656 4616
rect 7331 4576 7656 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 7926 4604 7932 4616
rect 7887 4576 7932 4604
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8168 4576 8213 4604
rect 8168 4564 8174 4576
rect 8478 4564 8484 4616
rect 8536 4604 8542 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 8536 4576 9597 4604
rect 8536 4564 8542 4576
rect 9585 4573 9597 4576
rect 9631 4604 9643 4607
rect 10152 4604 10180 4644
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 11606 4672 11612 4684
rect 11567 4644 11612 4672
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 11716 4672 11744 4712
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 14093 4743 14151 4749
rect 14093 4740 14105 4743
rect 12124 4712 14105 4740
rect 12124 4700 12130 4712
rect 14093 4709 14105 4712
rect 14139 4740 14151 4743
rect 14737 4743 14795 4749
rect 14737 4740 14749 4743
rect 14139 4712 14749 4740
rect 14139 4709 14151 4712
rect 14093 4703 14151 4709
rect 14737 4709 14749 4712
rect 14783 4740 14795 4743
rect 17402 4740 17408 4752
rect 14783 4712 17408 4740
rect 14783 4709 14795 4712
rect 14737 4703 14795 4709
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 17586 4700 17592 4752
rect 17644 4740 17650 4752
rect 17957 4743 18015 4749
rect 17957 4740 17969 4743
rect 17644 4712 17969 4740
rect 17644 4700 17650 4712
rect 17957 4709 17969 4712
rect 18003 4709 18015 4743
rect 17957 4703 18015 4709
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18325 4743 18383 4749
rect 18325 4740 18337 4743
rect 18104 4712 18337 4740
rect 18104 4700 18110 4712
rect 18325 4709 18337 4712
rect 18371 4709 18383 4743
rect 18325 4703 18383 4709
rect 13541 4675 13599 4681
rect 11716 4644 11836 4672
rect 11808 4616 11836 4644
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 14458 4672 14464 4684
rect 13587 4644 14464 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 18138 4672 18144 4684
rect 18099 4644 18144 4672
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 9631 4576 10180 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11698 4604 11704 4616
rect 11204 4576 11249 4604
rect 11659 4576 11704 4604
rect 11204 4564 11210 4576
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11790 4564 11796 4616
rect 11848 4604 11854 4616
rect 11848 4576 11941 4604
rect 11848 4564 11854 4576
rect 12250 4564 12256 4616
rect 12308 4564 12314 4616
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12400 4576 12817 4604
rect 12400 4564 12406 4576
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13814 4604 13820 4616
rect 13771 4576 13820 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14001 4607 14059 4613
rect 14001 4573 14013 4607
rect 14047 4604 14059 4607
rect 14274 4604 14280 4616
rect 14047 4576 14280 4604
rect 14047 4573 14059 4576
rect 14001 4567 14059 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4604 15071 4607
rect 15102 4604 15108 4616
rect 15059 4576 15108 4604
rect 15059 4573 15071 4576
rect 15013 4567 15071 4573
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 6365 4539 6423 4545
rect 5184 4508 6316 4536
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 5184 4468 5212 4508
rect 6288 4480 6316 4508
rect 6365 4505 6377 4539
rect 6411 4536 6423 4539
rect 6546 4536 6552 4548
rect 6411 4508 6552 4536
rect 6411 4505 6423 4508
rect 6365 4499 6423 4505
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 6696 4508 6741 4536
rect 6696 4496 6702 4508
rect 7466 4496 7472 4548
rect 7524 4536 7530 4548
rect 8665 4539 8723 4545
rect 8665 4536 8677 4539
rect 7524 4508 8677 4536
rect 7524 4496 7530 4508
rect 8665 4505 8677 4508
rect 8711 4505 8723 4539
rect 8665 4499 8723 4505
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 9674 4536 9680 4548
rect 9539 4508 9680 4536
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 11241 4539 11299 4545
rect 11241 4505 11253 4539
rect 11287 4536 11299 4539
rect 11606 4536 11612 4548
rect 11287 4508 11612 4536
rect 11287 4505 11299 4508
rect 11241 4499 11299 4505
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 12268 4536 12296 4564
rect 18506 4536 18512 4548
rect 11716 4508 13584 4536
rect 18467 4508 18512 4536
rect 2915 4440 5212 4468
rect 5261 4471 5319 4477
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 5350 4468 5356 4480
rect 5307 4440 5356 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 5500 4440 6101 4468
rect 5500 4428 5506 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 6270 4428 6276 4480
rect 6328 4428 6334 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 8294 4468 8300 4480
rect 6880 4440 8300 4468
rect 6880 4428 6886 4440
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 8849 4471 8907 4477
rect 8849 4468 8861 4471
rect 8444 4440 8861 4468
rect 8444 4428 8450 4440
rect 8849 4437 8861 4440
rect 8895 4437 8907 4471
rect 8849 4431 8907 4437
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 10962 4468 10968 4480
rect 9088 4440 10968 4468
rect 9088 4428 9094 4440
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 11716 4468 11744 4508
rect 12250 4468 12256 4480
rect 11388 4440 11744 4468
rect 12211 4440 12256 4468
rect 11388 4428 11394 4440
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 13556 4468 13584 4508
rect 18506 4496 18512 4508
rect 18564 4496 18570 4548
rect 13998 4468 14004 4480
rect 13556 4440 14004 4468
rect 13998 4428 14004 4440
rect 14056 4468 14062 4480
rect 15470 4468 15476 4480
rect 14056 4440 15476 4468
rect 14056 4428 14062 4440
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 3786 4264 3792 4276
rect 3528 4236 3792 4264
rect 3528 4137 3556 4236
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 6362 4264 6368 4276
rect 4856 4236 6368 4264
rect 4856 4224 4862 4236
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 7653 4267 7711 4273
rect 7653 4233 7665 4267
rect 7699 4264 7711 4267
rect 7926 4264 7932 4276
rect 7699 4236 7932 4264
rect 7699 4233 7711 4236
rect 7653 4227 7711 4233
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 8662 4224 8668 4276
rect 8720 4224 8726 4276
rect 9122 4264 9128 4276
rect 9083 4236 9128 4264
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 10965 4267 11023 4273
rect 10965 4233 10977 4267
rect 11011 4264 11023 4267
rect 11238 4264 11244 4276
rect 11011 4236 11244 4264
rect 11011 4233 11023 4236
rect 10965 4227 11023 4233
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 13906 4264 13912 4276
rect 11348 4236 13912 4264
rect 4893 4199 4951 4205
rect 4893 4165 4905 4199
rect 4939 4165 4951 4199
rect 4893 4159 4951 4165
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 4908 4128 4936 4159
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 6380 4196 6408 4224
rect 8680 4196 8708 4224
rect 5408 4168 6132 4196
rect 6380 4168 7779 4196
rect 8680 4168 10640 4196
rect 5408 4156 5414 4168
rect 5258 4128 5264 4140
rect 4908 4100 5264 4128
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 3528 4060 3556 4091
rect 2087 4032 3556 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4908 4060 4936 4100
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5500 4100 5672 4128
rect 5500 4088 5506 4100
rect 4212 4032 4936 4060
rect 5077 4063 5135 4069
rect 4212 4020 4218 4032
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5534 4060 5540 4072
rect 5123 4032 5540 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 1578 3992 1584 4004
rect 1539 3964 1584 3992
rect 1578 3952 1584 3964
rect 1636 3952 1642 4004
rect 2222 3952 2228 4004
rect 2280 4001 2286 4004
rect 2280 3995 2344 4001
rect 2280 3961 2298 3995
rect 2332 3961 2344 3995
rect 2280 3955 2344 3961
rect 3758 3995 3816 4001
rect 3758 3961 3770 3995
rect 3804 3961 3816 3995
rect 3758 3955 3816 3961
rect 2280 3952 2286 3955
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2130 3924 2136 3936
rect 1995 3896 2136 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 3418 3924 3424 3936
rect 3379 3896 3424 3924
rect 3418 3884 3424 3896
rect 3476 3924 3482 3936
rect 3773 3924 3801 3955
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 5092 3992 5120 4023
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5644 4060 5672 4100
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5776 4100 6009 4128
rect 5776 4088 5782 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 6104 4128 6132 4168
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6104 4100 7021 4128
rect 5997 4091 6055 4097
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7751 4128 7779 4168
rect 7751 4100 7880 4128
rect 7009 4091 7067 4097
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 5644 4032 6837 4060
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 7282 4060 7288 4072
rect 7243 4032 7288 4060
rect 6825 4023 6883 4029
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4029 7803 4063
rect 7852 4060 7880 4100
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9784 4137 9812 4168
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9640 4100 9689 4128
rect 9640 4088 9646 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10612 4137 10640 4168
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 11348 4196 11376 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 14458 4264 14464 4276
rect 14419 4236 14464 4264
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 15470 4264 15476 4276
rect 15431 4236 15476 4264
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 10928 4168 11376 4196
rect 13541 4199 13599 4205
rect 10928 4156 10934 4168
rect 13541 4165 13553 4199
rect 13587 4196 13599 4199
rect 14369 4199 14427 4205
rect 13587 4168 13952 4196
rect 13587 4165 13599 4168
rect 13541 4159 13599 4165
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10376 4100 10517 4128
rect 10376 4088 10382 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11606 4128 11612 4140
rect 11204 4100 11612 4128
rect 11204 4088 11210 4100
rect 11606 4088 11612 4100
rect 11664 4128 11670 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11664 4100 11713 4128
rect 11664 4088 11670 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 13814 4128 13820 4140
rect 13775 4100 13820 4128
rect 11701 4091 11759 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 13924 4137 13952 4168
rect 14369 4165 14381 4199
rect 14415 4196 14427 4199
rect 17497 4199 17555 4205
rect 14415 4168 14964 4196
rect 14415 4165 14427 4168
rect 14369 4159 14427 4165
rect 14936 4137 14964 4168
rect 17497 4165 17509 4199
rect 17543 4165 17555 4199
rect 17497 4159 17555 4165
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 14921 4131 14979 4137
rect 13955 4100 14136 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 10410 4060 10416 4072
rect 7852 4032 8148 4060
rect 10371 4032 10416 4060
rect 7745 4023 7803 4029
rect 6917 3995 6975 4001
rect 6917 3992 6929 3995
rect 4764 3964 5120 3992
rect 5920 3964 6929 3992
rect 4764 3952 4770 3964
rect 3476 3896 3801 3924
rect 3476 3884 3482 3896
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 4672 3896 5457 3924
rect 4672 3884 4678 3896
rect 5445 3893 5457 3896
rect 5491 3924 5503 3927
rect 5718 3924 5724 3936
rect 5491 3896 5724 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 5920 3933 5948 3964
rect 6917 3961 6929 3964
rect 6963 3961 6975 3995
rect 7760 3992 7788 4023
rect 8018 4001 8024 4004
rect 8012 3992 8024 4001
rect 6917 3955 6975 3961
rect 7300 3964 7788 3992
rect 7979 3964 8024 3992
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3893 5963 3927
rect 6454 3924 6460 3936
rect 6415 3896 6460 3924
rect 5905 3887 5963 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 6730 3924 6736 3936
rect 6604 3896 6736 3924
rect 6604 3884 6610 3896
rect 6730 3884 6736 3896
rect 6788 3924 6794 3936
rect 7300 3924 7328 3964
rect 8012 3955 8024 3964
rect 8018 3952 8024 3955
rect 8076 3952 8082 4004
rect 8120 3992 8148 4032
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 11974 4069 11980 4072
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4060 11115 4063
rect 11103 4032 11928 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 11900 4004 11928 4032
rect 11968 4023 11980 4069
rect 12032 4060 12038 4072
rect 13998 4060 14004 4072
rect 12032 4032 12068 4060
rect 13959 4032 14004 4060
rect 11974 4020 11980 4023
rect 12032 4020 12038 4032
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14108 4060 14136 4100
rect 14921 4097 14933 4131
rect 14967 4097 14979 4131
rect 15102 4128 15108 4140
rect 15063 4100 15108 4128
rect 14921 4091 14979 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 15252 4100 16681 4128
rect 15252 4088 15258 4100
rect 16669 4097 16681 4100
rect 16715 4128 16727 4131
rect 17512 4128 17540 4159
rect 16715 4100 17356 4128
rect 17512 4100 18368 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 16574 4060 16580 4072
rect 14108 4032 14964 4060
rect 16535 4032 16580 4060
rect 11238 3992 11244 4004
rect 8120 3964 11244 3992
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 11882 3992 11888 4004
rect 11795 3964 11888 3992
rect 11882 3952 11888 3964
rect 11940 3992 11946 4004
rect 12158 3992 12164 4004
rect 11940 3964 12164 3992
rect 11940 3952 11946 3964
rect 12158 3952 12164 3964
rect 12216 3952 12222 4004
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 14936 3992 14964 4032
rect 16574 4020 16580 4032
rect 16632 4060 16638 4072
rect 17328 4069 17356 4100
rect 17037 4063 17095 4069
rect 17037 4060 17049 4063
rect 16632 4032 17049 4060
rect 16632 4020 16638 4032
rect 17037 4029 17049 4032
rect 17083 4029 17095 4063
rect 17037 4023 17095 4029
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17402 4020 17408 4072
rect 17460 4060 17466 4072
rect 18340 4069 18368 4100
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 17460 4032 17601 4060
rect 17460 4020 17466 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4029 18383 4063
rect 18325 4023 18383 4029
rect 16850 3992 16856 4004
rect 13780 3964 14872 3992
rect 14936 3964 16856 3992
rect 13780 3952 13786 3964
rect 7466 3924 7472 3936
rect 6788 3896 7328 3924
rect 7427 3896 7472 3924
rect 6788 3884 6794 3896
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9582 3924 9588 3936
rect 9272 3896 9317 3924
rect 9543 3896 9588 3924
rect 9272 3884 9278 3896
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 11204 3896 11345 3924
rect 11204 3884 11210 3896
rect 11333 3893 11345 3896
rect 11379 3893 11391 3927
rect 11333 3887 11391 3893
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11974 3924 11980 3936
rect 11480 3896 11980 3924
rect 11480 3884 11486 3896
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 12342 3884 12348 3936
rect 12400 3924 12406 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12400 3896 13093 3924
rect 12400 3884 12406 3896
rect 13081 3893 13093 3896
rect 13127 3893 13139 3927
rect 13262 3924 13268 3936
rect 13223 3896 13268 3924
rect 13081 3887 13139 3893
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 14844 3933 14872 3964
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 17957 3995 18015 4001
rect 17957 3992 17969 3995
rect 17236 3964 17969 3992
rect 14829 3927 14887 3933
rect 14829 3893 14841 3927
rect 14875 3924 14887 3927
rect 15381 3927 15439 3933
rect 15381 3924 15393 3927
rect 14875 3896 15393 3924
rect 14875 3893 14887 3896
rect 14829 3887 14887 3893
rect 15381 3893 15393 3896
rect 15427 3924 15439 3927
rect 16666 3924 16672 3936
rect 15427 3896 16672 3924
rect 15427 3893 15439 3896
rect 15381 3887 15439 3893
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 17236 3933 17264 3964
rect 17957 3961 17969 3964
rect 18003 3961 18015 3995
rect 18138 3992 18144 4004
rect 18099 3964 18144 3992
rect 17957 3955 18015 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18506 3992 18512 4004
rect 18467 3964 18512 3992
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 17221 3927 17279 3933
rect 17221 3893 17233 3927
rect 17267 3893 17279 3927
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17221 3887 17279 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 3326 3720 3332 3732
rect 1596 3692 3188 3720
rect 3287 3692 3332 3720
rect 1596 3661 1624 3692
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3621 1639 3655
rect 1581 3615 1639 3621
rect 2317 3655 2375 3661
rect 2317 3621 2329 3655
rect 2363 3652 2375 3655
rect 2590 3652 2596 3664
rect 2363 3624 2596 3652
rect 2363 3621 2375 3624
rect 2317 3615 2375 3621
rect 2590 3612 2596 3624
rect 2648 3612 2654 3664
rect 2866 3652 2872 3664
rect 2827 3624 2872 3652
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 3053 3655 3111 3661
rect 3053 3652 3065 3655
rect 3016 3624 3065 3652
rect 3016 3612 3022 3624
rect 3053 3621 3065 3624
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3553 2007 3587
rect 1949 3547 2007 3553
rect 1964 3448 1992 3547
rect 2406 3544 2412 3596
rect 2464 3584 2470 3596
rect 2685 3587 2743 3593
rect 2685 3584 2697 3587
rect 2464 3556 2697 3584
rect 2464 3544 2470 3556
rect 2685 3553 2697 3556
rect 2731 3553 2743 3587
rect 3160 3584 3188 3692
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4709 3723 4767 3729
rect 4709 3720 4721 3723
rect 3712 3692 4721 3720
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 3421 3655 3479 3661
rect 3421 3652 3433 3655
rect 3292 3624 3433 3652
rect 3292 3612 3298 3624
rect 3421 3621 3433 3624
rect 3467 3621 3479 3655
rect 3421 3615 3479 3621
rect 3712 3584 3740 3692
rect 4709 3689 4721 3692
rect 4755 3689 4767 3723
rect 4709 3683 4767 3689
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 6638 3720 6644 3732
rect 4948 3692 6644 3720
rect 4948 3680 4954 3692
rect 4154 3652 4160 3664
rect 3160 3556 3740 3584
rect 4080 3624 4160 3652
rect 2685 3547 2743 3553
rect 2498 3516 2504 3528
rect 2459 3488 2504 3516
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3694 3516 3700 3528
rect 3292 3488 3700 3516
rect 3292 3476 3298 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 4080 3525 4108 3624
rect 4154 3612 4160 3624
rect 4212 3612 4218 3664
rect 4246 3584 4252 3596
rect 4207 3556 4252 3584
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4893 3587 4951 3593
rect 4893 3553 4905 3587
rect 4939 3584 4951 3587
rect 5074 3584 5080 3596
rect 4939 3556 5080 3584
rect 4939 3553 4951 3556
rect 4893 3547 4951 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5175 3593 5203 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 7432 3692 7481 3720
rect 7432 3680 7438 3692
rect 7469 3689 7481 3692
rect 7515 3689 7527 3723
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7469 3683 7527 3689
rect 7576 3692 7941 3720
rect 6086 3612 6092 3664
rect 6144 3652 6150 3664
rect 7285 3655 7343 3661
rect 7285 3652 7297 3655
rect 6144 3624 7297 3652
rect 6144 3612 6150 3624
rect 7285 3621 7297 3624
rect 7331 3652 7343 3655
rect 7576 3652 7604 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8849 3723 8907 3729
rect 8849 3720 8861 3723
rect 8260 3692 8861 3720
rect 8260 3680 8266 3692
rect 8849 3689 8861 3692
rect 8895 3720 8907 3723
rect 9030 3720 9036 3732
rect 8895 3692 9036 3720
rect 8895 3689 8907 3692
rect 8849 3683 8907 3689
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9125 3723 9183 3729
rect 9125 3689 9137 3723
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 7331 3624 7604 3652
rect 7331 3621 7343 3624
rect 7285 3615 7343 3621
rect 7742 3612 7748 3664
rect 7800 3652 7806 3664
rect 8938 3652 8944 3664
rect 7800 3624 8248 3652
rect 7800 3612 7806 3624
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3553 5227 3587
rect 5169 3547 5227 3553
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 5517 3587 5575 3593
rect 5517 3584 5529 3587
rect 5408 3556 5529 3584
rect 5408 3544 5414 3556
rect 5517 3553 5529 3556
rect 5563 3553 5575 3587
rect 5517 3547 5575 3553
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6788 3556 6929 3584
rect 6788 3544 6794 3556
rect 6917 3553 6929 3556
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3584 7251 3587
rect 7558 3584 7564 3596
rect 7239 3556 7564 3584
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 1964 3420 3740 3448
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1489 3383 1547 3389
rect 1489 3380 1501 3383
rect 1452 3352 1501 3380
rect 1452 3340 1458 3352
rect 1489 3349 1501 3352
rect 1535 3349 1547 3383
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1489 3343 1547 3349
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2222 3380 2228 3392
rect 2183 3352 2228 3380
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 3712 3380 3740 3420
rect 3786 3408 3792 3460
rect 3844 3448 3850 3460
rect 4172 3448 4200 3479
rect 4985 3451 5043 3457
rect 4985 3448 4997 3451
rect 3844 3420 4200 3448
rect 4264 3420 4997 3448
rect 3844 3408 3850 3420
rect 4264 3380 4292 3420
rect 4985 3417 4997 3420
rect 5031 3417 5043 3451
rect 4985 3411 5043 3417
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5276 3448 5304 3479
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 7852 3516 7880 3547
rect 6696 3488 7880 3516
rect 6696 3476 6702 3488
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8220 3516 8248 3624
rect 8312 3624 8944 3652
rect 8312 3593 8340 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3553 8355 3587
rect 8297 3547 8355 3553
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3584 8631 3587
rect 9140 3584 9168 3683
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 9585 3723 9643 3729
rect 9585 3720 9597 3723
rect 9272 3692 9597 3720
rect 9272 3680 9278 3692
rect 9585 3689 9597 3692
rect 9631 3689 9643 3723
rect 9585 3683 9643 3689
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 10870 3720 10876 3732
rect 9732 3692 10180 3720
rect 10831 3692 10876 3720
rect 9732 3680 9738 3692
rect 9493 3655 9551 3661
rect 9493 3621 9505 3655
rect 9539 3652 9551 3655
rect 10042 3652 10048 3664
rect 9539 3624 10048 3652
rect 9539 3621 9551 3624
rect 9493 3615 9551 3621
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 10152 3661 10180 3692
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3720 11299 3723
rect 11698 3720 11704 3732
rect 11287 3692 11704 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 11977 3723 12035 3729
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 13170 3720 13176 3732
rect 12023 3692 13176 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 10137 3655 10195 3661
rect 10137 3621 10149 3655
rect 10183 3621 10195 3655
rect 10137 3615 10195 3621
rect 10686 3612 10692 3664
rect 10744 3652 10750 3664
rect 11992 3652 12020 3683
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13449 3723 13507 3729
rect 13449 3689 13461 3723
rect 13495 3720 13507 3723
rect 13906 3720 13912 3732
rect 13495 3692 13768 3720
rect 13867 3692 13912 3720
rect 13495 3689 13507 3692
rect 13449 3683 13507 3689
rect 10744 3624 12020 3652
rect 10744 3612 10750 3624
rect 12066 3612 12072 3664
rect 12124 3652 12130 3664
rect 13740 3652 13768 3692
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 15102 3680 15108 3732
rect 15160 3720 15166 3732
rect 15749 3723 15807 3729
rect 15749 3720 15761 3723
rect 15160 3692 15761 3720
rect 15160 3680 15166 3692
rect 15749 3689 15761 3692
rect 15795 3689 15807 3723
rect 15749 3683 15807 3689
rect 13814 3652 13820 3664
rect 12124 3624 12572 3652
rect 13727 3624 13820 3652
rect 12124 3612 12130 3624
rect 10502 3584 10508 3596
rect 8619 3556 9168 3584
rect 9232 3556 10508 3584
rect 8619 3553 8631 3556
rect 8573 3547 8631 3553
rect 9232 3516 9260 3556
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 10870 3544 10876 3596
rect 10928 3544 10934 3596
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11388 3556 11713 3584
rect 11388 3544 11394 3556
rect 11701 3553 11713 3556
rect 11747 3553 11759 3587
rect 11701 3547 11759 3553
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 12342 3593 12348 3596
rect 12325 3587 12348 3593
rect 12325 3584 12337 3587
rect 11940 3556 12337 3584
rect 11940 3544 11946 3556
rect 12325 3553 12337 3556
rect 12325 3547 12348 3553
rect 12342 3544 12348 3547
rect 12400 3544 12406 3596
rect 12544 3584 12572 3624
rect 13814 3612 13820 3624
rect 13872 3652 13878 3664
rect 14614 3655 14672 3661
rect 14614 3652 14626 3655
rect 13872 3624 14626 3652
rect 13872 3612 13878 3624
rect 14614 3621 14626 3624
rect 14660 3621 14672 3655
rect 16390 3652 16396 3664
rect 16351 3624 16396 3652
rect 14614 3615 14672 3621
rect 16390 3612 16396 3624
rect 16448 3652 16454 3664
rect 16448 3624 17632 3652
rect 16448 3612 16454 3624
rect 17604 3593 17632 3624
rect 17770 3612 17776 3664
rect 17828 3652 17834 3664
rect 17957 3655 18015 3661
rect 17957 3652 17969 3655
rect 17828 3624 17969 3652
rect 17828 3612 17834 3624
rect 17957 3621 17969 3624
rect 18003 3621 18015 3655
rect 17957 3615 18015 3621
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 12544 3556 16221 3584
rect 16209 3553 16221 3556
rect 16255 3584 16267 3587
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 16255 3556 16957 3584
rect 16255 3553 16267 3556
rect 16209 3547 16267 3553
rect 16945 3553 16957 3556
rect 16991 3553 17003 3587
rect 16945 3547 17003 3553
rect 17221 3587 17279 3593
rect 17221 3553 17233 3587
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 17589 3587 17647 3593
rect 17589 3553 17601 3587
rect 17635 3553 17647 3587
rect 18325 3587 18383 3593
rect 18325 3584 18337 3587
rect 17589 3547 17647 3553
rect 17788 3556 18337 3584
rect 8076 3488 8121 3516
rect 8220 3488 9260 3516
rect 8076 3476 8082 3488
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9548 3488 9689 3516
rect 9548 3476 9554 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 10594 3516 10600 3528
rect 10555 3488 10600 3516
rect 9677 3479 9735 3485
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3485 10839 3519
rect 10888 3516 10916 3544
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10888 3488 11437 3516
rect 10781 3479 10839 3485
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 7742 3448 7748 3460
rect 5224 3420 5304 3448
rect 6196 3420 7748 3448
rect 5224 3408 5230 3420
rect 6196 3392 6224 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 8757 3451 8815 3457
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 9306 3448 9312 3460
rect 8803 3420 9312 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 9306 3408 9312 3420
rect 9364 3408 9370 3460
rect 9398 3408 9404 3460
rect 9456 3448 9462 3460
rect 9953 3451 10011 3457
rect 9953 3448 9965 3451
rect 9456 3420 9965 3448
rect 9456 3408 9462 3420
rect 9953 3417 9965 3420
rect 9999 3417 10011 3451
rect 9953 3411 10011 3417
rect 10796 3448 10824 3479
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11664 3488 12081 3516
rect 11664 3476 11670 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 14366 3516 14372 3528
rect 14327 3488 14372 3516
rect 12069 3479 12127 3485
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 16666 3516 16672 3528
rect 16579 3488 16672 3516
rect 16666 3476 16672 3488
rect 16724 3516 16730 3528
rect 17236 3516 17264 3547
rect 16724 3488 17264 3516
rect 16724 3476 16730 3488
rect 10870 3448 10876 3460
rect 10796 3420 10876 3448
rect 4614 3380 4620 3392
rect 3712 3352 4292 3380
rect 4575 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 5442 3380 5448 3392
rect 4764 3352 5448 3380
rect 4764 3340 4770 3352
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 6178 3340 6184 3392
rect 6236 3340 6242 3392
rect 6638 3380 6644 3392
rect 6599 3352 6644 3380
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 7009 3383 7067 3389
rect 6788 3352 6833 3380
rect 6788 3340 6794 3352
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 7190 3380 7196 3392
rect 7055 3352 7196 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8662 3380 8668 3392
rect 8527 3352 8668 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 9674 3380 9680 3392
rect 8996 3352 9680 3380
rect 8996 3340 9002 3352
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 10413 3383 10471 3389
rect 10413 3349 10425 3383
rect 10459 3380 10471 3383
rect 10796 3380 10824 3420
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 10962 3408 10968 3460
rect 11020 3448 11026 3460
rect 11517 3451 11575 3457
rect 11517 3448 11529 3451
rect 11020 3420 11529 3448
rect 11020 3408 11026 3420
rect 11517 3417 11529 3420
rect 11563 3448 11575 3451
rect 16758 3448 16764 3460
rect 11563 3420 12112 3448
rect 11563 3417 11575 3420
rect 11517 3411 11575 3417
rect 10459 3352 10824 3380
rect 12084 3380 12112 3420
rect 13556 3420 13860 3448
rect 12342 3380 12348 3392
rect 12084 3352 12348 3380
rect 10459 3349 10471 3352
rect 10413 3343 10471 3349
rect 12342 3340 12348 3352
rect 12400 3380 12406 3392
rect 13556 3380 13584 3420
rect 12400 3352 13584 3380
rect 13633 3383 13691 3389
rect 12400 3340 12406 3352
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 13722 3380 13728 3392
rect 13679 3352 13728 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13832 3380 13860 3420
rect 16408 3420 16764 3448
rect 16408 3380 16436 3420
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 17788 3457 17816 3556
rect 18325 3553 18337 3556
rect 18371 3553 18383 3587
rect 18325 3547 18383 3553
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 17920 3488 18521 3516
rect 17920 3476 17926 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 17773 3451 17831 3457
rect 17773 3417 17785 3451
rect 17819 3417 17831 3451
rect 18138 3448 18144 3460
rect 18099 3420 18144 3448
rect 17773 3411 17831 3417
rect 18138 3408 18144 3420
rect 18196 3408 18202 3460
rect 16850 3380 16856 3392
rect 13832 3352 16436 3380
rect 16811 3352 16856 3380
rect 16850 3340 16856 3352
rect 16908 3340 16914 3392
rect 17129 3383 17187 3389
rect 17129 3349 17141 3383
rect 17175 3380 17187 3383
rect 17310 3380 17316 3392
rect 17175 3352 17316 3380
rect 17175 3349 17187 3352
rect 17129 3343 17187 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17405 3383 17463 3389
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 18322 3380 18328 3392
rect 17451 3352 18328 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 1636 3148 3740 3176
rect 1636 3136 1642 3148
rect 2869 3111 2927 3117
rect 2869 3077 2881 3111
rect 2915 3077 2927 3111
rect 3712 3108 3740 3148
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 3844 3148 3893 3176
rect 3844 3136 3850 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 3881 3139 3939 3145
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3176 4031 3179
rect 4246 3176 4252 3188
rect 4019 3148 4252 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 5994 3176 6000 3188
rect 4580 3148 6000 3176
rect 4580 3136 4586 3148
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 7929 3179 7987 3185
rect 6196 3148 7604 3176
rect 5629 3111 5687 3117
rect 5629 3108 5641 3111
rect 3712 3080 5641 3108
rect 2869 3071 2927 3077
rect 5629 3077 5641 3080
rect 5675 3077 5687 3111
rect 5629 3071 5687 3077
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2884 2972 2912 3071
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3418 3040 3424 3052
rect 3375 3012 3424 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3418 3000 3424 3012
rect 3476 3040 3482 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 3476 3012 4629 3040
rect 3476 3000 3482 3012
rect 4617 3009 4629 3012
rect 4663 3040 4675 3043
rect 4890 3040 4896 3052
rect 4663 3012 4896 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5092 3012 5273 3040
rect 1995 2944 2912 2972
rect 3053 2975 3111 2981
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 3053 2941 3065 2975
rect 3099 2972 3111 2975
rect 3510 2972 3516 2984
rect 3099 2944 3516 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 3752 2944 4353 2972
rect 3752 2932 3758 2944
rect 4341 2941 4353 2944
rect 4387 2972 4399 2975
rect 4706 2972 4712 2984
rect 4387 2944 4712 2972
rect 4387 2941 4399 2944
rect 4341 2935 4399 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 5092 2972 5120 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5408 3012 5453 3040
rect 5408 3000 5414 3012
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6196 3040 6224 3148
rect 5776 3012 6224 3040
rect 5776 3000 5782 3012
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 7576 3040 7604 3148
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8018 3176 8024 3188
rect 7975 3148 8024 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8938 3176 8944 3188
rect 8899 3148 8944 3176
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 10410 3176 10416 3188
rect 10091 3148 10416 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 10410 3136 10416 3148
rect 10468 3176 10474 3188
rect 11054 3176 11060 3188
rect 10468 3148 11060 3176
rect 10468 3136 10474 3148
rect 11054 3136 11060 3148
rect 11112 3176 11118 3188
rect 11974 3176 11980 3188
rect 11112 3148 11980 3176
rect 11112 3136 11118 3148
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 12124 3148 13553 3176
rect 12124 3136 12130 3148
rect 13541 3145 13553 3148
rect 13587 3176 13599 3179
rect 13725 3179 13783 3185
rect 13725 3176 13737 3179
rect 13587 3148 13737 3176
rect 13587 3145 13599 3148
rect 13541 3139 13599 3145
rect 13725 3145 13737 3148
rect 13771 3145 13783 3179
rect 13725 3139 13783 3145
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14826 3176 14832 3188
rect 13872 3148 14832 3176
rect 13872 3136 13878 3148
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 15562 3176 15568 3188
rect 15523 3148 15568 3176
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 11882 3108 11888 3120
rect 9232 3080 11888 3108
rect 9232 3049 9260 3080
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 12802 3108 12808 3120
rect 11992 3080 12808 3108
rect 9217 3043 9275 3049
rect 6328 3012 6684 3040
rect 7576 3012 8984 3040
rect 6328 3000 6334 3012
rect 4856 2944 5120 2972
rect 5169 2975 5227 2981
rect 4856 2932 4862 2944
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5810 2972 5816 2984
rect 5215 2944 5816 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6089 2975 6147 2981
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 6178 2972 6184 2984
rect 6135 2944 6184 2972
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 6546 2972 6552 2984
rect 6507 2944 6552 2972
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6656 2972 6684 3012
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 6656 2944 8217 2972
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 8205 2935 8263 2941
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 8846 2972 8852 2984
rect 8803 2944 8852 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 382 2864 388 2916
rect 440 2904 446 2916
rect 1397 2907 1455 2913
rect 1397 2904 1409 2907
rect 440 2876 1409 2904
rect 440 2864 446 2876
rect 1397 2873 1409 2876
rect 1443 2873 1455 2907
rect 1762 2904 1768 2916
rect 1723 2876 1768 2904
rect 1397 2867 1455 2873
rect 1762 2864 1768 2876
rect 1820 2864 1826 2916
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 2317 2907 2375 2913
rect 2317 2904 2329 2907
rect 2188 2876 2329 2904
rect 2188 2864 2194 2876
rect 2317 2873 2329 2876
rect 2363 2873 2375 2907
rect 2317 2867 2375 2873
rect 2685 2907 2743 2913
rect 2685 2873 2697 2907
rect 2731 2904 2743 2907
rect 2731 2876 5948 2904
rect 2731 2873 2743 2876
rect 2685 2867 2743 2873
rect 2222 2836 2228 2848
rect 2183 2808 2228 2836
rect 2222 2796 2228 2808
rect 2280 2796 2286 2848
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 2774 2836 2780 2848
rect 2639 2808 2780 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 3421 2839 3479 2845
rect 3421 2836 3433 2839
rect 3292 2808 3433 2836
rect 3292 2796 3298 2808
rect 3421 2805 3433 2808
rect 3467 2805 3479 2839
rect 3421 2799 3479 2805
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 4522 2836 4528 2848
rect 4479 2808 4528 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 4798 2836 4804 2848
rect 4759 2808 4804 2836
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 5350 2836 5356 2848
rect 4948 2808 5356 2836
rect 4948 2796 4954 2808
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 5920 2845 5948 2876
rect 6638 2864 6644 2916
rect 6696 2904 6702 2916
rect 6794 2907 6852 2913
rect 6794 2904 6806 2907
rect 6696 2876 6806 2904
rect 6696 2864 6702 2876
rect 6794 2873 6806 2876
rect 6840 2873 6852 2907
rect 6794 2867 6852 2873
rect 7650 2864 7656 2916
rect 7708 2904 7714 2916
rect 8496 2904 8524 2935
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 8956 2972 8984 3012
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 9217 3003 9275 3009
rect 9324 3012 10609 3040
rect 9324 2972 9352 3012
rect 10597 3009 10609 3012
rect 10643 3040 10655 3043
rect 10686 3040 10692 3052
rect 10643 3012 10692 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 11054 3040 11060 3052
rect 10827 3012 11060 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 11054 3000 11060 3012
rect 11112 3040 11118 3052
rect 11790 3040 11796 3052
rect 11112 3012 11796 3040
rect 11112 3000 11118 3012
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11992 3049 12020 3080
rect 12802 3068 12808 3080
rect 12860 3068 12866 3120
rect 13170 3108 13176 3120
rect 13131 3080 13176 3108
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 13262 3068 13268 3120
rect 13320 3108 13326 3120
rect 13909 3111 13967 3117
rect 13909 3108 13921 3111
rect 13320 3080 13921 3108
rect 13320 3068 13326 3080
rect 13909 3077 13921 3080
rect 13955 3077 13967 3111
rect 13909 3071 13967 3077
rect 16850 3068 16856 3120
rect 16908 3108 16914 3120
rect 17770 3108 17776 3120
rect 16908 3080 17264 3108
rect 17731 3080 17776 3108
rect 16908 3068 16914 3080
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12158 3000 12164 3052
rect 12216 3040 12222 3052
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 12216 3012 16037 3040
rect 12216 3000 12222 3012
rect 16025 3009 16037 3012
rect 16071 3040 16083 3043
rect 16071 3012 17172 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 8956 2944 9352 2972
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 11517 2975 11575 2981
rect 9447 2944 11468 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 7708 2876 8524 2904
rect 9309 2907 9367 2913
rect 7708 2864 7714 2876
rect 9309 2873 9321 2907
rect 9355 2904 9367 2907
rect 9858 2904 9864 2916
rect 9355 2876 9864 2904
rect 9355 2873 9367 2876
rect 9309 2867 9367 2873
rect 9858 2864 9864 2876
rect 9916 2864 9922 2916
rect 10318 2864 10324 2916
rect 10376 2904 10382 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 10376 2876 10977 2904
rect 10376 2864 10382 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 10965 2867 11023 2873
rect 11149 2907 11207 2913
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 11440 2904 11468 2944
rect 11517 2941 11529 2975
rect 11563 2972 11575 2975
rect 12250 2972 12256 2984
rect 11563 2944 12256 2972
rect 11563 2941 11575 2944
rect 11517 2935 11575 2941
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12618 2932 12624 2984
rect 12676 2972 12682 2984
rect 13081 2975 13139 2981
rect 13081 2972 13093 2975
rect 12676 2944 13093 2972
rect 12676 2932 12682 2944
rect 13081 2941 13093 2944
rect 13127 2941 13139 2975
rect 13081 2935 13139 2941
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 13228 2944 13369 2972
rect 13228 2932 13234 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 14093 2975 14151 2981
rect 14093 2972 14105 2975
rect 13688 2944 14105 2972
rect 13688 2932 13694 2944
rect 14093 2941 14105 2944
rect 14139 2941 14151 2975
rect 16298 2972 16304 2984
rect 16259 2944 16304 2972
rect 14093 2935 14151 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2972 16819 2975
rect 17034 2972 17040 2984
rect 16807 2944 17040 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17144 2981 17172 3012
rect 17236 2981 17264 3080
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17368 3012 17632 3040
rect 17368 3000 17374 3012
rect 17604 2981 17632 3012
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 17736 3012 18521 3040
rect 17736 3000 17742 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 17589 2975 17647 2981
rect 17589 2941 17601 2975
rect 17635 2941 17647 2975
rect 17957 2975 18015 2981
rect 17957 2972 17969 2975
rect 17589 2935 17647 2941
rect 17696 2944 17969 2972
rect 11882 2904 11888 2916
rect 11195 2876 11376 2904
rect 11440 2876 11888 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 5905 2839 5963 2845
rect 5905 2805 5917 2839
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 6052 2808 6193 2836
rect 6052 2796 6058 2808
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 6181 2799 6239 2805
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 8021 2839 8079 2845
rect 8021 2836 8033 2839
rect 6328 2808 8033 2836
rect 6328 2796 6334 2808
rect 8021 2805 8033 2808
rect 8067 2805 8079 2839
rect 8294 2836 8300 2848
rect 8255 2808 8300 2836
rect 8021 2799 8079 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 8570 2836 8576 2848
rect 8531 2808 8576 2836
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 10134 2836 10140 2848
rect 10095 2808 10140 2836
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 11348 2845 11376 2876
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 12158 2864 12164 2916
rect 12216 2904 12222 2916
rect 12529 2907 12587 2913
rect 12529 2904 12541 2907
rect 12216 2876 12541 2904
rect 12216 2864 12222 2876
rect 12529 2873 12541 2876
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 12713 2907 12771 2913
rect 12713 2873 12725 2907
rect 12759 2873 12771 2907
rect 12713 2867 12771 2873
rect 10505 2839 10563 2845
rect 10505 2836 10517 2839
rect 10468 2808 10517 2836
rect 10468 2796 10474 2808
rect 10505 2805 10517 2808
rect 10551 2805 10563 2839
rect 10505 2799 10563 2805
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2805 11391 2839
rect 11333 2799 11391 2805
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12342 2836 12348 2848
rect 12115 2808 12348 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12728 2836 12756 2867
rect 12802 2864 12808 2916
rect 12860 2904 12866 2916
rect 13648 2904 13676 2932
rect 12860 2876 13676 2904
rect 12860 2864 12866 2876
rect 15838 2864 15844 2916
rect 15896 2904 15902 2916
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 15896 2876 16497 2904
rect 15896 2864 15902 2876
rect 16485 2873 16497 2876
rect 16531 2904 16543 2907
rect 16531 2876 17264 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 17236 2848 17264 2876
rect 17494 2864 17500 2916
rect 17552 2904 17558 2916
rect 17696 2904 17724 2944
rect 17957 2941 17969 2944
rect 18003 2941 18015 2975
rect 18322 2972 18328 2984
rect 18283 2944 18328 2972
rect 17957 2935 18015 2941
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 17552 2876 17724 2904
rect 17552 2864 17558 2876
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12492 2808 12537 2836
rect 12728 2808 12909 2836
rect 12492 2796 12498 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 15746 2836 15752 2848
rect 15707 2808 15752 2836
rect 12897 2799 12955 2805
rect 15746 2796 15752 2808
rect 15804 2796 15810 2848
rect 16114 2836 16120 2848
rect 16075 2808 16120 2836
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 16942 2836 16948 2848
rect 16903 2808 16948 2836
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17218 2796 17224 2848
rect 17276 2796 17282 2848
rect 17402 2836 17408 2848
rect 17363 2808 17408 2836
rect 17402 2796 17408 2808
rect 17460 2796 17466 2848
rect 17586 2796 17592 2848
rect 17644 2836 17650 2848
rect 18049 2839 18107 2845
rect 18049 2836 18061 2839
rect 17644 2808 18061 2836
rect 17644 2796 17650 2808
rect 18049 2805 18061 2808
rect 18095 2805 18107 2839
rect 18049 2799 18107 2805
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 4249 2635 4307 2641
rect 4249 2601 4261 2635
rect 4295 2632 4307 2635
rect 4709 2635 4767 2641
rect 4709 2632 4721 2635
rect 4295 2604 4721 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 4709 2601 4721 2604
rect 4755 2601 4767 2635
rect 4709 2595 4767 2601
rect 4798 2592 4804 2644
rect 4856 2632 4862 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 4856 2604 5181 2632
rect 4856 2592 4862 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5169 2595 5227 2601
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6454 2632 6460 2644
rect 5951 2604 6460 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 8846 2632 8852 2644
rect 7392 2604 8852 2632
rect 1210 2524 1216 2576
rect 1268 2564 1274 2576
rect 2133 2567 2191 2573
rect 2133 2564 2145 2567
rect 1268 2536 2145 2564
rect 1268 2524 1274 2536
rect 2133 2533 2145 2536
rect 2179 2533 2191 2567
rect 2314 2564 2320 2576
rect 2275 2536 2320 2564
rect 2133 2527 2191 2533
rect 2314 2524 2320 2536
rect 2372 2524 2378 2576
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 4614 2564 4620 2576
rect 4203 2536 4620 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 6270 2564 6276 2576
rect 4724 2536 6276 2564
rect 2038 2496 2044 2508
rect 1999 2468 2044 2496
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2682 2496 2688 2508
rect 2643 2468 2688 2496
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2465 3295 2499
rect 3510 2496 3516 2508
rect 3471 2468 3516 2496
rect 3237 2459 3295 2465
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 1946 2428 1952 2440
rect 1903 2400 1952 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 1946 2388 1952 2400
rect 2004 2388 2010 2440
rect 3252 2428 3280 2459
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 4724 2496 4752 2536
rect 6270 2524 6276 2536
rect 6328 2524 6334 2576
rect 6362 2524 6368 2576
rect 6420 2564 6426 2576
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 6420 2536 6745 2564
rect 6420 2524 6426 2536
rect 6733 2533 6745 2536
rect 6779 2533 6791 2567
rect 7392 2564 7420 2604
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 9088 2604 9597 2632
rect 9088 2592 9094 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9858 2632 9864 2644
rect 9819 2604 9864 2632
rect 9585 2595 9643 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 10192 2604 10241 2632
rect 10192 2592 10198 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10229 2595 10287 2601
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2632 10379 2635
rect 10410 2632 10416 2644
rect 10367 2604 10416 2632
rect 10367 2601 10379 2604
rect 10321 2595 10379 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11146 2632 11152 2644
rect 11103 2604 11152 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2601 11483 2635
rect 11698 2632 11704 2644
rect 11659 2604 11704 2632
rect 11425 2595 11483 2601
rect 6733 2527 6791 2533
rect 6932 2536 7420 2564
rect 6932 2508 6960 2536
rect 7466 2524 7472 2576
rect 7524 2564 7530 2576
rect 8205 2567 8263 2573
rect 8205 2564 8217 2567
rect 7524 2536 8217 2564
rect 7524 2524 7530 2536
rect 8205 2533 8217 2536
rect 8251 2533 8263 2567
rect 8389 2567 8447 2573
rect 8389 2564 8401 2567
rect 8205 2527 8263 2533
rect 8312 2536 8401 2564
rect 5074 2496 5080 2508
rect 4540 2468 4752 2496
rect 5035 2468 5080 2496
rect 4065 2431 4123 2437
rect 2056 2400 3188 2428
rect 3252 2400 3924 2428
rect 1489 2363 1547 2369
rect 1489 2329 1501 2363
rect 1535 2360 1547 2363
rect 2056 2360 2084 2400
rect 1535 2332 2084 2360
rect 1535 2329 1547 2332
rect 1489 2323 1547 2329
rect 2130 2320 2136 2372
rect 2188 2360 2194 2372
rect 2501 2363 2559 2369
rect 2501 2360 2513 2363
rect 2188 2332 2513 2360
rect 2188 2320 2194 2332
rect 2501 2329 2513 2332
rect 2547 2329 2559 2363
rect 3050 2360 3056 2372
rect 3011 2332 3056 2360
rect 2501 2323 2559 2329
rect 3050 2320 3056 2332
rect 3108 2320 3114 2372
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 2958 2292 2964 2304
rect 2096 2264 2964 2292
rect 2096 2252 2102 2264
rect 2958 2252 2964 2264
rect 3016 2252 3022 2304
rect 3160 2292 3188 2400
rect 3697 2363 3755 2369
rect 3697 2329 3709 2363
rect 3743 2360 3755 2363
rect 3786 2360 3792 2372
rect 3743 2332 3792 2360
rect 3743 2329 3755 2332
rect 3697 2323 3755 2329
rect 3786 2320 3792 2332
rect 3844 2320 3850 2372
rect 3896 2360 3924 2400
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4430 2428 4436 2440
rect 4111 2400 4436 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 4540 2360 4568 2468
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5813 2499 5871 2505
rect 5813 2496 5825 2499
rect 5184 2468 5825 2496
rect 5184 2428 5212 2468
rect 5813 2465 5825 2468
rect 5859 2465 5871 2499
rect 6914 2496 6920 2508
rect 6827 2468 6920 2496
rect 5813 2459 5871 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 8312 2496 8340 2536
rect 8389 2533 8401 2536
rect 8435 2533 8447 2567
rect 8570 2564 8576 2576
rect 8531 2536 8576 2564
rect 8389 2527 8447 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 8662 2524 8668 2576
rect 8720 2564 8726 2576
rect 8941 2567 8999 2573
rect 8941 2564 8953 2567
rect 8720 2536 8953 2564
rect 8720 2524 8726 2536
rect 8941 2533 8953 2536
rect 8987 2533 8999 2567
rect 8941 2527 8999 2533
rect 9306 2524 9312 2576
rect 9364 2564 9370 2576
rect 9401 2567 9459 2573
rect 9401 2564 9413 2567
rect 9364 2536 9413 2564
rect 9364 2524 9370 2536
rect 9401 2533 9413 2536
rect 9447 2533 9459 2567
rect 9401 2527 9459 2533
rect 10965 2567 11023 2573
rect 10965 2533 10977 2567
rect 11011 2564 11023 2567
rect 11330 2564 11336 2576
rect 11011 2536 11336 2564
rect 11011 2533 11023 2536
rect 10965 2527 11023 2533
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 11440 2564 11468 2595
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12345 2635 12403 2641
rect 12345 2601 12357 2635
rect 12391 2632 12403 2635
rect 12434 2632 12440 2644
rect 12391 2604 12440 2632
rect 12391 2601 12403 2604
rect 12345 2595 12403 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 13449 2635 13507 2641
rect 13449 2601 13461 2635
rect 13495 2601 13507 2635
rect 14553 2635 14611 2641
rect 14553 2632 14565 2635
rect 13449 2595 13507 2601
rect 14108 2604 14565 2632
rect 12253 2567 12311 2573
rect 12253 2564 12265 2567
rect 11440 2536 12265 2564
rect 12253 2533 12265 2536
rect 12299 2533 12311 2567
rect 12253 2527 12311 2533
rect 13265 2567 13323 2573
rect 13265 2533 13277 2567
rect 13311 2564 13323 2567
rect 13464 2564 13492 2595
rect 14108 2573 14136 2604
rect 14553 2601 14565 2604
rect 14599 2601 14611 2635
rect 15197 2635 15255 2641
rect 15197 2632 15209 2635
rect 14553 2595 14611 2601
rect 15028 2604 15209 2632
rect 15028 2573 15056 2604
rect 15197 2601 15209 2604
rect 15243 2601 15255 2635
rect 15654 2632 15660 2644
rect 15615 2604 15660 2632
rect 15197 2595 15255 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 17494 2632 17500 2644
rect 16255 2604 17500 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 13311 2536 13492 2564
rect 14093 2567 14151 2573
rect 13311 2533 13323 2536
rect 13265 2527 13323 2533
rect 14093 2533 14105 2567
rect 14139 2533 14151 2567
rect 14093 2527 14151 2533
rect 15013 2567 15071 2573
rect 15013 2533 15025 2567
rect 15059 2533 15071 2567
rect 15013 2527 15071 2533
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 16393 2567 16451 2573
rect 15620 2536 16068 2564
rect 15620 2524 15626 2536
rect 11054 2496 11060 2508
rect 7024 2468 8340 2496
rect 8404 2468 9628 2496
rect 4632 2400 5212 2428
rect 4632 2369 4660 2400
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 5721 2431 5779 2437
rect 5316 2400 5361 2428
rect 5316 2388 5322 2400
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 6638 2428 6644 2440
rect 5767 2400 6644 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7024 2428 7052 2468
rect 6788 2400 7052 2428
rect 7745 2431 7803 2437
rect 6788 2388 6794 2400
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 8404 2428 8432 2468
rect 7791 2400 8432 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 8536 2400 9229 2428
rect 8536 2388 8542 2400
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 9600 2428 9628 2468
rect 10888 2468 11060 2496
rect 10226 2428 10232 2440
rect 9600 2400 10232 2428
rect 9217 2391 9275 2397
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10888 2437 10916 2468
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11514 2496 11520 2508
rect 11475 2468 11520 2496
rect 11514 2456 11520 2468
rect 11572 2456 11578 2508
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 11756 2468 12909 2496
rect 11756 2456 11762 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 13412 2468 13645 2496
rect 13412 2456 13418 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 14642 2456 14648 2508
rect 14700 2496 14706 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14700 2468 14749 2496
rect 14700 2456 14706 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 15378 2496 15384 2508
rect 15339 2468 15384 2496
rect 14737 2459 14795 2465
rect 15378 2456 15384 2468
rect 15436 2456 15442 2508
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 15654 2496 15660 2508
rect 15519 2468 15660 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 15749 2499 15807 2505
rect 15749 2465 15761 2499
rect 15795 2496 15807 2499
rect 15838 2496 15844 2508
rect 15795 2468 15844 2496
rect 15795 2465 15807 2468
rect 15749 2459 15807 2465
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 16040 2505 16068 2536
rect 16393 2533 16405 2567
rect 16439 2564 16451 2567
rect 16942 2564 16948 2576
rect 16439 2536 16948 2564
rect 16439 2533 16451 2536
rect 16393 2527 16451 2533
rect 16942 2524 16948 2536
rect 17000 2524 17006 2576
rect 17402 2524 17408 2576
rect 17460 2564 17466 2576
rect 17589 2567 17647 2573
rect 17589 2564 17601 2567
rect 17460 2536 17601 2564
rect 17460 2524 17466 2536
rect 17589 2533 17601 2536
rect 17635 2533 17647 2567
rect 17589 2527 17647 2533
rect 18230 2524 18236 2576
rect 18288 2564 18294 2576
rect 18325 2567 18383 2573
rect 18325 2564 18337 2567
rect 18288 2536 18337 2564
rect 18288 2524 18294 2536
rect 18325 2533 18337 2536
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 16025 2499 16083 2505
rect 16025 2465 16037 2499
rect 16071 2465 16083 2499
rect 16025 2459 16083 2465
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 16853 2499 16911 2505
rect 16853 2496 16865 2499
rect 16632 2468 16865 2496
rect 16632 2456 16638 2468
rect 16853 2465 16865 2468
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17221 2499 17279 2505
rect 17221 2496 17233 2499
rect 17092 2468 17233 2496
rect 17092 2456 17098 2468
rect 17221 2465 17233 2468
rect 17267 2465 17279 2499
rect 17221 2459 17279 2465
rect 17957 2499 18015 2505
rect 17957 2465 17969 2499
rect 18003 2465 18015 2499
rect 17957 2459 18015 2465
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10873 2431 10931 2437
rect 10551 2400 10824 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 3896 2332 4568 2360
rect 4617 2363 4675 2369
rect 4617 2329 4629 2363
rect 4663 2329 4675 2363
rect 4617 2323 4675 2329
rect 4890 2320 4896 2372
rect 4948 2360 4954 2372
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 4948 2332 6561 2360
rect 4948 2320 4954 2332
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 6549 2323 6607 2329
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 8757 2363 8815 2369
rect 8757 2360 8769 2363
rect 7616 2332 8769 2360
rect 7616 2320 7622 2332
rect 8757 2329 8769 2332
rect 8803 2329 8815 2363
rect 8757 2323 8815 2329
rect 5074 2292 5080 2304
rect 3160 2264 5080 2292
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 6270 2292 6276 2304
rect 6231 2264 6276 2292
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 6420 2264 8125 2292
rect 6420 2252 6426 2264
rect 8113 2261 8125 2264
rect 8159 2261 8171 2295
rect 10796 2292 10824 2400
rect 10873 2397 10885 2431
rect 10919 2397 10931 2431
rect 12434 2428 12440 2440
rect 12395 2400 12440 2428
rect 10873 2391 10931 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 11238 2320 11244 2372
rect 11296 2360 11302 2372
rect 12713 2363 12771 2369
rect 12713 2360 12725 2363
rect 11296 2332 12725 2360
rect 11296 2320 11302 2332
rect 12713 2329 12725 2332
rect 12759 2329 12771 2363
rect 13078 2360 13084 2372
rect 13039 2332 13084 2360
rect 12713 2323 12771 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 13906 2360 13912 2372
rect 13867 2332 13912 2360
rect 13906 2320 13912 2332
rect 13964 2320 13970 2372
rect 14826 2360 14832 2372
rect 14787 2332 14832 2360
rect 14826 2320 14832 2332
rect 14884 2320 14890 2372
rect 15286 2320 15292 2372
rect 15344 2360 15350 2372
rect 15933 2363 15991 2369
rect 15933 2360 15945 2363
rect 15344 2332 15945 2360
rect 15344 2320 15350 2332
rect 15933 2329 15945 2332
rect 15979 2329 15991 2363
rect 15933 2323 15991 2329
rect 16574 2320 16580 2372
rect 16632 2360 16638 2372
rect 17405 2363 17463 2369
rect 16632 2332 16677 2360
rect 16632 2320 16638 2332
rect 17405 2329 17417 2363
rect 17451 2360 17463 2363
rect 17972 2360 18000 2459
rect 18506 2360 18512 2372
rect 17451 2332 18000 2360
rect 18467 2332 18512 2360
rect 17451 2329 17463 2332
rect 17405 2323 17463 2329
rect 18506 2320 18512 2332
rect 18564 2320 18570 2372
rect 11422 2292 11428 2304
rect 10796 2264 11428 2292
rect 8113 2255 8171 2261
rect 11422 2252 11428 2264
rect 11480 2292 11486 2304
rect 12434 2292 12440 2304
rect 11480 2264 12440 2292
rect 11480 2252 11486 2264
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 16666 2252 16672 2304
rect 16724 2292 16730 2304
rect 16761 2295 16819 2301
rect 16761 2292 16773 2295
rect 16724 2264 16773 2292
rect 16724 2252 16730 2264
rect 16761 2261 16773 2264
rect 16807 2261 16819 2295
rect 16761 2255 16819 2261
rect 17494 2252 17500 2304
rect 17552 2292 17558 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17552 2264 17693 2292
rect 17552 2252 17558 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 18049 2295 18107 2301
rect 18049 2292 18061 2295
rect 17828 2264 18061 2292
rect 17828 2252 17834 2264
rect 18049 2261 18061 2264
rect 18095 2261 18107 2295
rect 18049 2255 18107 2261
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 3510 2048 3516 2100
rect 3568 2088 3574 2100
rect 8294 2088 8300 2100
rect 3568 2060 8300 2088
rect 3568 2048 3574 2060
rect 8294 2048 8300 2060
rect 8352 2048 8358 2100
rect 2958 1980 2964 2032
rect 3016 2020 3022 2032
rect 6914 2020 6920 2032
rect 3016 1992 6920 2020
rect 3016 1980 3022 1992
rect 6914 1980 6920 1992
rect 6972 1980 6978 2032
rect 2682 1912 2688 1964
rect 2740 1952 2746 1964
rect 7282 1952 7288 1964
rect 2740 1924 7288 1952
rect 2740 1912 2746 1924
rect 7282 1912 7288 1924
rect 7340 1912 7346 1964
rect 1946 1844 1952 1896
rect 2004 1884 2010 1896
rect 5902 1884 5908 1896
rect 2004 1856 5908 1884
rect 2004 1844 2010 1856
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 6270 1844 6276 1896
rect 6328 1884 6334 1896
rect 7650 1884 7656 1896
rect 6328 1856 7656 1884
rect 6328 1844 6334 1856
rect 7650 1844 7656 1856
rect 7708 1844 7714 1896
rect 5074 1776 5080 1828
rect 5132 1816 5138 1828
rect 10502 1816 10508 1828
rect 5132 1788 10508 1816
rect 5132 1776 5138 1788
rect 10502 1776 10508 1788
rect 10560 1776 10566 1828
rect 9674 1708 9680 1760
rect 9732 1748 9738 1760
rect 19426 1748 19432 1760
rect 9732 1720 19432 1748
rect 9732 1708 9738 1720
rect 19426 1708 19432 1720
rect 19484 1708 19490 1760
rect 17218 1504 17224 1556
rect 17276 1544 17282 1556
rect 17586 1544 17592 1556
rect 17276 1516 17592 1544
rect 17276 1504 17282 1516
rect 17586 1504 17592 1516
rect 17644 1504 17650 1556
<< via1 >>
rect 15292 14900 15344 14952
rect 17776 14900 17828 14952
rect 2320 14832 2372 14884
rect 12716 14832 12768 14884
rect 15476 14832 15528 14884
rect 16396 14832 16448 14884
rect 4068 14764 4120 14816
rect 17224 14764 17276 14816
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 2596 14560 2648 14612
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 7748 14560 7800 14612
rect 1860 14535 1912 14544
rect 1860 14501 1869 14535
rect 1869 14501 1903 14535
rect 1903 14501 1912 14535
rect 1860 14492 1912 14501
rect 2228 14535 2280 14544
rect 2228 14501 2237 14535
rect 2237 14501 2271 14535
rect 2271 14501 2280 14535
rect 2228 14492 2280 14501
rect 3608 14535 3660 14544
rect 3608 14501 3617 14535
rect 3617 14501 3651 14535
rect 3651 14501 3660 14535
rect 3608 14492 3660 14501
rect 5540 14535 5592 14544
rect 5540 14501 5549 14535
rect 5549 14501 5583 14535
rect 5583 14501 5592 14535
rect 5540 14492 5592 14501
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2504 14424 2556 14476
rect 2872 14424 2924 14476
rect 2964 14424 3016 14476
rect 2688 14356 2740 14408
rect 3240 14356 3292 14408
rect 3424 14424 3476 14476
rect 9956 14535 10008 14544
rect 9956 14501 9965 14535
rect 9965 14501 9999 14535
rect 9999 14501 10008 14535
rect 9956 14492 10008 14501
rect 12164 14535 12216 14544
rect 12164 14501 12173 14535
rect 12173 14501 12207 14535
rect 12207 14501 12216 14535
rect 12164 14492 12216 14501
rect 14372 14492 14424 14544
rect 3516 14356 3568 14408
rect 11520 14424 11572 14476
rect 12348 14467 12400 14476
rect 12348 14433 12357 14467
rect 12357 14433 12391 14467
rect 12391 14433 12400 14467
rect 12348 14424 12400 14433
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 15016 14424 15068 14476
rect 16580 14560 16632 14612
rect 16212 14492 16264 14544
rect 16396 14492 16448 14544
rect 17408 14492 17460 14544
rect 18052 14535 18104 14544
rect 18052 14501 18061 14535
rect 18061 14501 18095 14535
rect 18095 14501 18104 14535
rect 18052 14492 18104 14501
rect 17224 14467 17276 14476
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 2504 14288 2556 14340
rect 3608 14288 3660 14340
rect 3332 14220 3384 14272
rect 8208 14288 8260 14340
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 15200 14288 15252 14340
rect 17224 14433 17233 14467
rect 17233 14433 17267 14467
rect 17267 14433 17276 14467
rect 17224 14424 17276 14433
rect 17684 14467 17736 14476
rect 17684 14433 17693 14467
rect 17693 14433 17727 14467
rect 17727 14433 17736 14467
rect 17684 14424 17736 14433
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 16120 14356 16172 14408
rect 16672 14288 16724 14340
rect 14924 14220 14976 14272
rect 15384 14263 15436 14272
rect 15384 14229 15393 14263
rect 15393 14229 15427 14263
rect 15427 14229 15436 14263
rect 15384 14220 15436 14229
rect 18788 14356 18840 14408
rect 17224 14288 17276 14340
rect 18052 14288 18104 14340
rect 18144 14220 18196 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 1492 14016 1544 14068
rect 3240 14016 3292 14068
rect 3516 14059 3568 14068
rect 3516 14025 3525 14059
rect 3525 14025 3559 14059
rect 3559 14025 3568 14059
rect 3516 14016 3568 14025
rect 11520 14016 11572 14068
rect 12072 14016 12124 14068
rect 14740 14016 14792 14068
rect 15016 14059 15068 14068
rect 15016 14025 15025 14059
rect 15025 14025 15059 14059
rect 15059 14025 15068 14059
rect 15016 14016 15068 14025
rect 15292 14016 15344 14068
rect 15476 14016 15528 14068
rect 17960 14016 18012 14068
rect 8116 13948 8168 14000
rect 14924 13948 14976 14000
rect 16396 13948 16448 14000
rect 16488 13948 16540 14000
rect 2688 13880 2740 13932
rect 5632 13880 5684 13932
rect 10508 13880 10560 13932
rect 15384 13880 15436 13932
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 1124 13744 1176 13796
rect 1952 13744 2004 13796
rect 2872 13812 2924 13864
rect 11704 13812 11756 13864
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 15016 13744 15068 13796
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 2596 13676 2648 13728
rect 5080 13676 5132 13728
rect 5172 13676 5224 13728
rect 15292 13676 15344 13728
rect 15844 13787 15896 13796
rect 15844 13753 15853 13787
rect 15853 13753 15887 13787
rect 15887 13753 15896 13787
rect 15844 13744 15896 13753
rect 16028 13744 16080 13796
rect 17316 13880 17368 13932
rect 16948 13812 17000 13864
rect 17776 13880 17828 13932
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 17960 13812 18012 13864
rect 18420 13855 18472 13864
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 17592 13744 17644 13796
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 1952 13472 2004 13524
rect 3056 13472 3108 13524
rect 3332 13472 3384 13524
rect 3700 13472 3752 13524
rect 1860 13447 1912 13456
rect 1860 13413 1869 13447
rect 1869 13413 1903 13447
rect 1903 13413 1912 13447
rect 1860 13404 1912 13413
rect 6368 13404 6420 13456
rect 13820 13472 13872 13524
rect 14372 13472 14424 13524
rect 15108 13472 15160 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 15844 13472 15896 13524
rect 16396 13472 16448 13524
rect 16580 13515 16632 13524
rect 16580 13481 16589 13515
rect 16589 13481 16623 13515
rect 16623 13481 16632 13515
rect 16580 13472 16632 13481
rect 16764 13472 16816 13524
rect 17592 13472 17644 13524
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 3332 13336 3384 13388
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 4988 13336 5040 13388
rect 5080 13336 5132 13388
rect 11520 13404 11572 13456
rect 6644 13336 6696 13388
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 11888 13336 11940 13388
rect 14740 13379 14792 13388
rect 14740 13345 14749 13379
rect 14749 13345 14783 13379
rect 14783 13345 14792 13379
rect 14740 13336 14792 13345
rect 15200 13404 15252 13456
rect 3056 13268 3108 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 7472 13268 7524 13320
rect 8024 13268 8076 13320
rect 8852 13268 8904 13320
rect 9588 13268 9640 13320
rect 3240 13200 3292 13252
rect 4620 13200 4672 13252
rect 8484 13200 8536 13252
rect 13360 13268 13412 13320
rect 15660 13268 15712 13320
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 4344 13175 4396 13184
rect 4344 13141 4353 13175
rect 4353 13141 4387 13175
rect 4387 13141 4396 13175
rect 4344 13132 4396 13141
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 8944 13132 8996 13184
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 11520 13175 11572 13184
rect 9220 13132 9272 13141
rect 11520 13141 11529 13175
rect 11529 13141 11563 13175
rect 11563 13141 11572 13175
rect 11520 13132 11572 13141
rect 14096 13200 14148 13252
rect 14556 13200 14608 13252
rect 14832 13200 14884 13252
rect 15292 13200 15344 13252
rect 15384 13243 15436 13252
rect 15384 13209 15393 13243
rect 15393 13209 15427 13243
rect 15427 13209 15436 13243
rect 16212 13336 16264 13388
rect 17040 13447 17092 13456
rect 17040 13413 17049 13447
rect 17049 13413 17083 13447
rect 17083 13413 17092 13447
rect 17040 13404 17092 13413
rect 17684 13379 17736 13388
rect 16396 13268 16448 13320
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 17960 13268 18012 13320
rect 15384 13200 15436 13209
rect 15016 13132 15068 13184
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 4712 12928 4764 12980
rect 6644 12971 6696 12980
rect 6644 12937 6653 12971
rect 6653 12937 6687 12971
rect 6687 12937 6696 12971
rect 6644 12928 6696 12937
rect 8300 12928 8352 12980
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 12348 12928 12400 12980
rect 8116 12903 8168 12912
rect 1400 12792 1452 12844
rect 8116 12869 8125 12903
rect 8125 12869 8159 12903
rect 8159 12869 8168 12903
rect 8116 12860 8168 12869
rect 8576 12860 8628 12912
rect 11152 12860 11204 12912
rect 14740 12928 14792 12980
rect 14832 12928 14884 12980
rect 15660 12928 15712 12980
rect 16212 12928 16264 12980
rect 2872 12724 2924 12776
rect 5080 12792 5132 12844
rect 5540 12792 5592 12844
rect 5908 12792 5960 12844
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 1492 12699 1544 12708
rect 1492 12665 1501 12699
rect 1501 12665 1535 12699
rect 1535 12665 1544 12699
rect 1492 12656 1544 12665
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 3516 12656 3568 12708
rect 5816 12656 5868 12708
rect 6368 12656 6420 12708
rect 7748 12767 7800 12776
rect 7748 12733 7766 12767
rect 7766 12733 7800 12767
rect 7748 12724 7800 12733
rect 2228 12588 2280 12640
rect 4436 12588 4488 12640
rect 5724 12588 5776 12640
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 9496 12656 9548 12708
rect 10416 12724 10468 12776
rect 10692 12724 10744 12776
rect 13360 12724 13412 12776
rect 14004 12860 14056 12912
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 17500 12792 17552 12844
rect 11520 12656 11572 12708
rect 10600 12588 10652 12640
rect 11428 12631 11480 12640
rect 11428 12597 11437 12631
rect 11437 12597 11471 12631
rect 11471 12597 11480 12631
rect 11428 12588 11480 12597
rect 12072 12631 12124 12640
rect 12072 12597 12081 12631
rect 12081 12597 12115 12631
rect 12115 12597 12124 12631
rect 12072 12588 12124 12597
rect 14004 12656 14056 12708
rect 15108 12699 15160 12708
rect 14096 12588 14148 12640
rect 14280 12631 14332 12640
rect 14280 12597 14289 12631
rect 14289 12597 14323 12631
rect 14323 12597 14332 12631
rect 15108 12665 15117 12699
rect 15117 12665 15151 12699
rect 15151 12665 15160 12699
rect 15108 12656 15160 12665
rect 14280 12588 14332 12597
rect 14924 12588 14976 12640
rect 15660 12724 15712 12776
rect 16580 12724 16632 12776
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 18512 12767 18564 12776
rect 18512 12733 18521 12767
rect 18521 12733 18555 12767
rect 18555 12733 18564 12767
rect 18512 12724 18564 12733
rect 15476 12656 15528 12708
rect 16488 12588 16540 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 18972 12495 19024 12504
rect 18972 12461 18981 12495
rect 18981 12461 19015 12495
rect 19015 12461 19024 12495
rect 18972 12452 19024 12461
rect 3516 12427 3568 12436
rect 3516 12393 3525 12427
rect 3525 12393 3559 12427
rect 3559 12393 3568 12427
rect 3516 12384 3568 12393
rect 4896 12384 4948 12436
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 5080 12384 5132 12393
rect 6736 12384 6788 12436
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 9588 12427 9640 12436
rect 9588 12393 9597 12427
rect 9597 12393 9631 12427
rect 9631 12393 9640 12427
rect 9588 12384 9640 12393
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 1400 12248 1452 12300
rect 2228 12248 2280 12300
rect 3516 12248 3568 12300
rect 3700 12248 3752 12300
rect 4712 12248 4764 12300
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 3884 12180 3936 12232
rect 2872 12044 2924 12096
rect 3700 12044 3752 12096
rect 4252 12044 4304 12096
rect 4896 12180 4948 12232
rect 7288 12316 7340 12368
rect 7748 12359 7800 12368
rect 7748 12325 7757 12359
rect 7757 12325 7791 12359
rect 7791 12325 7800 12359
rect 7748 12316 7800 12325
rect 9404 12316 9456 12368
rect 9496 12316 9548 12368
rect 5540 12180 5592 12232
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 8484 12180 8536 12232
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9772 12248 9824 12300
rect 10784 12316 10836 12368
rect 11428 12316 11480 12368
rect 13360 12384 13412 12436
rect 12072 12316 12124 12368
rect 13268 12316 13320 12368
rect 17868 12384 17920 12436
rect 18420 12384 18472 12436
rect 14556 12316 14608 12368
rect 15292 12316 15344 12368
rect 15660 12316 15712 12368
rect 16580 12316 16632 12368
rect 16856 12316 16908 12368
rect 17316 12316 17368 12368
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 10416 12223 10468 12232
rect 4988 12112 5040 12164
rect 6184 12112 6236 12164
rect 5448 12044 5500 12096
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 6000 12044 6052 12096
rect 6828 12044 6880 12096
rect 8392 12112 8444 12164
rect 8668 12044 8720 12096
rect 9220 12044 9272 12096
rect 9588 12112 9640 12164
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 11888 12248 11940 12300
rect 12532 12248 12584 12300
rect 10324 12112 10376 12164
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 17776 12248 17828 12300
rect 14556 12112 14608 12164
rect 16856 12180 16908 12232
rect 16580 12112 16632 12164
rect 12072 12044 12124 12096
rect 13912 12044 13964 12096
rect 14924 12044 14976 12096
rect 15108 12044 15160 12096
rect 16212 12044 16264 12096
rect 18328 12087 18380 12096
rect 18328 12053 18337 12087
rect 18337 12053 18371 12087
rect 18371 12053 18380 12087
rect 18328 12044 18380 12053
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 1952 11840 2004 11892
rect 3608 11840 3660 11892
rect 4712 11883 4764 11892
rect 2780 11704 2832 11756
rect 1768 11611 1820 11620
rect 1768 11577 1777 11611
rect 1777 11577 1811 11611
rect 1811 11577 1820 11611
rect 1768 11568 1820 11577
rect 2044 11611 2096 11620
rect 2044 11577 2053 11611
rect 2053 11577 2087 11611
rect 2087 11577 2096 11611
rect 2044 11568 2096 11577
rect 4436 11772 4488 11824
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 5448 11840 5500 11892
rect 8852 11883 8904 11892
rect 6368 11772 6420 11824
rect 6736 11772 6788 11824
rect 8852 11849 8861 11883
rect 8861 11849 8895 11883
rect 8895 11849 8904 11883
rect 8852 11840 8904 11849
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 9772 11840 9824 11892
rect 10324 11840 10376 11892
rect 11888 11772 11940 11824
rect 12532 11840 12584 11892
rect 14280 11840 14332 11892
rect 13820 11772 13872 11824
rect 14096 11772 14148 11824
rect 14832 11840 14884 11892
rect 15476 11840 15528 11892
rect 14556 11772 14608 11824
rect 16028 11772 16080 11824
rect 4252 11704 4304 11756
rect 5540 11704 5592 11756
rect 6644 11704 6696 11756
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 10784 11704 10836 11756
rect 12072 11704 12124 11756
rect 13636 11704 13688 11756
rect 15292 11747 15344 11756
rect 3240 11636 3292 11688
rect 4804 11636 4856 11688
rect 6000 11636 6052 11688
rect 6368 11636 6420 11688
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 8484 11636 8536 11688
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 9404 11636 9456 11688
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 12256 11679 12308 11688
rect 12256 11645 12265 11679
rect 12265 11645 12299 11679
rect 12299 11645 12308 11679
rect 12256 11636 12308 11645
rect 14556 11636 14608 11688
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 16672 11840 16724 11892
rect 17040 11840 17092 11892
rect 17316 11840 17368 11892
rect 17500 11840 17552 11892
rect 17592 11840 17644 11892
rect 18052 11840 18104 11892
rect 16764 11704 16816 11756
rect 17592 11747 17644 11756
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 17776 11704 17828 11756
rect 16488 11636 16540 11688
rect 16580 11636 16632 11688
rect 4160 11568 4212 11620
rect 4344 11568 4396 11620
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 3792 11500 3844 11552
rect 10692 11568 10744 11620
rect 13360 11568 13412 11620
rect 4804 11500 4856 11552
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 8116 11500 8168 11552
rect 8300 11500 8352 11552
rect 9036 11500 9088 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 9588 11500 9640 11552
rect 10968 11500 11020 11552
rect 11060 11500 11112 11552
rect 11244 11500 11296 11552
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12440 11500 12492 11509
rect 12716 11500 12768 11552
rect 13176 11500 13228 11552
rect 13452 11500 13504 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 14004 11543 14056 11552
rect 14004 11509 14013 11543
rect 14013 11509 14047 11543
rect 14047 11509 14056 11543
rect 14004 11500 14056 11509
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 16488 11500 16540 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 17316 11543 17368 11552
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 18144 11543 18196 11552
rect 18144 11509 18153 11543
rect 18153 11509 18187 11543
rect 18187 11509 18196 11543
rect 18144 11500 18196 11509
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 1584 11296 1636 11348
rect 4068 11296 4120 11348
rect 4252 11296 4304 11348
rect 4896 11296 4948 11348
rect 5172 11296 5224 11348
rect 9588 11296 9640 11348
rect 10416 11296 10468 11348
rect 4436 11228 4488 11280
rect 5540 11228 5592 11280
rect 5724 11228 5776 11280
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 3424 11203 3476 11212
rect 3424 11169 3442 11203
rect 3442 11169 3476 11203
rect 3424 11160 3476 11169
rect 6092 11160 6144 11212
rect 6552 11160 6604 11212
rect 7656 11160 7708 11212
rect 8300 11160 8352 11212
rect 8484 11203 8536 11212
rect 8484 11169 8493 11203
rect 8493 11169 8527 11203
rect 8527 11169 8536 11203
rect 8484 11160 8536 11169
rect 8852 11228 8904 11280
rect 10692 11271 10744 11280
rect 10692 11237 10701 11271
rect 10701 11237 10735 11271
rect 10735 11237 10744 11271
rect 10692 11228 10744 11237
rect 10968 11296 11020 11348
rect 11152 11296 11204 11348
rect 11428 11296 11480 11348
rect 12440 11296 12492 11348
rect 13176 11296 13228 11348
rect 14096 11296 14148 11348
rect 14188 11296 14240 11348
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 16764 11339 16816 11348
rect 16764 11305 16773 11339
rect 16773 11305 16807 11339
rect 16807 11305 16816 11339
rect 16764 11296 16816 11305
rect 11060 11203 11112 11212
rect 2320 11092 2372 11144
rect 3700 11135 3752 11144
rect 3700 11101 3709 11135
rect 3709 11101 3743 11135
rect 3743 11101 3752 11135
rect 3700 11092 3752 11101
rect 5632 11092 5684 11144
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 7380 11092 7432 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 11152 11160 11204 11212
rect 11888 11228 11940 11280
rect 12532 11228 12584 11280
rect 13360 11228 13412 11280
rect 12072 11160 12124 11212
rect 12624 11160 12676 11212
rect 13452 11160 13504 11212
rect 17040 11271 17092 11280
rect 17040 11237 17049 11271
rect 17049 11237 17083 11271
rect 17083 11237 17092 11271
rect 17040 11228 17092 11237
rect 17316 11296 17368 11348
rect 17684 11228 17736 11280
rect 18972 11271 19024 11280
rect 18972 11237 18981 11271
rect 18981 11237 19015 11271
rect 19015 11237 19024 11271
rect 18972 11228 19024 11237
rect 7840 11024 7892 11076
rect 2412 10956 2464 11008
rect 2504 10956 2556 11008
rect 4252 10956 4304 11008
rect 5080 10956 5132 11008
rect 6184 10956 6236 11008
rect 7472 10956 7524 11008
rect 11244 11092 11296 11144
rect 10692 11024 10744 11076
rect 11520 11092 11572 11144
rect 11796 11092 11848 11144
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 13176 11092 13228 11144
rect 13636 11092 13688 11144
rect 14372 11135 14424 11144
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 9128 10956 9180 11008
rect 11888 10999 11940 11008
rect 11888 10965 11897 10999
rect 11897 10965 11931 10999
rect 11931 10965 11940 10999
rect 11888 10956 11940 10965
rect 13728 11024 13780 11076
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 13544 10956 13596 11008
rect 13820 10956 13872 11008
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 15016 11160 15068 11212
rect 16028 11160 16080 11212
rect 16488 11160 16540 11212
rect 17960 11203 18012 11212
rect 15108 11092 15160 11144
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 17500 11092 17552 11144
rect 18420 11092 18472 11144
rect 18512 11067 18564 11076
rect 18512 11033 18521 11067
rect 18521 11033 18555 11067
rect 18555 11033 18564 11067
rect 18512 11024 18564 11033
rect 16580 10956 16632 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 1860 10752 1912 10804
rect 2320 10795 2372 10804
rect 2320 10761 2329 10795
rect 2329 10761 2363 10795
rect 2363 10761 2372 10795
rect 2320 10752 2372 10761
rect 3424 10616 3476 10668
rect 5356 10752 5408 10804
rect 7564 10752 7616 10804
rect 7840 10795 7892 10804
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 11520 10752 11572 10804
rect 16856 10752 16908 10804
rect 17592 10752 17644 10804
rect 2596 10548 2648 10600
rect 3608 10548 3660 10600
rect 3792 10548 3844 10600
rect 6368 10548 6420 10600
rect 7472 10548 7524 10600
rect 10508 10684 10560 10736
rect 11244 10684 11296 10736
rect 12072 10684 12124 10736
rect 15016 10684 15068 10736
rect 16212 10659 16264 10668
rect 16212 10625 16221 10659
rect 16221 10625 16255 10659
rect 16255 10625 16264 10659
rect 16212 10616 16264 10625
rect 16488 10616 16540 10668
rect 1860 10412 1912 10464
rect 2136 10412 2188 10464
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 5080 10480 5132 10532
rect 3792 10412 3844 10421
rect 6000 10412 6052 10464
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 6736 10523 6788 10532
rect 6736 10489 6770 10523
rect 6770 10489 6788 10523
rect 6736 10480 6788 10489
rect 7748 10480 7800 10532
rect 10416 10548 10468 10600
rect 10968 10548 11020 10600
rect 11060 10548 11112 10600
rect 11520 10548 11572 10600
rect 11980 10548 12032 10600
rect 9680 10523 9732 10532
rect 7840 10412 7892 10464
rect 8576 10412 8628 10464
rect 9680 10489 9692 10523
rect 9692 10489 9732 10523
rect 9680 10480 9732 10489
rect 11612 10480 11664 10532
rect 12624 10480 12676 10532
rect 13544 10480 13596 10532
rect 17776 10480 17828 10532
rect 13452 10412 13504 10464
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 16028 10412 16080 10464
rect 17592 10412 17644 10464
rect 18604 10412 18656 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 3332 10251 3384 10260
rect 3332 10217 3341 10251
rect 3341 10217 3375 10251
rect 3375 10217 3384 10251
rect 3332 10208 3384 10217
rect 3792 10208 3844 10260
rect 2780 10140 2832 10192
rect 6000 10208 6052 10260
rect 6276 10208 6328 10260
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 7932 10208 7984 10260
rect 8392 10208 8444 10260
rect 9588 10251 9640 10260
rect 9588 10217 9597 10251
rect 9597 10217 9631 10251
rect 9631 10217 9640 10251
rect 9588 10208 9640 10217
rect 5172 10140 5224 10192
rect 5356 10140 5408 10192
rect 2412 10072 2464 10124
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 5632 10115 5684 10124
rect 5632 10081 5641 10115
rect 5641 10081 5675 10115
rect 5675 10081 5684 10115
rect 5632 10072 5684 10081
rect 5080 10047 5132 10056
rect 4160 9979 4212 9988
rect 4160 9945 4169 9979
rect 4169 9945 4203 9979
rect 4203 9945 4212 9979
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 7472 10140 7524 10192
rect 8208 10140 8260 10192
rect 10324 10140 10376 10192
rect 12716 10208 12768 10260
rect 14372 10208 14424 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 17408 10251 17460 10260
rect 17408 10217 17417 10251
rect 17417 10217 17451 10251
rect 17451 10217 17460 10251
rect 17408 10208 17460 10217
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 11888 10140 11940 10192
rect 7104 10072 7156 10124
rect 7748 10072 7800 10124
rect 7840 10072 7892 10124
rect 9496 10072 9548 10124
rect 10508 10072 10560 10124
rect 12072 10072 12124 10124
rect 12716 10072 12768 10124
rect 13452 10140 13504 10192
rect 13268 10072 13320 10124
rect 16948 10140 17000 10192
rect 18604 10140 18656 10192
rect 6736 10047 6788 10056
rect 6736 10013 6745 10047
rect 6745 10013 6779 10047
rect 6779 10013 6788 10047
rect 6736 10004 6788 10013
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 8668 10047 8720 10056
rect 4160 9936 4212 9945
rect 2320 9868 2372 9920
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2964 9911 3016 9920
rect 2780 9868 2832 9877
rect 2964 9877 2973 9911
rect 2973 9877 3007 9911
rect 3007 9877 3016 9911
rect 2964 9868 3016 9877
rect 3240 9868 3292 9920
rect 5172 9868 5224 9920
rect 6460 9868 6512 9920
rect 7104 9868 7156 9920
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 7564 9868 7616 9877
rect 8024 9868 8076 9920
rect 8208 9868 8260 9920
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 11244 10004 11296 10056
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 12256 10047 12308 10056
rect 8392 9936 8444 9988
rect 9772 9936 9824 9988
rect 10508 9936 10560 9988
rect 10784 9936 10836 9988
rect 11152 9936 11204 9988
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 15016 10047 15068 10056
rect 13728 10004 13780 10013
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 15660 10004 15712 10056
rect 16028 10004 16080 10056
rect 17592 10072 17644 10124
rect 18512 10115 18564 10124
rect 18512 10081 18521 10115
rect 18521 10081 18555 10115
rect 18555 10081 18564 10115
rect 18512 10072 18564 10081
rect 12624 9936 12676 9988
rect 8852 9868 8904 9920
rect 11612 9868 11664 9920
rect 12992 9868 13044 9920
rect 13268 9868 13320 9920
rect 13360 9868 13412 9920
rect 14648 9868 14700 9920
rect 14740 9868 14792 9920
rect 15016 9868 15068 9920
rect 16672 9936 16724 9988
rect 17868 10004 17920 10056
rect 17776 9936 17828 9988
rect 18420 10004 18472 10056
rect 17868 9868 17920 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 3608 9664 3660 9716
rect 3792 9707 3844 9716
rect 3792 9673 3801 9707
rect 3801 9673 3835 9707
rect 3835 9673 3844 9707
rect 3792 9664 3844 9673
rect 4344 9664 4396 9716
rect 2780 9596 2832 9648
rect 3884 9596 3936 9648
rect 3976 9596 4028 9648
rect 5172 9596 5224 9648
rect 2964 9528 3016 9580
rect 2228 9503 2280 9512
rect 2228 9469 2237 9503
rect 2237 9469 2271 9503
rect 2271 9469 2280 9503
rect 2228 9460 2280 9469
rect 3148 9460 3200 9512
rect 4988 9528 5040 9580
rect 5540 9596 5592 9648
rect 5724 9596 5776 9648
rect 8392 9664 8444 9716
rect 8576 9664 8628 9716
rect 6920 9596 6972 9648
rect 7656 9639 7708 9648
rect 7656 9605 7665 9639
rect 7665 9605 7699 9639
rect 7699 9605 7708 9639
rect 7656 9596 7708 9605
rect 8300 9596 8352 9648
rect 3976 9503 4028 9512
rect 2872 9392 2924 9444
rect 3332 9435 3384 9444
rect 3332 9401 3341 9435
rect 3341 9401 3375 9435
rect 3375 9401 3384 9435
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4620 9460 4672 9512
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 6092 9528 6144 9580
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7840 9528 7892 9580
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 13452 9664 13504 9716
rect 13728 9707 13780 9716
rect 13728 9673 13737 9707
rect 13737 9673 13771 9707
rect 13771 9673 13780 9707
rect 13728 9664 13780 9673
rect 13820 9664 13872 9716
rect 11060 9596 11112 9648
rect 12072 9596 12124 9648
rect 15660 9664 15712 9716
rect 16396 9664 16448 9716
rect 16672 9664 16724 9716
rect 17132 9664 17184 9716
rect 17592 9664 17644 9716
rect 8208 9528 8260 9537
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 5816 9460 5868 9469
rect 6276 9460 6328 9512
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 3332 9392 3384 9401
rect 3516 9392 3568 9444
rect 8576 9460 8628 9512
rect 8668 9460 8720 9512
rect 9772 9460 9824 9512
rect 10692 9503 10744 9512
rect 10692 9469 10710 9503
rect 10710 9469 10744 9503
rect 10692 9460 10744 9469
rect 11796 9460 11848 9512
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 3976 9324 4028 9376
rect 8024 9435 8076 9444
rect 8024 9401 8033 9435
rect 8033 9401 8067 9435
rect 8067 9401 8076 9435
rect 12624 9435 12676 9444
rect 8024 9392 8076 9401
rect 12624 9401 12658 9435
rect 12658 9401 12676 9435
rect 12624 9392 12676 9401
rect 13820 9435 13872 9444
rect 13820 9401 13829 9435
rect 13829 9401 13863 9435
rect 13863 9401 13872 9435
rect 13820 9392 13872 9401
rect 4712 9324 4764 9376
rect 5080 9324 5132 9376
rect 5540 9324 5592 9376
rect 5908 9324 5960 9376
rect 6092 9324 6144 9376
rect 7288 9324 7340 9376
rect 7932 9324 7984 9376
rect 8300 9324 8352 9376
rect 9680 9324 9732 9376
rect 11244 9324 11296 9376
rect 11612 9324 11664 9376
rect 11888 9324 11940 9376
rect 12348 9324 12400 9376
rect 13452 9324 13504 9376
rect 14740 9460 14792 9512
rect 15200 9392 15252 9444
rect 16488 9460 16540 9512
rect 16028 9392 16080 9444
rect 16212 9392 16264 9444
rect 17408 9392 17460 9444
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 17500 9324 17552 9376
rect 17776 9324 17828 9376
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 2780 9120 2832 9172
rect 3884 9120 3936 9172
rect 4712 9120 4764 9172
rect 3700 9052 3752 9104
rect 4344 9052 4396 9104
rect 6184 9120 6236 9172
rect 7288 9120 7340 9172
rect 8208 9163 8260 9172
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 8576 9120 8628 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9956 9163 10008 9172
rect 9128 9120 9180 9129
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 11244 9120 11296 9172
rect 11428 9120 11480 9172
rect 11520 9120 11572 9172
rect 12072 9120 12124 9172
rect 12256 9120 12308 9172
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 12716 9120 12768 9172
rect 13176 9120 13228 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 13728 9120 13780 9172
rect 8116 9052 8168 9104
rect 8484 9052 8536 9104
rect 11152 9052 11204 9104
rect 1492 9027 1544 9036
rect 1492 8993 1501 9027
rect 1501 8993 1535 9027
rect 1535 8993 1544 9027
rect 1492 8984 1544 8993
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 2320 8984 2372 9036
rect 2780 8984 2832 9036
rect 3976 8984 4028 9036
rect 4620 8984 4672 9036
rect 4712 8984 4764 9036
rect 5632 8984 5684 9036
rect 6092 8984 6144 9036
rect 6368 8984 6420 9036
rect 7840 8984 7892 9036
rect 8300 8984 8352 9036
rect 11612 8984 11664 9036
rect 12348 9052 12400 9104
rect 15660 9120 15712 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 17592 9120 17644 9172
rect 17868 9163 17920 9172
rect 17868 9129 17877 9163
rect 17877 9129 17911 9163
rect 17911 9129 17920 9163
rect 17868 9120 17920 9129
rect 17960 9120 18012 9172
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6276 8916 6328 8968
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 7932 8916 7984 8968
rect 10232 8959 10284 8968
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 5448 8848 5500 8900
rect 3332 8780 3384 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 6736 8823 6788 8832
rect 6736 8789 6745 8823
rect 6745 8789 6779 8823
rect 6779 8789 6788 8823
rect 6736 8780 6788 8789
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8484 8823 8536 8832
rect 8300 8780 8352 8789
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 10416 8823 10468 8832
rect 10416 8789 10425 8823
rect 10425 8789 10459 8823
rect 10459 8789 10468 8823
rect 10416 8780 10468 8789
rect 10692 8848 10744 8900
rect 11060 8916 11112 8968
rect 11520 8916 11572 8968
rect 13820 8984 13872 9036
rect 14832 9027 14884 9036
rect 14832 8993 14841 9027
rect 14841 8993 14875 9027
rect 14875 8993 14884 9027
rect 14832 8984 14884 8993
rect 13452 8959 13504 8968
rect 12532 8848 12584 8900
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 15016 8959 15068 8968
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 17224 9052 17276 9104
rect 15476 8984 15528 9036
rect 16028 9027 16080 9036
rect 16028 8993 16037 9027
rect 16037 8993 16071 9027
rect 16071 8993 16080 9027
rect 16028 8984 16080 8993
rect 15016 8916 15068 8925
rect 13636 8848 13688 8900
rect 14556 8848 14608 8900
rect 12348 8780 12400 8832
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 14372 8780 14424 8832
rect 17408 8891 17460 8900
rect 17408 8857 17417 8891
rect 17417 8857 17451 8891
rect 17451 8857 17460 8891
rect 17408 8848 17460 8857
rect 16948 8780 17000 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2136 8576 2188 8628
rect 3056 8576 3108 8628
rect 5724 8576 5776 8628
rect 6276 8619 6328 8628
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 8024 8576 8076 8628
rect 11796 8576 11848 8628
rect 3148 8508 3200 8560
rect 3332 8508 3384 8560
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 3516 8440 3568 8492
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 3884 8440 3936 8492
rect 4436 8440 4488 8492
rect 4620 8440 4672 8492
rect 4988 8508 5040 8560
rect 5448 8508 5500 8560
rect 5632 8508 5684 8560
rect 2872 8347 2924 8356
rect 2872 8313 2881 8347
rect 2881 8313 2915 8347
rect 2915 8313 2924 8347
rect 2872 8304 2924 8313
rect 4344 8372 4396 8424
rect 5264 8440 5316 8492
rect 5908 8440 5960 8492
rect 9680 8508 9732 8560
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 6368 8372 6420 8424
rect 4436 8304 4488 8356
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 5632 8304 5684 8356
rect 6276 8304 6328 8356
rect 8484 8304 8536 8356
rect 10968 8440 11020 8492
rect 12624 8440 12676 8492
rect 13728 8440 13780 8492
rect 14372 8508 14424 8560
rect 14464 8440 14516 8492
rect 9772 8372 9824 8424
rect 13544 8372 13596 8424
rect 16396 8508 16448 8560
rect 15568 8440 15620 8492
rect 15752 8440 15804 8492
rect 18420 8576 18472 8628
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 16212 8372 16264 8424
rect 16948 8372 17000 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 1676 8236 1728 8288
rect 3516 8236 3568 8288
rect 4160 8236 4212 8288
rect 5264 8236 5316 8288
rect 5724 8236 5776 8288
rect 6460 8236 6512 8288
rect 8668 8236 8720 8288
rect 9036 8236 9088 8288
rect 9404 8236 9456 8288
rect 10324 8304 10376 8356
rect 11520 8304 11572 8356
rect 12072 8304 12124 8356
rect 12716 8304 12768 8356
rect 11244 8236 11296 8288
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 12256 8279 12308 8288
rect 12256 8245 12265 8279
rect 12265 8245 12299 8279
rect 12299 8245 12308 8279
rect 12256 8236 12308 8245
rect 13176 8236 13228 8288
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 13544 8236 13596 8288
rect 13636 8236 13688 8288
rect 16488 8304 16540 8356
rect 17316 8304 17368 8356
rect 17868 8372 17920 8424
rect 18144 8372 18196 8424
rect 18420 8415 18472 8424
rect 18420 8381 18429 8415
rect 18429 8381 18463 8415
rect 18463 8381 18472 8415
rect 18420 8372 18472 8381
rect 17960 8347 18012 8356
rect 17960 8313 17969 8347
rect 17969 8313 18003 8347
rect 18003 8313 18012 8347
rect 17960 8304 18012 8313
rect 14556 8236 14608 8288
rect 16672 8236 16724 8288
rect 17592 8279 17644 8288
rect 17592 8245 17601 8279
rect 17601 8245 17635 8279
rect 17635 8245 17644 8279
rect 17592 8236 17644 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 5724 8032 5776 8084
rect 5816 8032 5868 8084
rect 6276 8075 6328 8084
rect 6276 8041 6285 8075
rect 6285 8041 6319 8075
rect 6319 8041 6328 8075
rect 6276 8032 6328 8041
rect 1676 7964 1728 8016
rect 3424 8007 3476 8016
rect 2964 7896 3016 7948
rect 2320 7828 2372 7880
rect 3424 7973 3433 8007
rect 3433 7973 3467 8007
rect 3467 7973 3476 8007
rect 3424 7964 3476 7973
rect 6644 8032 6696 8084
rect 4620 7896 4672 7948
rect 5908 7896 5960 7948
rect 8024 8032 8076 8084
rect 8484 8032 8536 8084
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 4712 7828 4764 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 4160 7760 4212 7812
rect 5908 7760 5960 7812
rect 7104 7828 7156 7880
rect 8392 7964 8444 8016
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 9312 7964 9364 8016
rect 9404 7964 9456 8016
rect 11520 7964 11572 8016
rect 12532 8032 12584 8084
rect 13176 8032 13228 8084
rect 16488 8032 16540 8084
rect 16764 8032 16816 8084
rect 17224 8075 17276 8084
rect 17224 8041 17233 8075
rect 17233 8041 17267 8075
rect 17267 8041 17276 8075
rect 17224 8032 17276 8041
rect 13544 7964 13596 8016
rect 14464 7964 14516 8016
rect 17868 7964 17920 8016
rect 18604 7964 18656 8016
rect 8392 7828 8444 7880
rect 11060 7896 11112 7948
rect 15200 7896 15252 7948
rect 15476 7939 15528 7948
rect 15476 7905 15494 7939
rect 15494 7905 15528 7939
rect 15476 7896 15528 7905
rect 15660 7896 15712 7948
rect 17224 7896 17276 7948
rect 3792 7692 3844 7744
rect 4252 7692 4304 7744
rect 4620 7692 4672 7744
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 9772 7760 9824 7812
rect 11152 7760 11204 7812
rect 13544 7828 13596 7880
rect 13912 7871 13964 7880
rect 13912 7837 13921 7871
rect 13921 7837 13955 7871
rect 13955 7837 13964 7871
rect 13912 7828 13964 7837
rect 12624 7760 12676 7812
rect 9036 7692 9088 7744
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 11244 7735 11296 7744
rect 9128 7692 9180 7701
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 13452 7692 13504 7744
rect 13728 7692 13780 7744
rect 14464 7760 14516 7812
rect 17960 7803 18012 7812
rect 17960 7769 17969 7803
rect 17969 7769 18003 7803
rect 18003 7769 18012 7803
rect 17960 7760 18012 7769
rect 15016 7692 15068 7744
rect 18144 7735 18196 7744
rect 18144 7701 18153 7735
rect 18153 7701 18187 7735
rect 18187 7701 18196 7735
rect 18144 7692 18196 7701
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 2320 7488 2372 7540
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 5908 7488 5960 7540
rect 6460 7531 6512 7540
rect 6460 7497 6469 7531
rect 6469 7497 6503 7531
rect 6503 7497 6512 7531
rect 6460 7488 6512 7497
rect 6736 7488 6788 7540
rect 7472 7488 7524 7540
rect 8760 7488 8812 7540
rect 3056 7463 3108 7472
rect 3056 7429 3065 7463
rect 3065 7429 3099 7463
rect 3099 7429 3108 7463
rect 3056 7420 3108 7429
rect 2688 7352 2740 7404
rect 4988 7420 5040 7472
rect 6828 7420 6880 7472
rect 8484 7463 8536 7472
rect 4436 7352 4488 7404
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 1676 7284 1728 7336
rect 3516 7284 3568 7336
rect 3608 7284 3660 7336
rect 3792 7284 3844 7336
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 4528 7284 4580 7336
rect 6736 7352 6788 7404
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7840 7352 7892 7404
rect 6368 7284 6420 7336
rect 6644 7284 6696 7336
rect 2504 7216 2556 7268
rect 3240 7259 3292 7268
rect 3240 7225 3249 7259
rect 3249 7225 3283 7259
rect 3283 7225 3292 7259
rect 3240 7216 3292 7225
rect 7564 7216 7616 7268
rect 7656 7259 7708 7268
rect 7656 7225 7665 7259
rect 7665 7225 7699 7259
rect 7699 7225 7708 7259
rect 8484 7429 8493 7463
rect 8493 7429 8527 7463
rect 8527 7429 8536 7463
rect 8484 7420 8536 7429
rect 9772 7352 9824 7404
rect 11612 7352 11664 7404
rect 12256 7488 12308 7540
rect 12716 7488 12768 7540
rect 13912 7488 13964 7540
rect 15200 7488 15252 7540
rect 17132 7488 17184 7540
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 17868 7488 17920 7540
rect 12532 7420 12584 7472
rect 12716 7352 12768 7404
rect 13636 7352 13688 7404
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 8668 7284 8720 7336
rect 9312 7284 9364 7336
rect 13544 7327 13596 7336
rect 7656 7216 7708 7225
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 4160 7148 4212 7200
rect 4252 7148 4304 7200
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 6092 7148 6144 7200
rect 8116 7148 8168 7200
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 9496 7148 9548 7200
rect 10232 7216 10284 7268
rect 10968 7216 11020 7268
rect 11244 7216 11296 7268
rect 11336 7148 11388 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 12624 7216 12676 7268
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 13820 7284 13872 7336
rect 14464 7420 14516 7472
rect 16672 7420 16724 7472
rect 18144 7420 18196 7472
rect 15476 7352 15528 7404
rect 16580 7352 16632 7404
rect 18512 7395 18564 7404
rect 17224 7284 17276 7336
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 17868 7327 17920 7336
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 13176 7148 13228 7200
rect 13268 7148 13320 7200
rect 13544 7148 13596 7200
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 15752 7148 15804 7157
rect 16488 7216 16540 7268
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 1584 6944 1636 6996
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2044 6944 2096 6996
rect 2688 6944 2740 6996
rect 4252 6987 4304 6996
rect 4252 6953 4261 6987
rect 4261 6953 4295 6987
rect 4295 6953 4304 6987
rect 4252 6944 4304 6953
rect 4804 6944 4856 6996
rect 8392 6944 8444 6996
rect 10416 6944 10468 6996
rect 2412 6876 2464 6928
rect 4344 6919 4396 6928
rect 4344 6885 4353 6919
rect 4353 6885 4387 6919
rect 4387 6885 4396 6919
rect 4344 6876 4396 6885
rect 4988 6876 5040 6928
rect 5448 6876 5500 6928
rect 6460 6876 6512 6928
rect 6552 6876 6604 6928
rect 8116 6876 8168 6928
rect 8484 6876 8536 6928
rect 12256 6944 12308 6996
rect 13544 6944 13596 6996
rect 10968 6876 11020 6928
rect 11428 6919 11480 6928
rect 11428 6885 11437 6919
rect 11437 6885 11471 6919
rect 11471 6885 11480 6919
rect 11428 6876 11480 6885
rect 11704 6919 11756 6928
rect 11704 6885 11713 6919
rect 11713 6885 11747 6919
rect 11747 6885 11756 6919
rect 11704 6876 11756 6885
rect 12624 6876 12676 6928
rect 2044 6808 2096 6860
rect 3148 6808 3200 6860
rect 4436 6808 4488 6860
rect 5080 6851 5132 6860
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 5724 6808 5776 6860
rect 6736 6808 6788 6860
rect 3332 6672 3384 6724
rect 6644 6740 6696 6792
rect 5632 6715 5684 6724
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 5632 6681 5641 6715
rect 5641 6681 5675 6715
rect 5675 6681 5684 6715
rect 5632 6672 5684 6681
rect 6828 6672 6880 6724
rect 8024 6808 8076 6860
rect 9680 6808 9732 6860
rect 4344 6604 4396 6656
rect 5172 6604 5224 6656
rect 5816 6604 5868 6656
rect 9588 6740 9640 6792
rect 8760 6672 8812 6724
rect 10232 6672 10284 6724
rect 8484 6604 8536 6656
rect 9588 6604 9640 6656
rect 11152 6604 11204 6656
rect 11980 6740 12032 6792
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 12992 6851 13044 6860
rect 12992 6817 13001 6851
rect 13001 6817 13035 6851
rect 13035 6817 13044 6851
rect 12992 6808 13044 6817
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 14188 6808 14240 6860
rect 15752 6944 15804 6996
rect 17224 6987 17276 6996
rect 17224 6953 17233 6987
rect 17233 6953 17267 6987
rect 17267 6953 17276 6987
rect 17224 6944 17276 6953
rect 17500 6987 17552 6996
rect 17500 6953 17509 6987
rect 17509 6953 17543 6987
rect 17543 6953 17552 6987
rect 17500 6944 17552 6953
rect 17868 6944 17920 6996
rect 18052 6876 18104 6928
rect 18144 6851 18196 6860
rect 18144 6817 18153 6851
rect 18153 6817 18187 6851
rect 18187 6817 18196 6851
rect 18144 6808 18196 6817
rect 18328 6851 18380 6860
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 15016 6783 15068 6792
rect 13544 6672 13596 6724
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 15108 6672 15160 6724
rect 15568 6672 15620 6724
rect 15936 6715 15988 6724
rect 15936 6681 15945 6715
rect 15945 6681 15979 6715
rect 15979 6681 15988 6715
rect 15936 6672 15988 6681
rect 16488 6672 16540 6724
rect 17960 6672 18012 6724
rect 18512 6715 18564 6724
rect 18512 6681 18521 6715
rect 18521 6681 18555 6715
rect 18555 6681 18564 6715
rect 18512 6672 18564 6681
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 14832 6604 14884 6656
rect 16120 6604 16172 6656
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 2872 6332 2924 6384
rect 3516 6307 3568 6316
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 2688 6196 2740 6248
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 3608 6196 3660 6248
rect 4160 6196 4212 6248
rect 5816 6307 5868 6316
rect 4804 6196 4856 6248
rect 5172 6239 5224 6248
rect 5172 6205 5190 6239
rect 5190 6205 5224 6239
rect 5448 6239 5500 6248
rect 5172 6196 5224 6205
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 2412 6060 2464 6112
rect 4712 6128 4764 6180
rect 5540 6128 5592 6180
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 8392 6400 8444 6452
rect 8116 6332 8168 6384
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 8300 6196 8352 6248
rect 6828 6128 6880 6180
rect 3976 6060 4028 6112
rect 6184 6060 6236 6112
rect 6460 6060 6512 6112
rect 7932 6060 7984 6112
rect 9128 6128 9180 6180
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 8576 6060 8628 6112
rect 9496 6128 9548 6180
rect 11060 6400 11112 6452
rect 11152 6400 11204 6452
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 12992 6400 13044 6452
rect 13636 6443 13688 6452
rect 13636 6409 13645 6443
rect 13645 6409 13679 6443
rect 13679 6409 13688 6443
rect 13636 6400 13688 6409
rect 10140 6332 10192 6384
rect 10600 6332 10652 6384
rect 11520 6264 11572 6316
rect 11980 6264 12032 6316
rect 13544 6264 13596 6316
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 11796 6196 11848 6248
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 12164 6196 12216 6248
rect 9864 6060 9916 6112
rect 10968 6060 11020 6112
rect 12348 6103 12400 6112
rect 12348 6069 12357 6103
rect 12357 6069 12391 6103
rect 12391 6069 12400 6103
rect 12348 6060 12400 6069
rect 14924 6196 14976 6248
rect 16948 6400 17000 6452
rect 18328 6400 18380 6452
rect 15200 6196 15252 6248
rect 13176 6171 13228 6180
rect 13176 6137 13185 6171
rect 13185 6137 13219 6171
rect 13219 6137 13228 6171
rect 13176 6128 13228 6137
rect 14464 6128 14516 6180
rect 14832 6128 14884 6180
rect 18420 6196 18472 6248
rect 14556 6060 14608 6112
rect 14740 6060 14792 6112
rect 14924 6060 14976 6112
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 18512 6171 18564 6180
rect 18052 6103 18104 6112
rect 15476 6060 15528 6069
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 18512 6137 18521 6171
rect 18521 6137 18555 6171
rect 18555 6137 18564 6171
rect 18512 6128 18564 6137
rect 18420 6060 18472 6112
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 3792 5856 3844 5908
rect 4068 5856 4120 5908
rect 4344 5899 4396 5908
rect 4344 5865 4353 5899
rect 4353 5865 4387 5899
rect 4387 5865 4396 5899
rect 4344 5856 4396 5865
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 4896 5856 4948 5908
rect 5264 5856 5316 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 3976 5788 4028 5840
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 3240 5720 3292 5772
rect 3700 5720 3752 5772
rect 4344 5720 4396 5772
rect 8484 5856 8536 5908
rect 8116 5788 8168 5840
rect 9772 5856 9824 5908
rect 13544 5899 13596 5908
rect 9680 5788 9732 5840
rect 10140 5788 10192 5840
rect 11152 5788 11204 5840
rect 4896 5720 4948 5772
rect 5632 5720 5684 5772
rect 6828 5720 6880 5772
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 3056 5584 3108 5636
rect 4344 5584 4396 5636
rect 5172 5584 5224 5636
rect 7472 5720 7524 5772
rect 7840 5720 7892 5772
rect 9036 5720 9088 5772
rect 9404 5720 9456 5772
rect 10600 5720 10652 5772
rect 11060 5720 11112 5772
rect 11336 5720 11388 5772
rect 11980 5720 12032 5772
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 13820 5856 13872 5908
rect 14280 5856 14332 5908
rect 14832 5899 14884 5908
rect 14832 5865 14841 5899
rect 14841 5865 14875 5899
rect 14875 5865 14884 5899
rect 14832 5856 14884 5865
rect 15200 5856 15252 5908
rect 17316 5856 17368 5908
rect 18420 5856 18472 5908
rect 12532 5788 12584 5840
rect 12624 5788 12676 5840
rect 14004 5720 14056 5772
rect 14096 5720 14148 5772
rect 14832 5720 14884 5772
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 16764 5720 16816 5772
rect 18052 5788 18104 5840
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 9864 5652 9916 5704
rect 14464 5652 14516 5704
rect 15108 5652 15160 5704
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 3792 5516 3844 5568
rect 10324 5516 10376 5568
rect 10692 5516 10744 5568
rect 11888 5584 11940 5636
rect 12164 5584 12216 5636
rect 11336 5559 11388 5568
rect 11336 5525 11345 5559
rect 11345 5525 11379 5559
rect 11379 5525 11388 5559
rect 11336 5516 11388 5525
rect 11704 5516 11756 5568
rect 14832 5584 14884 5636
rect 18512 5627 18564 5636
rect 18512 5593 18521 5627
rect 18521 5593 18555 5627
rect 18555 5593 18564 5627
rect 18512 5584 18564 5593
rect 13636 5516 13688 5568
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 14464 5516 14516 5568
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 1584 5312 1636 5364
rect 2044 5312 2096 5364
rect 3700 5312 3752 5364
rect 5172 5312 5224 5364
rect 5448 5312 5500 5364
rect 6552 5355 6604 5364
rect 3608 5244 3660 5296
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 8392 5312 8444 5364
rect 9128 5312 9180 5364
rect 9772 5312 9824 5364
rect 2964 5176 3016 5228
rect 3516 5176 3568 5228
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 7656 5244 7708 5296
rect 9220 5244 9272 5296
rect 16580 5312 16632 5364
rect 3148 5108 3200 5160
rect 3792 5108 3844 5160
rect 4252 5108 4304 5160
rect 4528 5108 4580 5160
rect 5264 5108 5316 5160
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 5908 5108 5960 5160
rect 8300 5108 8352 5160
rect 8576 5176 8628 5228
rect 8760 5176 8812 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 13820 5219 13872 5228
rect 9220 5108 9272 5160
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 10876 5108 10928 5160
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 16212 5244 16264 5296
rect 15568 5219 15620 5228
rect 13820 5176 13872 5185
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 16488 5176 16540 5228
rect 2964 5040 3016 5092
rect 4712 5040 4764 5092
rect 2228 4972 2280 5024
rect 2780 4972 2832 5024
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 4068 4972 4120 5024
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 5356 4972 5408 5024
rect 13452 5040 13504 5092
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 7840 5015 7892 5024
rect 7840 4981 7849 5015
rect 7849 4981 7883 5015
rect 7883 4981 7892 5015
rect 7840 4972 7892 4981
rect 8116 4972 8168 5024
rect 8300 4972 8352 5024
rect 9036 4972 9088 5024
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 10508 4972 10560 5024
rect 10692 4972 10744 5024
rect 12348 4972 12400 5024
rect 12532 4972 12584 5024
rect 12624 4972 12676 5024
rect 14372 5108 14424 5160
rect 14464 5040 14516 5092
rect 14372 4972 14424 5024
rect 14740 4972 14792 5024
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 18052 5108 18104 5160
rect 15108 5040 15160 5092
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 4068 4768 4120 4820
rect 4252 4768 4304 4820
rect 1400 4743 1452 4752
rect 1400 4709 1409 4743
rect 1409 4709 1443 4743
rect 1443 4709 1452 4743
rect 1400 4700 1452 4709
rect 1952 4675 2004 4684
rect 1952 4641 1961 4675
rect 1961 4641 1995 4675
rect 1995 4641 2004 4675
rect 1952 4632 2004 4641
rect 3148 4700 3200 4752
rect 4804 4700 4856 4752
rect 5080 4700 5132 4752
rect 8116 4768 8168 4820
rect 3056 4632 3108 4684
rect 3884 4675 3936 4684
rect 3884 4641 3893 4675
rect 3893 4641 3927 4675
rect 3927 4641 3936 4675
rect 3884 4632 3936 4641
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6368 4632 6420 4684
rect 6828 4700 6880 4752
rect 9404 4768 9456 4820
rect 11980 4768 12032 4820
rect 12256 4768 12308 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 14832 4811 14884 4820
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 16120 4768 16172 4820
rect 10692 4700 10744 4752
rect 11336 4700 11388 4752
rect 7380 4632 7432 4684
rect 9220 4632 9272 4684
rect 9772 4632 9824 4684
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 5264 4564 5316 4616
rect 5540 4564 5592 4616
rect 7656 4564 7708 4616
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 8484 4564 8536 4616
rect 11428 4632 11480 4684
rect 11612 4675 11664 4684
rect 11612 4641 11621 4675
rect 11621 4641 11655 4675
rect 11655 4641 11664 4675
rect 11612 4632 11664 4641
rect 12072 4700 12124 4752
rect 17408 4743 17460 4752
rect 17408 4709 17417 4743
rect 17417 4709 17451 4743
rect 17451 4709 17460 4743
rect 17408 4700 17460 4709
rect 17592 4700 17644 4752
rect 18052 4700 18104 4752
rect 14464 4632 14516 4684
rect 18144 4675 18196 4684
rect 18144 4641 18153 4675
rect 18153 4641 18187 4675
rect 18187 4641 18196 4675
rect 18144 4632 18196 4641
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11704 4607 11756 4616
rect 11152 4564 11204 4573
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 12256 4564 12308 4616
rect 12348 4564 12400 4616
rect 13820 4564 13872 4616
rect 14280 4564 14332 4616
rect 15108 4564 15160 4616
rect 6552 4496 6604 4548
rect 6644 4539 6696 4548
rect 6644 4505 6653 4539
rect 6653 4505 6687 4539
rect 6687 4505 6696 4539
rect 6644 4496 6696 4505
rect 7472 4496 7524 4548
rect 9680 4496 9732 4548
rect 11612 4496 11664 4548
rect 18512 4539 18564 4548
rect 5356 4428 5408 4480
rect 5448 4428 5500 4480
rect 6276 4428 6328 4480
rect 6828 4428 6880 4480
rect 8300 4471 8352 4480
rect 8300 4437 8309 4471
rect 8309 4437 8343 4471
rect 8343 4437 8352 4471
rect 8300 4428 8352 4437
rect 8392 4428 8444 4480
rect 9036 4428 9088 4480
rect 10968 4428 11020 4480
rect 11336 4428 11388 4480
rect 12256 4471 12308 4480
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 12256 4428 12308 4437
rect 18512 4505 18521 4539
rect 18521 4505 18555 4539
rect 18555 4505 18564 4539
rect 18512 4496 18564 4505
rect 14004 4428 14056 4480
rect 15476 4428 15528 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 3792 4224 3844 4276
rect 4804 4224 4856 4276
rect 6368 4224 6420 4276
rect 7932 4224 7984 4276
rect 8668 4224 8720 4276
rect 9128 4267 9180 4276
rect 9128 4233 9137 4267
rect 9137 4233 9171 4267
rect 9171 4233 9180 4267
rect 9128 4224 9180 4233
rect 11244 4224 11296 4276
rect 5356 4156 5408 4208
rect 5264 4131 5316 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 4160 4020 4212 4072
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5448 4088 5500 4140
rect 5540 4063 5592 4072
rect 1584 3995 1636 4004
rect 1584 3961 1593 3995
rect 1593 3961 1627 3995
rect 1627 3961 1636 3995
rect 1584 3952 1636 3961
rect 2228 3952 2280 4004
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 2136 3884 2188 3936
rect 3424 3927 3476 3936
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 4712 3952 4764 4004
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 5724 4088 5776 4140
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 9588 4088 9640 4140
rect 10324 4088 10376 4140
rect 10876 4156 10928 4208
rect 13912 4224 13964 4276
rect 14464 4267 14516 4276
rect 14464 4233 14473 4267
rect 14473 4233 14507 4267
rect 14507 4233 14516 4267
rect 14464 4224 14516 4233
rect 15476 4267 15528 4276
rect 15476 4233 15485 4267
rect 15485 4233 15519 4267
rect 15519 4233 15528 4267
rect 15476 4224 15528 4233
rect 11152 4088 11204 4140
rect 11612 4088 11664 4140
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 10416 4063 10468 4072
rect 3424 3884 3476 3893
rect 4620 3884 4672 3936
rect 5724 3884 5776 3936
rect 8024 3995 8076 4004
rect 6460 3927 6512 3936
rect 6460 3893 6469 3927
rect 6469 3893 6503 3927
rect 6503 3893 6512 3927
rect 6460 3884 6512 3893
rect 6552 3884 6604 3936
rect 6736 3884 6788 3936
rect 8024 3961 8058 3995
rect 8058 3961 8076 3995
rect 8024 3952 8076 3961
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10416 4020 10468 4029
rect 11980 4063 12032 4072
rect 11980 4029 12014 4063
rect 12014 4029 12032 4063
rect 14004 4063 14056 4072
rect 11980 4020 12032 4029
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 15200 4088 15252 4140
rect 16580 4063 16632 4072
rect 11244 3952 11296 4004
rect 11888 3952 11940 4004
rect 12164 3952 12216 4004
rect 13728 3952 13780 4004
rect 16580 4029 16589 4063
rect 16589 4029 16623 4063
rect 16623 4029 16632 4063
rect 16580 4020 16632 4029
rect 17408 4020 17460 4072
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9588 3927 9640 3936
rect 9220 3884 9272 3893
rect 9588 3893 9597 3927
rect 9597 3893 9631 3927
rect 9631 3893 9640 3927
rect 9588 3884 9640 3893
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 11152 3884 11204 3936
rect 11428 3884 11480 3936
rect 11980 3884 12032 3936
rect 12348 3884 12400 3936
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 16856 3952 16908 4004
rect 16672 3884 16724 3936
rect 18144 3995 18196 4004
rect 18144 3961 18153 3995
rect 18153 3961 18187 3995
rect 18187 3961 18196 3995
rect 18144 3952 18196 3961
rect 18512 3995 18564 4004
rect 18512 3961 18521 3995
rect 18521 3961 18555 3995
rect 18555 3961 18564 3995
rect 18512 3952 18564 3961
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 3332 3723 3384 3732
rect 2596 3612 2648 3664
rect 2872 3655 2924 3664
rect 2872 3621 2881 3655
rect 2881 3621 2915 3655
rect 2915 3621 2924 3655
rect 2872 3612 2924 3621
rect 2964 3612 3016 3664
rect 2412 3544 2464 3596
rect 3332 3689 3341 3723
rect 3341 3689 3375 3723
rect 3375 3689 3384 3723
rect 3332 3680 3384 3689
rect 3240 3612 3292 3664
rect 4896 3680 4948 3732
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 3240 3476 3292 3528
rect 3700 3519 3752 3528
rect 3700 3485 3709 3519
rect 3709 3485 3743 3519
rect 3743 3485 3752 3519
rect 3700 3476 3752 3485
rect 4160 3612 4212 3664
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 5080 3544 5132 3596
rect 6644 3680 6696 3732
rect 7380 3680 7432 3732
rect 6092 3612 6144 3664
rect 8208 3680 8260 3732
rect 9036 3680 9088 3732
rect 7748 3612 7800 3664
rect 5356 3544 5408 3596
rect 6736 3544 6788 3596
rect 7564 3544 7616 3596
rect 1400 3340 1452 3392
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 3792 3408 3844 3460
rect 5172 3408 5224 3460
rect 6644 3476 6696 3528
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8944 3612 8996 3664
rect 9220 3680 9272 3732
rect 9680 3680 9732 3732
rect 10876 3723 10928 3732
rect 10048 3612 10100 3664
rect 10876 3689 10885 3723
rect 10885 3689 10919 3723
rect 10919 3689 10928 3723
rect 10876 3680 10928 3689
rect 11704 3680 11756 3732
rect 10692 3612 10744 3664
rect 13176 3680 13228 3732
rect 13912 3723 13964 3732
rect 12072 3612 12124 3664
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 15108 3680 15160 3732
rect 10508 3544 10560 3596
rect 10876 3544 10928 3596
rect 11336 3544 11388 3596
rect 11888 3544 11940 3596
rect 12348 3587 12400 3596
rect 12348 3553 12371 3587
rect 12371 3553 12400 3587
rect 12348 3544 12400 3553
rect 13820 3612 13872 3664
rect 16396 3655 16448 3664
rect 16396 3621 16405 3655
rect 16405 3621 16439 3655
rect 16439 3621 16448 3655
rect 16396 3612 16448 3621
rect 17776 3612 17828 3664
rect 8024 3476 8076 3485
rect 9496 3476 9548 3528
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 7748 3408 7800 3460
rect 9312 3408 9364 3460
rect 9404 3408 9456 3460
rect 11612 3476 11664 3528
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 4620 3383 4672 3392
rect 4620 3349 4629 3383
rect 4629 3349 4663 3383
rect 4663 3349 4672 3383
rect 4620 3340 4672 3349
rect 4712 3340 4764 3392
rect 5448 3340 5500 3392
rect 6184 3340 6236 3392
rect 6644 3383 6696 3392
rect 6644 3349 6653 3383
rect 6653 3349 6687 3383
rect 6687 3349 6696 3383
rect 6644 3340 6696 3349
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 7196 3340 7248 3392
rect 8668 3340 8720 3392
rect 8944 3340 8996 3392
rect 9680 3340 9732 3392
rect 10876 3408 10928 3460
rect 10968 3408 11020 3460
rect 12348 3340 12400 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 16764 3408 16816 3460
rect 17868 3476 17920 3528
rect 18144 3451 18196 3460
rect 18144 3417 18153 3451
rect 18153 3417 18187 3451
rect 18187 3417 18196 3451
rect 18144 3408 18196 3417
rect 16856 3383 16908 3392
rect 16856 3349 16865 3383
rect 16865 3349 16899 3383
rect 16899 3349 16908 3383
rect 16856 3340 16908 3349
rect 17316 3340 17368 3392
rect 18328 3340 18380 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 1584 3136 1636 3188
rect 3792 3136 3844 3188
rect 4252 3136 4304 3188
rect 4528 3136 4580 3188
rect 6000 3136 6052 3188
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 3424 3000 3476 3052
rect 4896 3000 4948 3052
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 3700 2932 3752 2984
rect 4712 2932 4764 2984
rect 4804 2932 4856 2984
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 5724 3000 5776 3052
rect 6276 3000 6328 3052
rect 8024 3136 8076 3188
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 10416 3136 10468 3188
rect 11060 3136 11112 3188
rect 11980 3136 12032 3188
rect 12072 3136 12124 3188
rect 13820 3136 13872 3188
rect 14832 3136 14884 3188
rect 15568 3179 15620 3188
rect 15568 3145 15577 3179
rect 15577 3145 15611 3179
rect 15611 3145 15620 3179
rect 15568 3136 15620 3145
rect 11888 3068 11940 3120
rect 5816 2975 5868 2984
rect 5816 2941 5825 2975
rect 5825 2941 5859 2975
rect 5859 2941 5868 2975
rect 5816 2932 5868 2941
rect 6184 2932 6236 2984
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 388 2864 440 2916
rect 1768 2907 1820 2916
rect 1768 2873 1777 2907
rect 1777 2873 1811 2907
rect 1811 2873 1820 2907
rect 1768 2864 1820 2873
rect 2136 2864 2188 2916
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 2780 2796 2832 2848
rect 3240 2796 3292 2848
rect 4528 2796 4580 2848
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 4896 2796 4948 2848
rect 5356 2796 5408 2848
rect 6644 2864 6696 2916
rect 7656 2864 7708 2916
rect 8852 2932 8904 2984
rect 10692 3000 10744 3052
rect 11060 3000 11112 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 12808 3068 12860 3120
rect 13176 3111 13228 3120
rect 13176 3077 13185 3111
rect 13185 3077 13219 3111
rect 13219 3077 13228 3111
rect 13176 3068 13228 3077
rect 13268 3068 13320 3120
rect 16856 3068 16908 3120
rect 17776 3111 17828 3120
rect 12164 3000 12216 3052
rect 9864 2864 9916 2916
rect 10324 2864 10376 2916
rect 12256 2932 12308 2984
rect 12624 2932 12676 2984
rect 13176 2932 13228 2984
rect 13636 2932 13688 2984
rect 16304 2975 16356 2984
rect 16304 2941 16313 2975
rect 16313 2941 16347 2975
rect 16347 2941 16356 2975
rect 16304 2932 16356 2941
rect 17040 2932 17092 2984
rect 17776 3077 17785 3111
rect 17785 3077 17819 3111
rect 17819 3077 17828 3111
rect 17776 3068 17828 3077
rect 17316 3000 17368 3052
rect 17684 3000 17736 3052
rect 6000 2796 6052 2848
rect 6276 2796 6328 2848
rect 8300 2839 8352 2848
rect 8300 2805 8309 2839
rect 8309 2805 8343 2839
rect 8343 2805 8352 2839
rect 8300 2796 8352 2805
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 10140 2839 10192 2848
rect 10140 2805 10149 2839
rect 10149 2805 10183 2839
rect 10183 2805 10192 2839
rect 10140 2796 10192 2805
rect 10416 2796 10468 2848
rect 11888 2864 11940 2916
rect 12164 2864 12216 2916
rect 12348 2796 12400 2848
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12808 2864 12860 2916
rect 15844 2864 15896 2916
rect 17500 2864 17552 2916
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 12440 2796 12492 2805
rect 15752 2839 15804 2848
rect 15752 2805 15761 2839
rect 15761 2805 15795 2839
rect 15795 2805 15804 2839
rect 15752 2796 15804 2805
rect 16120 2839 16172 2848
rect 16120 2805 16129 2839
rect 16129 2805 16163 2839
rect 16163 2805 16172 2839
rect 16120 2796 16172 2805
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 16948 2796 17000 2805
rect 17224 2796 17276 2848
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 17408 2796 17460 2805
rect 17592 2796 17644 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 4804 2592 4856 2644
rect 6460 2592 6512 2644
rect 1216 2524 1268 2576
rect 2320 2567 2372 2576
rect 2320 2533 2329 2567
rect 2329 2533 2363 2567
rect 2363 2533 2372 2567
rect 2320 2524 2372 2533
rect 4620 2524 4672 2576
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 3516 2499 3568 2508
rect 1952 2388 2004 2440
rect 3516 2465 3525 2499
rect 3525 2465 3559 2499
rect 3559 2465 3568 2499
rect 3516 2456 3568 2465
rect 6276 2524 6328 2576
rect 6368 2524 6420 2576
rect 8852 2592 8904 2644
rect 9036 2592 9088 2644
rect 9864 2635 9916 2644
rect 9864 2601 9873 2635
rect 9873 2601 9907 2635
rect 9907 2601 9916 2635
rect 9864 2592 9916 2601
rect 10140 2592 10192 2644
rect 10416 2592 10468 2644
rect 11152 2592 11204 2644
rect 11704 2635 11756 2644
rect 7472 2524 7524 2576
rect 5080 2499 5132 2508
rect 2136 2320 2188 2372
rect 3056 2363 3108 2372
rect 3056 2329 3065 2363
rect 3065 2329 3099 2363
rect 3099 2329 3108 2363
rect 3056 2320 3108 2329
rect 2044 2252 2096 2304
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 3792 2320 3844 2372
rect 4436 2388 4488 2440
rect 5080 2465 5089 2499
rect 5089 2465 5123 2499
rect 5123 2465 5132 2499
rect 5080 2456 5132 2465
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 8576 2567 8628 2576
rect 8576 2533 8585 2567
rect 8585 2533 8619 2567
rect 8619 2533 8628 2567
rect 8576 2524 8628 2533
rect 8668 2524 8720 2576
rect 9312 2524 9364 2576
rect 11336 2524 11388 2576
rect 11704 2601 11713 2635
rect 11713 2601 11747 2635
rect 11747 2601 11756 2635
rect 11704 2592 11756 2601
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 12440 2592 12492 2644
rect 15660 2635 15712 2644
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 17500 2592 17552 2644
rect 15568 2524 15620 2576
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 6644 2388 6696 2440
rect 6736 2388 6788 2440
rect 8484 2388 8536 2440
rect 10232 2388 10284 2440
rect 11060 2456 11112 2508
rect 11520 2499 11572 2508
rect 11520 2465 11529 2499
rect 11529 2465 11563 2499
rect 11563 2465 11572 2499
rect 11520 2456 11572 2465
rect 11704 2456 11756 2508
rect 13360 2456 13412 2508
rect 14648 2456 14700 2508
rect 15384 2499 15436 2508
rect 15384 2465 15393 2499
rect 15393 2465 15427 2499
rect 15427 2465 15436 2499
rect 15384 2456 15436 2465
rect 15660 2456 15712 2508
rect 15844 2456 15896 2508
rect 16948 2524 17000 2576
rect 17408 2524 17460 2576
rect 18236 2524 18288 2576
rect 16580 2456 16632 2508
rect 17040 2456 17092 2508
rect 4896 2320 4948 2372
rect 7564 2320 7616 2372
rect 5080 2252 5132 2304
rect 6276 2295 6328 2304
rect 6276 2261 6285 2295
rect 6285 2261 6319 2295
rect 6319 2261 6328 2295
rect 6276 2252 6328 2261
rect 6368 2252 6420 2304
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 11244 2320 11296 2372
rect 13084 2363 13136 2372
rect 13084 2329 13093 2363
rect 13093 2329 13127 2363
rect 13127 2329 13136 2363
rect 13084 2320 13136 2329
rect 13912 2363 13964 2372
rect 13912 2329 13921 2363
rect 13921 2329 13955 2363
rect 13955 2329 13964 2363
rect 13912 2320 13964 2329
rect 14832 2363 14884 2372
rect 14832 2329 14841 2363
rect 14841 2329 14875 2363
rect 14875 2329 14884 2363
rect 14832 2320 14884 2329
rect 15292 2320 15344 2372
rect 16580 2363 16632 2372
rect 16580 2329 16589 2363
rect 16589 2329 16623 2363
rect 16623 2329 16632 2363
rect 16580 2320 16632 2329
rect 18512 2363 18564 2372
rect 18512 2329 18521 2363
rect 18521 2329 18555 2363
rect 18555 2329 18564 2363
rect 18512 2320 18564 2329
rect 11428 2252 11480 2304
rect 12440 2252 12492 2304
rect 16672 2252 16724 2304
rect 17500 2252 17552 2304
rect 17776 2252 17828 2304
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 3516 2048 3568 2100
rect 8300 2048 8352 2100
rect 2964 1980 3016 2032
rect 6920 1980 6972 2032
rect 2688 1912 2740 1964
rect 7288 1912 7340 1964
rect 1952 1844 2004 1896
rect 5908 1844 5960 1896
rect 6276 1844 6328 1896
rect 7656 1844 7708 1896
rect 5080 1776 5132 1828
rect 10508 1776 10560 1828
rect 9680 1708 9732 1760
rect 19432 1708 19484 1760
rect 17224 1504 17276 1556
rect 17592 1504 17644 1556
<< metal2 >>
rect 1122 16400 1178 17200
rect 3054 16416 3110 16425
rect 1136 13802 1164 16400
rect 3330 16400 3386 17200
rect 3514 16824 3570 16833
rect 3514 16759 3570 16768
rect 3054 16351 3110 16360
rect 2962 16008 3018 16017
rect 2962 15943 3018 15952
rect 2502 15600 2558 15609
rect 2502 15535 2558 15544
rect 2226 15192 2282 15201
rect 2226 15127 2282 15136
rect 1858 14784 1914 14793
rect 1858 14719 1914 14728
rect 1872 14550 1900 14719
rect 2240 14550 2268 15127
rect 2320 14884 2372 14890
rect 2320 14826 2372 14832
rect 1860 14544 1912 14550
rect 2228 14544 2280 14550
rect 1860 14486 1912 14492
rect 2226 14512 2228 14521
rect 2280 14512 2282 14521
rect 1492 14476 1544 14482
rect 2226 14447 2282 14456
rect 1492 14418 1544 14424
rect 1504 14385 1532 14418
rect 1490 14376 1546 14385
rect 1490 14311 1546 14320
rect 1676 14340 1728 14346
rect 1504 14074 1532 14311
rect 1676 14282 1728 14288
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1688 13977 1716 14282
rect 1490 13968 1546 13977
rect 1490 13903 1546 13912
rect 1674 13968 1730 13977
rect 1674 13903 1730 13912
rect 1504 13870 1532 13903
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1124 13796 1176 13802
rect 1124 13738 1176 13744
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 1858 13560 1914 13569
rect 1964 13530 1992 13738
rect 2332 13734 2360 14826
rect 2516 14482 2544 15535
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 1858 13495 1914 13504
rect 1952 13524 2004 13530
rect 1872 13462 1900 13495
rect 1952 13466 2004 13472
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1504 13161 1532 13330
rect 1490 13152 1546 13161
rect 1490 13087 1546 13096
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12306 1440 12786
rect 1858 12744 1914 12753
rect 1492 12708 1544 12714
rect 1858 12679 1860 12688
rect 1492 12650 1544 12656
rect 1912 12679 1914 12688
rect 1860 12650 1912 12656
rect 1504 12345 1532 12650
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 1490 12336 1546 12345
rect 1400 12300 1452 12306
rect 2240 12306 2268 12582
rect 1490 12271 1546 12280
rect 2228 12300 2280 12306
rect 1400 12242 1452 12248
rect 2228 12242 2280 12248
rect 1412 11393 1440 12242
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1398 11384 1454 11393
rect 1596 11354 1624 12038
rect 1964 11898 1992 12038
rect 2240 11937 2268 12242
rect 2226 11928 2282 11937
rect 1952 11892 2004 11898
rect 2226 11863 2282 11872
rect 1952 11834 2004 11840
rect 1768 11620 1820 11626
rect 1768 11562 1820 11568
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1398 11319 1454 11328
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1688 10713 1716 11494
rect 1674 10704 1730 10713
rect 1674 10639 1730 10648
rect 1780 10169 1808 11562
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 10810 1900 11154
rect 2056 10985 2084 11562
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2042 10976 2098 10985
rect 2042 10911 2098 10920
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1860 10464 1912 10470
rect 1858 10432 1860 10441
rect 2136 10464 2188 10470
rect 1912 10432 1914 10441
rect 2136 10406 2188 10412
rect 1858 10367 1914 10376
rect 1766 10160 1822 10169
rect 1766 10095 1822 10104
rect 2148 9042 2176 10406
rect 2240 9518 2268 11018
rect 2332 10810 2360 11086
rect 2516 11014 2544 14282
rect 2608 13734 2636 14554
rect 2976 14482 3004 15943
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 13938 2728 14350
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2884 13870 2912 14418
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 3068 13530 3096 16351
rect 3344 14498 3372 16400
rect 3344 14482 3464 14498
rect 3344 14476 3476 14482
rect 3344 14470 3424 14476
rect 3424 14418 3476 14424
rect 3528 14414 3556 16759
rect 5538 16400 5594 17200
rect 7746 16400 7802 17200
rect 9954 16400 10010 17200
rect 12162 16400 12218 17200
rect 14370 16400 14426 17200
rect 16486 16824 16542 16833
rect 16486 16759 16542 16768
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14618 4108 14758
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 5552 14550 5580 16400
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 7760 14618 7788 16400
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 9968 14550 9996 16400
rect 12176 14550 12204 16400
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 3608 14544 3660 14550
rect 3606 14512 3608 14521
rect 5540 14544 5592 14550
rect 3660 14512 3662 14521
rect 5540 14486 5592 14492
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 3606 14447 3662 14456
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3252 14074 3280 14350
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3344 13530 3372 14214
rect 3528 14074 3556 14350
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12102 2912 12718
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2424 10130 2452 10950
rect 2608 10606 2636 11494
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2792 10198 2820 11698
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 10577 2912 11494
rect 3068 10577 3096 13262
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3252 11694 3280 13194
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3344 11558 3372 13330
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3436 11336 3464 13126
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3528 12442 3556 12650
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3344 11308 3464 11336
rect 2870 10568 2926 10577
rect 2870 10503 2926 10512
rect 3054 10568 3110 10577
rect 3344 10554 3372 11308
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3436 10674 3464 11154
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3344 10526 3464 10554
rect 3054 10503 3110 10512
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2318 10024 2374 10033
rect 2318 9959 2374 9968
rect 2332 9926 2360 9959
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2332 9042 2360 9862
rect 2792 9654 2820 9862
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 1504 8945 1532 8978
rect 1490 8936 1546 8945
rect 1412 8894 1490 8922
rect 1412 7546 1440 8894
rect 1490 8871 1546 8880
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1676 8288 1728 8294
rect 1676 8230 1728 8236
rect 1688 8022 1716 8230
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1504 7313 1532 7686
rect 1688 7342 1716 7958
rect 1584 7336 1636 7342
rect 1490 7304 1546 7313
rect 1584 7278 1636 7284
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1490 7239 1546 7248
rect 1596 7002 1624 7278
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1766 6896 1822 6905
rect 1766 6831 1768 6840
rect 1820 6831 1822 6840
rect 1768 6802 1820 6808
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6497 1532 6598
rect 1490 6488 1546 6497
rect 1490 6423 1546 6432
rect 1492 6112 1544 6118
rect 1860 6112 1912 6118
rect 1492 6054 1544 6060
rect 1858 6080 1860 6089
rect 1912 6080 1914 6089
rect 1504 5545 1532 6054
rect 1858 6015 1914 6024
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1490 5536 1546 5545
rect 1490 5471 1546 5480
rect 1596 5370 1624 5646
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1872 4826 1900 5063
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1400 4752 1452 4758
rect 1398 4720 1400 4729
rect 1452 4720 1454 4729
rect 1964 4690 1992 8774
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2042 7032 2098 7041
rect 2042 6967 2044 6976
rect 2096 6967 2098 6976
rect 2044 6938 2096 6944
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 5370 2084 6802
rect 2148 6254 2176 8570
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2332 7546 2360 7822
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2332 7018 2360 7482
rect 2516 7274 2544 7686
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2332 6990 2452 7018
rect 2424 6934 2452 6990
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2136 6248 2188 6254
rect 2134 6216 2136 6225
rect 2188 6216 2190 6225
rect 2134 6151 2190 6160
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 1398 4655 1454 4664
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 2240 4622 2268 4966
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1584 4004 1636 4010
rect 1584 3946 1636 3952
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 388 2916 440 2922
rect 388 2858 440 2864
rect 400 800 428 2858
rect 1216 2576 1268 2582
rect 1216 2518 1268 2524
rect 1228 800 1256 2518
rect 1412 1057 1440 3334
rect 1504 2281 1532 3878
rect 1596 3194 1624 3946
rect 1780 3233 1808 4014
rect 2240 4010 2268 4558
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1766 3224 1822 3233
rect 1584 3188 1636 3194
rect 1766 3159 1822 3168
rect 1584 3130 1636 3136
rect 1584 2984 1636 2990
rect 1582 2952 1584 2961
rect 1636 2952 1638 2961
rect 1582 2887 1638 2896
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 1490 2272 1546 2281
rect 1490 2207 1546 2216
rect 1398 1048 1454 1057
rect 1398 983 1454 992
rect 386 0 442 800
rect 1214 0 1270 800
rect 1780 649 1808 2858
rect 1872 1873 1900 3334
rect 2148 2922 2176 3878
rect 2424 3602 2452 6054
rect 2608 3777 2636 9318
rect 2792 9178 2820 9590
rect 2884 9450 2912 10503
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9586 3004 9862
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8498 2820 8978
rect 3068 8634 3096 10503
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3160 9518 3188 10406
rect 3344 10266 3372 10406
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 9353 3188 9454
rect 3146 9344 3202 9353
rect 3146 9279 3202 9288
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3148 8560 3200 8566
rect 3054 8528 3110 8537
rect 2780 8492 2832 8498
rect 3148 8502 3200 8508
rect 3054 8463 3110 8472
rect 2780 8434 2832 8440
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 7721 2912 8298
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2870 7712 2926 7721
rect 2870 7647 2926 7656
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2700 7002 2728 7346
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2976 6458 3004 7890
rect 3068 7478 3096 8463
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 3160 6866 3188 8502
rect 3252 7274 3280 9862
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3344 9450 3372 9687
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8566 3372 8774
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3436 8242 3464 10526
rect 3528 9568 3556 12242
rect 3620 11898 3648 14282
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 5630 13968 5686 13977
rect 5630 13903 5632 13912
rect 5684 13903 5686 13912
rect 5632 13874 5684 13880
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3712 12306 3740 13466
rect 5092 13394 5120 13670
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3884 12232 3936 12238
rect 3882 12200 3884 12209
rect 3936 12200 3938 12209
rect 3882 12135 3938 12144
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3620 10606 3648 11834
rect 3712 11150 3740 12038
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 4264 11762 4292 12038
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4356 11626 4384 13126
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4448 11830 4476 12582
rect 4632 12434 4660 13194
rect 4724 12986 4752 13330
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4908 12442 4936 13262
rect 4540 12406 4660 12434
rect 4896 12436 4948 12442
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3606 10296 3662 10305
rect 3606 10231 3662 10240
rect 3620 9722 3648 10231
rect 3712 10033 3740 11086
rect 3804 10606 3832 11494
rect 4068 11348 4120 11354
rect 4172 11336 4200 11562
rect 4252 11348 4304 11354
rect 4172 11308 4252 11336
rect 4068 11290 4120 11296
rect 4252 11290 4304 11296
rect 4080 11234 4108 11290
rect 4448 11286 4476 11766
rect 4436 11280 4488 11286
rect 4080 11206 4384 11234
rect 4436 11222 4488 11228
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 10266 3832 10406
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 4066 10160 4122 10169
rect 4066 10095 4068 10104
rect 4120 10095 4122 10104
rect 4068 10066 4120 10072
rect 3698 10024 3754 10033
rect 3698 9959 3754 9968
rect 4158 10024 4214 10033
rect 4158 9959 4160 9968
rect 4212 9959 4214 9968
rect 4160 9930 4212 9936
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3528 9540 3648 9568
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3528 8498 3556 9386
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3344 8214 3464 8242
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3344 6882 3372 8214
rect 3422 8120 3478 8129
rect 3422 8055 3478 8064
rect 3436 8022 3464 8055
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3528 7868 3556 8230
rect 3436 7840 3556 7868
rect 3436 7313 3464 7840
rect 3514 7712 3570 7721
rect 3514 7647 3570 7656
rect 3528 7546 3556 7647
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3620 7342 3648 9540
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3712 8498 3740 9046
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3804 7750 3832 9658
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3896 9178 3924 9590
rect 3988 9518 4016 9590
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3988 9042 4016 9318
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3882 8528 3938 8537
rect 3882 8463 3884 8472
rect 3936 8463 3938 8472
rect 3884 8434 3936 8440
rect 3896 7857 3924 8434
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3882 7848 3938 7857
rect 4172 7818 4200 8230
rect 3882 7783 3938 7792
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4264 7750 4292 10950
rect 4356 10248 4384 11206
rect 4356 10220 4476 10248
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4356 9722 4384 10066
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4356 8430 4384 9046
rect 4448 8498 4476 10220
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 3698 7440 3754 7449
rect 3698 7375 3754 7384
rect 3516 7336 3568 7342
rect 3422 7304 3478 7313
rect 3516 7278 3568 7284
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3422 7239 3478 7248
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3252 6854 3372 6882
rect 3146 6760 3202 6769
rect 3146 6695 3202 6704
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2700 4593 2728 6190
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2884 4978 2912 6326
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5234 3004 5510
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2976 5098 3004 5170
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2686 4584 2742 4593
rect 2686 4519 2742 4528
rect 2594 3768 2650 3777
rect 2594 3703 2650 3712
rect 2596 3664 2648 3670
rect 2792 3618 2820 4966
rect 2884 4950 3004 4978
rect 2870 3904 2926 3913
rect 2870 3839 2926 3848
rect 2884 3670 2912 3839
rect 2976 3670 3004 4950
rect 3068 4690 3096 5578
rect 3160 5166 3188 6695
rect 3252 5778 3280 6854
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3344 6254 3372 6666
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3252 5681 3280 5714
rect 3238 5672 3294 5681
rect 3238 5607 3294 5616
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3160 4758 3188 4966
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 3252 3670 3280 5510
rect 3436 4468 3464 7239
rect 3528 6322 3556 7278
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3620 6254 3648 7142
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3712 5778 3740 7375
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 4068 7336 4120 7342
rect 4264 7290 4292 7686
rect 4068 7278 4120 7284
rect 3804 5914 3832 7278
rect 4080 6905 4108 7278
rect 4172 7262 4292 7290
rect 4172 7206 4200 7262
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 7002 4292 7142
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4356 6934 4384 8366
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4448 7886 4476 8298
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7410 4476 7822
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4344 6928 4396 6934
rect 4066 6896 4122 6905
rect 4344 6870 4396 6876
rect 4448 6866 4476 7346
rect 4540 7342 4568 12406
rect 4896 12378 4948 12384
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4618 12200 4674 12209
rect 4618 12135 4674 12144
rect 4632 10441 4660 12135
rect 4724 11898 4752 12242
rect 4908 12238 4936 12378
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 5000 12170 5028 13330
rect 5092 12850 5120 13330
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5092 12442 5120 12786
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4804 11688 4856 11694
rect 5184 11642 5212 13670
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 4804 11630 4856 11636
rect 4816 11558 4844 11630
rect 5092 11614 5212 11642
rect 5092 11558 5120 11614
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 4618 10432 4674 10441
rect 4618 10367 4674 10376
rect 4632 9518 4660 10367
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 9178 4752 9318
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4724 9042 4752 9114
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4632 8922 4660 8978
rect 4710 8936 4766 8945
rect 4632 8894 4710 8922
rect 4710 8871 4766 8880
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 7993 4660 8434
rect 4724 8362 4752 8871
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4618 7984 4674 7993
rect 4618 7919 4620 7928
rect 4672 7919 4674 7928
rect 4620 7890 4672 7896
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4066 6831 4122 6840
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3988 5846 4016 6054
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3792 5568 3844 5574
rect 4080 5556 4108 5850
rect 4172 5817 4200 6190
rect 4356 5914 4384 6598
rect 4434 6216 4490 6225
rect 4434 6151 4490 6160
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4158 5808 4214 5817
rect 4158 5743 4214 5752
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5642 4384 5714
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4080 5528 4292 5556
rect 3792 5510 3844 5516
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3528 4622 3556 5170
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3436 4440 3556 4468
rect 3330 4312 3386 4321
rect 3330 4247 3386 4256
rect 3344 3738 3372 4247
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 2648 3612 2820 3618
rect 2596 3606 2820 3612
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 2412 3596 2464 3602
rect 2608 3590 2820 3606
rect 2412 3538 2464 3544
rect 2504 3528 2556 3534
rect 2502 3496 2504 3505
rect 3240 3528 3292 3534
rect 2556 3496 2558 3505
rect 3240 3470 3292 3476
rect 2502 3431 2558 3440
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3097 2268 3334
rect 2226 3088 2282 3097
rect 2226 3023 2282 3032
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 3252 2854 3280 3470
rect 3436 3058 3464 3878
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3528 2990 3556 4440
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 2228 2848 2280 2854
rect 2780 2848 2832 2854
rect 2228 2790 2280 2796
rect 2318 2816 2374 2825
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1964 1902 1992 2382
rect 2056 2310 2084 2450
rect 2136 2372 2188 2378
rect 2136 2314 2188 2320
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 1952 1896 2004 1902
rect 1858 1864 1914 1873
rect 1952 1838 2004 1844
rect 1858 1799 1914 1808
rect 2148 800 2176 2314
rect 2240 1465 2268 2790
rect 2780 2790 2832 2796
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 2318 2751 2374 2760
rect 2332 2582 2360 2751
rect 2792 2689 2820 2790
rect 3620 2774 3648 5238
rect 3712 4672 3740 5306
rect 3804 5166 3832 5510
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4264 5166 4292 5528
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4826 4108 4966
rect 4264 4826 4292 5102
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3882 4720 3938 4729
rect 3712 4664 3882 4672
rect 3712 4644 3884 4664
rect 3804 4282 3832 4644
rect 3936 4655 3938 4664
rect 3884 4626 3936 4632
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 3698 3904 3754 3913
rect 3698 3839 3754 3848
rect 3712 3534 3740 3839
rect 4172 3670 4200 4014
rect 4356 3913 4384 5578
rect 4448 5234 4476 6151
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4540 5166 4568 5646
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4632 4978 4660 7686
rect 4724 6186 4752 7822
rect 4816 7206 4844 11494
rect 5184 11354 5212 11494
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 4908 9625 4936 11290
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10538 5120 10950
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10062 5120 10474
rect 5172 10192 5224 10198
rect 5276 10180 5304 13126
rect 5920 12850 5948 13126
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5552 12238 5580 12786
rect 6380 12714 6408 13398
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6656 12986 6684 13330
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11898 5488 12038
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5552 11762 5580 12174
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5736 11286 5764 12582
rect 5828 12434 5856 12650
rect 5828 12406 5948 12434
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5368 10198 5396 10746
rect 5224 10152 5304 10180
rect 5356 10192 5408 10198
rect 5172 10134 5224 10140
rect 5356 10134 5408 10140
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9674 5120 9998
rect 5184 9926 5212 10134
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5552 9738 5580 11222
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 10305 5672 11086
rect 5722 10704 5778 10713
rect 5722 10639 5778 10648
rect 5630 10296 5686 10305
rect 5630 10231 5686 10240
rect 5736 10180 5764 10639
rect 5828 10305 5856 12038
rect 5814 10296 5870 10305
rect 5814 10231 5870 10240
rect 5736 10152 5856 10180
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5000 9646 5120 9674
rect 5184 9710 5580 9738
rect 5184 9654 5212 9710
rect 5172 9648 5224 9654
rect 4894 9616 4950 9625
rect 5000 9586 5028 9646
rect 5172 9590 5224 9596
rect 5540 9648 5592 9654
rect 5644 9636 5672 10066
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5736 9654 5764 9998
rect 5592 9608 5672 9636
rect 5724 9648 5776 9654
rect 5540 9590 5592 9596
rect 5724 9590 5776 9596
rect 4894 9551 4950 9560
rect 4988 9580 5040 9586
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 7002 4844 7142
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4724 5098 4752 5850
rect 4816 5273 4844 6190
rect 4908 5914 4936 9551
rect 4988 9522 5040 9528
rect 5000 9353 5028 9522
rect 5828 9518 5856 10152
rect 5816 9512 5868 9518
rect 5736 9460 5816 9466
rect 5920 9489 5948 12406
rect 6182 12200 6238 12209
rect 6182 12135 6184 12144
rect 6236 12135 6238 12144
rect 6184 12106 6236 12112
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11694 6040 12038
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 10266 6040 10406
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6104 10010 6132 11154
rect 6196 11014 6224 12106
rect 6380 11830 6408 12650
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6368 11688 6420 11694
rect 6564 11665 6592 12582
rect 6656 12238 6684 12922
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6644 12232 6696 12238
rect 6748 12209 6776 12378
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 6644 12174 6696 12180
rect 6734 12200 6790 12209
rect 6656 11762 6684 12174
rect 6734 12135 6790 12144
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6368 11630 6420 11636
rect 6550 11656 6606 11665
rect 6184 11008 6236 11014
rect 6380 10996 6408 11630
rect 6550 11591 6606 11600
rect 6564 11218 6592 11591
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6656 11150 6684 11698
rect 6460 11144 6512 11150
rect 6458 11112 6460 11121
rect 6644 11144 6696 11150
rect 6512 11112 6514 11121
rect 6514 11070 6592 11098
rect 6644 11086 6696 11092
rect 6458 11047 6514 11056
rect 6380 10968 6500 10996
rect 6184 10950 6236 10956
rect 6274 10704 6330 10713
rect 6274 10639 6330 10648
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6012 9982 6132 10010
rect 5736 9454 5868 9460
rect 5906 9480 5962 9489
rect 5736 9438 5856 9454
rect 5080 9376 5132 9382
rect 4986 9344 5042 9353
rect 5080 9318 5132 9324
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 4986 9279 5042 9288
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5000 7478 5028 8502
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4802 5264 4858 5273
rect 4802 5199 4858 5208
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4804 5024 4856 5030
rect 4632 4950 4752 4978
rect 4804 4966 4856 4972
rect 4618 4584 4674 4593
rect 4618 4519 4674 4528
rect 4632 3942 4660 4519
rect 4724 4010 4752 4950
rect 4816 4758 4844 4966
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4620 3936 4672 3942
rect 4342 3904 4398 3913
rect 4620 3878 4672 3884
rect 4342 3839 4398 3848
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3698 3224 3754 3233
rect 3804 3194 3832 3402
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4264 3194 4292 3538
rect 4434 3496 4490 3505
rect 4434 3431 4490 3440
rect 3698 3159 3754 3168
rect 3792 3188 3844 3194
rect 3712 2990 3740 3159
rect 3792 3130 3844 3136
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3344 2746 3648 2774
rect 2778 2680 2834 2689
rect 2778 2615 2834 2624
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2700 1970 2728 2450
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2976 2038 3004 2246
rect 2964 2032 3016 2038
rect 2964 1974 3016 1980
rect 2688 1964 2740 1970
rect 2688 1906 2740 1912
rect 2226 1456 2282 1465
rect 2226 1391 2282 1400
rect 3068 800 3096 2314
rect 1766 640 1822 649
rect 1766 575 1822 584
rect 2134 0 2190 800
rect 3054 0 3110 800
rect 3344 241 3372 2746
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3528 2106 3556 2450
rect 4448 2446 4476 3431
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4540 2854 4568 3130
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4632 2582 4660 3334
rect 4724 2990 4752 3334
rect 4816 2990 4844 4218
rect 4908 3738 4936 5714
rect 5000 4593 5028 6870
rect 5092 6866 5120 9318
rect 5448 8900 5500 8906
rect 5368 8860 5448 8888
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8498 5304 8774
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5368 8430 5396 8860
rect 5448 8842 5500 8848
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5092 4758 5120 6802
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 6254 5212 6598
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5276 6100 5304 8230
rect 5184 6072 5304 6100
rect 5184 5642 5212 6072
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 4752 5132 4758
rect 5184 4729 5212 5306
rect 5276 5166 5304 5850
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5368 5030 5396 8366
rect 5460 7041 5488 8502
rect 5446 7032 5502 7041
rect 5446 6967 5502 6976
rect 5460 6934 5488 6967
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5552 6610 5580 9318
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8566 5672 8978
rect 5736 8634 5764 9438
rect 5906 9415 5962 9424
rect 5920 9382 5948 9415
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 6730 5672 8298
rect 5736 8294 5764 8570
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5828 8090 5856 8910
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5736 6866 5764 8026
rect 5920 7954 5948 8434
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5920 7818 5948 7890
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5920 7546 5948 7754
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5552 6582 5672 6610
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5460 5370 5488 6190
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5552 5914 5580 6122
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5644 5778 5672 6582
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5736 4808 5764 6802
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 6322 5856 6598
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6012 5250 6040 9982
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6104 9382 6132 9522
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 9042 6132 9318
rect 6196 9178 6224 10406
rect 6288 10266 6316 10639
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6288 9353 6316 9454
rect 6274 9344 6330 9353
rect 6274 9279 6330 9288
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6380 9042 6408 10542
rect 6472 9926 6500 10968
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9081 6500 9862
rect 6458 9072 6514 9081
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6368 9036 6420 9042
rect 6458 9007 6514 9016
rect 6368 8978 6420 8984
rect 6276 8968 6328 8974
rect 6090 8936 6146 8945
rect 6276 8910 6328 8916
rect 6090 8871 6146 8880
rect 6104 7585 6132 8871
rect 6288 8634 6316 8910
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 8430 6408 8978
rect 6460 8968 6512 8974
rect 6458 8936 6460 8945
rect 6512 8936 6514 8945
rect 6458 8871 6514 8880
rect 6368 8424 6420 8430
rect 6182 8392 6238 8401
rect 6368 8366 6420 8372
rect 6182 8327 6238 8336
rect 6276 8356 6328 8362
rect 6196 7970 6224 8327
rect 6276 8298 6328 8304
rect 6288 8090 6316 8298
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6196 7942 6316 7970
rect 6090 7576 6146 7585
rect 6090 7511 6146 7520
rect 6104 7206 6132 7511
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 5644 4780 5764 4808
rect 5828 5222 6040 5250
rect 5080 4694 5132 4700
rect 5170 4720 5226 4729
rect 4986 4584 5042 4593
rect 4986 4519 5042 4528
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5092 3602 5120 4694
rect 5170 4655 5226 4664
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5184 3466 5212 4655
rect 5264 4616 5316 4622
rect 5540 4616 5592 4622
rect 5264 4558 5316 4564
rect 5538 4584 5540 4593
rect 5592 4584 5594 4593
rect 5276 4146 5304 4558
rect 5538 4519 5594 4528
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5368 4214 5396 4422
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4908 2854 4936 2994
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4816 2650 4844 2790
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3804 1170 3832 2314
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 3804 1142 4016 1170
rect 3988 800 4016 1142
rect 4908 800 4936 2314
rect 5092 2310 5120 2450
rect 5276 2446 5304 4082
rect 5368 3602 5396 4150
rect 5460 4146 5488 4422
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5540 4072 5592 4078
rect 5538 4040 5540 4049
rect 5592 4040 5594 4049
rect 5538 3975 5594 3984
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 3505 5396 3538
rect 5354 3496 5410 3505
rect 5644 3482 5672 4780
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5736 4146 5764 4626
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3641 5764 3878
rect 5722 3632 5778 3641
rect 5722 3567 5778 3576
rect 5354 3431 5410 3440
rect 5460 3454 5764 3482
rect 5460 3398 5488 3454
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5736 3058 5764 3454
rect 5828 3097 5856 5222
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5814 3088 5870 3097
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5724 3052 5776 3058
rect 5814 3023 5870 3032
rect 5724 2994 5776 3000
rect 5368 2854 5396 2994
rect 5828 2990 5856 3023
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5092 1834 5120 2246
rect 5920 1902 5948 5102
rect 6104 4536 6132 7142
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 4690 6224 6054
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6288 4570 6316 7942
rect 6380 7342 6408 8366
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6472 7546 6500 8230
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6564 7154 6592 11070
rect 6748 10996 6776 11766
rect 6840 11694 6868 12038
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6656 10968 6776 10996
rect 6656 9874 6684 10968
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6748 10062 6776 10474
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 7300 10146 7328 12310
rect 7484 11694 7512 13262
rect 7760 12782 7788 14214
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12850 8064 13262
rect 8128 12918 8156 13942
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 11937 7788 12310
rect 7746 11928 7802 11937
rect 7746 11863 7802 11872
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10266 7420 11086
rect 7484 11014 7512 11630
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11393 8156 11494
rect 8114 11384 8170 11393
rect 8114 11319 8170 11328
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10606 7512 10950
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7472 10192 7524 10198
rect 7104 10124 7156 10130
rect 7300 10118 7420 10146
rect 7472 10134 7524 10140
rect 7104 10066 7156 10072
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6656 9846 6776 9874
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 8090 6684 9454
rect 6748 9160 6776 9846
rect 6932 9654 6960 9998
rect 7116 9926 7144 10066
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7300 9382 7328 9522
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7288 9172 7340 9178
rect 6748 9132 6868 9160
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8084 6696 8090
rect 6748 8072 6776 8774
rect 6840 8401 6868 9132
rect 7288 9114 7340 9120
rect 6826 8392 6882 8401
rect 6826 8327 6882 8336
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 6748 8044 6868 8072
rect 6644 8026 6696 8032
rect 6656 7342 6684 8026
rect 6840 7993 6868 8044
rect 6826 7984 6882 7993
rect 6826 7919 6882 7928
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7546 6776 7822
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6840 7478 6868 7919
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 7116 7410 7144 7822
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6380 7126 6592 7154
rect 6380 4690 6408 7126
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6472 6118 6500 6870
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6564 5370 6592 6870
rect 6748 6866 6776 7346
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6032 4508 6132 4536
rect 6196 4542 6316 4570
rect 6032 4468 6060 4508
rect 6012 4440 6060 4468
rect 6012 3194 6040 4440
rect 6090 3904 6146 3913
rect 6090 3839 6146 3848
rect 6104 3670 6132 3839
rect 6092 3664 6144 3670
rect 6196 3641 6224 4542
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6092 3606 6144 3612
rect 6182 3632 6238 3641
rect 6182 3567 6238 3576
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6012 2854 6040 3130
rect 6196 2990 6224 3334
rect 6288 3058 6316 4422
rect 6380 4282 6408 4626
rect 6656 4554 6684 6734
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6840 6186 6868 6666
rect 6828 6180 6880 6186
rect 6748 6140 6828 6168
rect 6748 5760 6776 6140
rect 6828 6122 6880 6128
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 6828 5772 6880 5778
rect 6748 5732 6828 5760
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6564 4026 6592 4490
rect 6380 3998 6592 4026
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6288 2582 6316 2790
rect 6380 2582 6408 3998
rect 6748 3942 6776 5732
rect 6828 5714 6880 5720
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6840 4486 6868 4694
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 7300 4078 7328 9114
rect 7392 8809 7420 10118
rect 7484 9674 7512 10134
rect 7576 9926 7604 10746
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7484 9646 7604 9674
rect 7668 9654 7696 11154
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7852 10810 7880 11018
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7760 10130 7788 10474
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 10130 7880 10406
rect 7944 10266 7972 11086
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7378 8800 7434 8809
rect 7378 8735 7434 8744
rect 7392 7886 7420 8735
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7449 7420 7822
rect 7484 7546 7512 7890
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7378 7440 7434 7449
rect 7576 7426 7604 9646
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7378 7375 7434 7384
rect 7484 7398 7604 7426
rect 7392 4808 7420 7375
rect 7484 5778 7512 7398
rect 7654 7304 7710 7313
rect 7564 7268 7616 7274
rect 7654 7239 7656 7248
rect 7564 7210 7616 7216
rect 7708 7239 7710 7248
rect 7656 7210 7708 7216
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7392 4780 7512 4808
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6472 2650 6500 3878
rect 6564 2990 6592 3878
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6734 3768 6790 3777
rect 6644 3732 6696 3738
rect 6886 3760 7182 3780
rect 7392 3738 7420 4626
rect 7484 4554 7512 4780
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 6734 3703 6790 3712
rect 7380 3732 7432 3738
rect 6644 3674 6696 3680
rect 6656 3534 6684 3674
rect 6748 3602 6776 3703
rect 7380 3674 7432 3680
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6656 2922 6684 3334
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6276 2576 6328 2582
rect 6276 2518 6328 2524
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6656 2446 6684 2858
rect 6748 2825 6776 3334
rect 7208 3074 7236 3334
rect 7208 3046 7328 3074
rect 6734 2816 6790 2825
rect 6734 2751 6790 2760
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 6288 1902 6316 2246
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 6276 1896 6328 1902
rect 6276 1838 6328 1844
rect 5080 1828 5132 1834
rect 5080 1770 5132 1776
rect 6380 1170 6408 2246
rect 5828 1142 6408 1170
rect 5828 800 5856 1142
rect 6748 800 6776 2382
rect 6932 2038 6960 2450
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 7300 1970 7328 3046
rect 7484 2582 7512 3878
rect 7576 3602 7604 7210
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7668 4622 7696 5238
rect 7760 5030 7788 10066
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 9042 7880 9522
rect 8036 9450 8064 9862
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8634 7880 8978
rect 7944 8974 7972 9318
rect 8128 9194 8156 11319
rect 8220 10198 8248 14282
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 11532 14074 11560 14418
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8312 11558 8340 12922
rect 8404 12170 8432 13330
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 12986 8524 13194
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8496 12238 8524 12922
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8588 12442 8616 12854
rect 8576 12436 8628 12442
rect 8628 12396 8800 12424
rect 8576 12378 8628 12384
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 8496 11694 8524 12174
rect 8680 12102 8708 12174
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9586 8248 9862
rect 8312 9654 8340 11154
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10266 8432 10950
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8390 10160 8446 10169
rect 8390 10095 8446 10104
rect 8404 9994 8432 10095
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8496 9738 8524 11154
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8404 9722 8524 9738
rect 8588 9722 8616 10406
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8392 9716 8524 9722
rect 8444 9710 8524 9716
rect 8576 9716 8628 9722
rect 8392 9658 8444 9664
rect 8576 9658 8628 9664
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8036 9166 8156 9194
rect 8220 9178 8248 9522
rect 8680 9518 8708 9998
rect 8576 9512 8628 9518
rect 8298 9480 8354 9489
rect 8576 9454 8628 9460
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8298 9415 8354 9424
rect 8312 9382 8340 9415
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 9172 8260 9178
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8036 8786 8064 9166
rect 8208 9114 8260 9120
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8206 9072 8262 9081
rect 7944 8758 8064 8786
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7944 8537 7972 8758
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7930 8528 7986 8537
rect 7930 8463 7986 8472
rect 7840 7404 7892 7410
rect 7944 7392 7972 8463
rect 8036 8090 8064 8570
rect 8128 8129 8156 9046
rect 8312 9042 8340 9318
rect 8588 9178 8616 9454
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8206 9007 8262 9016
rect 8300 9036 8352 9042
rect 8220 8820 8248 9007
rect 8300 8978 8352 8984
rect 8496 8838 8524 9046
rect 8300 8832 8352 8838
rect 8220 8792 8300 8820
rect 8484 8832 8536 8838
rect 8300 8774 8352 8780
rect 8482 8800 8484 8809
rect 8536 8800 8538 8809
rect 8114 8120 8170 8129
rect 8024 8084 8076 8090
rect 8114 8055 8170 8064
rect 8024 8026 8076 8032
rect 7892 7364 7972 7392
rect 7840 7346 7892 7352
rect 7944 6848 7972 7364
rect 8312 7313 8340 8774
rect 8482 8735 8538 8744
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8496 8090 8524 8298
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8404 7886 8432 7958
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8298 7304 8354 7313
rect 8220 7262 8298 7290
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6934 8156 7142
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8024 6860 8076 6866
rect 7944 6820 8024 6848
rect 8024 6802 8076 6808
rect 8128 6390 8156 6870
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5030 7880 5714
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7760 3670 7788 4966
rect 7944 4622 7972 6054
rect 8116 5840 8168 5846
rect 8114 5808 8116 5817
rect 8168 5808 8170 5817
rect 8114 5743 8170 5752
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8036 4604 8064 5170
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4826 8156 4966
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8116 4616 8168 4622
rect 8036 4576 8116 4604
rect 7944 4282 7972 4558
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8036 4010 8064 4576
rect 8116 4558 8168 4564
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7760 3466 7788 3606
rect 8036 3534 8064 3946
rect 8220 3738 8248 7262
rect 8298 7239 8354 7248
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 6254 8340 7142
rect 8404 7002 8432 7822
rect 8482 7576 8538 7585
rect 8482 7511 8538 7520
rect 8496 7478 8524 7511
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8496 6934 8524 7414
rect 8680 7342 8708 8230
rect 8772 7546 8800 12396
rect 8864 11898 8892 13262
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 8956 12434 8984 13126
rect 8956 12406 9076 12434
rect 8942 11928 8998 11937
rect 8852 11892 8904 11898
rect 8942 11863 8944 11872
rect 8852 11834 8904 11840
rect 8996 11863 8998 11872
rect 8944 11834 8996 11840
rect 8864 11286 8892 11834
rect 9048 11778 9076 12406
rect 9232 12102 9260 13126
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9508 12374 9536 12650
rect 9600 12442 9628 13262
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 8956 11750 9076 11778
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8484 6928 8536 6934
rect 8390 6896 8446 6905
rect 8484 6870 8536 6876
rect 8390 6831 8446 6840
rect 8404 6458 8432 6831
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8496 6322 8524 6598
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8312 5166 8340 6190
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5370 8432 6054
rect 8496 5914 8524 6258
rect 8588 6118 8616 7278
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8588 5710 8616 6054
rect 8576 5704 8628 5710
rect 8482 5672 8538 5681
rect 8576 5646 8628 5652
rect 8482 5607 8538 5616
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8390 5264 8446 5273
rect 8496 5250 8524 5607
rect 8496 5234 8616 5250
rect 8496 5228 8628 5234
rect 8496 5222 8576 5228
rect 8390 5199 8446 5208
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4486 8340 4966
rect 8404 4486 8432 5199
rect 8576 5170 8628 5176
rect 8484 4616 8536 4622
rect 8482 4584 8484 4593
rect 8536 4584 8538 4593
rect 8482 4519 8538 4528
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8680 4282 8708 7278
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8772 5234 8800 6666
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 8036 3194 8064 3470
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7288 1964 7340 1970
rect 7288 1906 7340 1912
rect 7576 800 7604 2314
rect 7668 1902 7696 2858
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8312 2106 8340 2790
rect 8588 2582 8616 2790
rect 8680 2582 8708 3334
rect 8864 2990 8892 9862
rect 8956 3670 8984 11750
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 8294 9076 11494
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9140 9178 9168 10950
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 7750 9076 8230
rect 9126 8120 9182 8129
rect 9126 8055 9182 8064
rect 9140 7750 9168 8055
rect 9232 7868 9260 12038
rect 9324 11694 9352 12174
rect 9416 11694 9444 12310
rect 9508 11762 9536 12310
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9586 12200 9642 12209
rect 9586 12135 9588 12144
rect 9640 12135 9642 12144
rect 9588 12106 9640 12112
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9600 11558 9628 12106
rect 9784 11898 9812 12242
rect 10428 12238 10456 12718
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10230 11928 10286 11937
rect 9772 11892 9824 11898
rect 10336 11898 10364 12106
rect 10230 11863 10286 11872
rect 10324 11892 10376 11898
rect 9772 11834 9824 11840
rect 10244 11694 10272 11863
rect 10324 11834 10376 11840
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9416 10713 9444 11494
rect 10428 11354 10456 12174
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 9402 10704 9458 10713
rect 9324 10662 9402 10690
rect 9324 8022 9352 10662
rect 9402 10639 9458 10648
rect 9600 10266 9628 11290
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10428 10606 10456 11290
rect 10520 10742 10548 13874
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11532 13190 11560 13398
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 8022 9444 8230
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9232 7840 9352 7868
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9048 6338 9076 7686
rect 9324 7342 9352 7840
rect 9312 7336 9364 7342
rect 9508 7290 9536 10066
rect 9692 10062 9720 10474
rect 10324 10192 10376 10198
rect 10322 10160 10324 10169
rect 10376 10160 10378 10169
rect 10520 10130 10548 10678
rect 10322 10095 10378 10104
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 9784 9518 9812 9930
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9954 9480 10010 9489
rect 9954 9415 10010 9424
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9312 7278 9364 7284
rect 9048 6310 9260 6338
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9048 5216 9076 5714
rect 9140 5370 9168 6122
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9232 5302 9260 6310
rect 9220 5296 9272 5302
rect 9324 5273 9352 7278
rect 9416 7262 9536 7290
rect 9416 5778 9444 7262
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 6186 9536 7142
rect 9600 6798 9628 8774
rect 9692 8566 9720 9318
rect 9968 9178 9996 9415
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9692 6866 9720 8502
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9784 7818 9812 8366
rect 10140 7880 10192 7886
rect 10244 7868 10272 8910
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10192 7840 10272 7868
rect 10140 7822 10192 7828
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7410 9812 7754
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9220 5238 9272 5244
rect 9310 5264 9366 5273
rect 9128 5228 9180 5234
rect 9048 5188 9128 5216
rect 9128 5170 9180 5176
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 4486 9076 4966
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9140 4282 9168 5170
rect 9232 5166 9260 5238
rect 9310 5199 9366 5208
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9232 4690 9260 5102
rect 9416 4826 9444 5714
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9034 3768 9090 3777
rect 9232 3738 9260 3878
rect 9034 3703 9036 3712
rect 9088 3703 9090 3712
rect 9220 3732 9272 3738
rect 9036 3674 9088 3680
rect 9220 3674 9272 3680
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3194 8984 3334
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8956 2774 8984 3130
rect 8864 2746 8984 2774
rect 8864 2650 8892 2746
rect 9048 2650 9076 3674
rect 9508 3534 9536 6122
rect 9600 4146 9628 6598
rect 9692 6100 9720 6802
rect 10244 6730 10272 7210
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 9864 6112 9916 6118
rect 9692 6072 9864 6100
rect 9864 6054 9916 6060
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9692 5166 9720 5782
rect 9784 5370 9812 5850
rect 9876 5710 9904 6054
rect 10152 5846 10180 6326
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9864 5704 9916 5710
rect 10336 5658 10364 8298
rect 10428 7002 10456 8774
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 9864 5646 9916 5652
rect 10244 5630 10364 5658
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3641 9628 3878
rect 9692 3738 9720 4490
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9586 3632 9642 3641
rect 9586 3567 9642 3576
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9324 2582 9352 3402
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 8496 800 8524 2382
rect 9416 800 9444 3402
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 1766 9720 3334
rect 9784 3194 9812 4626
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3670 10088 3878
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9876 2650 9904 2858
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10152 2650 10180 2790
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10244 2446 10272 5630
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10336 4146 10364 5510
rect 10520 5030 10548 9930
rect 10612 7936 10640 12582
rect 10704 11626 10732 12718
rect 10796 12374 10824 12786
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 11762 10824 12310
rect 10874 12200 10930 12209
rect 10874 12135 10930 12144
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10690 11520 10746 11529
rect 10690 11455 10746 11464
rect 10704 11286 10732 11455
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 9518 10732 11018
rect 10796 10810 10824 11698
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10784 9988 10836 9994
rect 10888 9976 10916 12135
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10980 11354 11008 11494
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11072 11218 11100 11494
rect 11164 11354 11192 12854
rect 11532 12714 11560 13126
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12374 11468 12582
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11716 12288 11744 13806
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12442 11928 13330
rect 12084 12646 12112 14010
rect 12360 12986 12388 14418
rect 12728 13870 12756 14826
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 14384 14550 14412 16400
rect 16394 15600 16450 15609
rect 16394 15535 16450 15544
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14752 14074 14780 14418
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14936 14006 14964 14214
rect 15028 14074 15056 14418
rect 15198 14376 15254 14385
rect 15198 14311 15200 14320
rect 15252 14311 15254 14320
rect 15200 14282 15252 14288
rect 15304 14074 15332 14894
rect 16408 14890 16436 15535
rect 15476 14884 15528 14890
rect 15476 14826 15528 14832
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 15396 13938 15424 14214
rect 15488 14074 15516 14826
rect 16408 14550 16436 14826
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15764 13926 16068 13954
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 13372 12782 13400 13262
rect 13832 12850 13860 13466
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 13372 12442 13400 12718
rect 14016 12714 14044 12854
rect 14108 12850 14136 13194
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 11888 12300 11940 12306
rect 11716 12260 11888 12288
rect 11334 11928 11390 11937
rect 11334 11863 11390 11872
rect 11244 11552 11296 11558
rect 11242 11520 11244 11529
rect 11296 11520 11298 11529
rect 11242 11455 11298 11464
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11242 11248 11298 11257
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11152 11212 11204 11218
rect 11242 11183 11298 11192
rect 11152 11154 11204 11160
rect 10968 10600 11020 10606
rect 11060 10600 11112 10606
rect 10968 10542 11020 10548
rect 11058 10568 11060 10577
rect 11112 10568 11114 10577
rect 10836 9948 10916 9976
rect 10784 9930 10836 9936
rect 10980 9586 11008 10542
rect 11058 10503 11114 10512
rect 11164 9994 11192 11154
rect 11256 11150 11284 11183
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11256 10062 11284 10678
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11060 9648 11112 9654
rect 11058 9616 11060 9625
rect 11112 9616 11114 9625
rect 10968 9580 11020 9586
rect 11058 9551 11114 9560
rect 10968 9522 11020 9528
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10704 8906 10732 9454
rect 11072 8974 11100 9551
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 9178 11284 9318
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11060 8968 11112 8974
rect 11164 8945 11192 9046
rect 11060 8910 11112 8916
rect 11150 8936 11206 8945
rect 10692 8900 10744 8906
rect 11150 8871 11206 8880
rect 10692 8842 10744 8848
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10612 7908 10824 7936
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10612 5778 10640 6326
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10428 4078 10456 4966
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10520 3505 10548 3538
rect 10612 3534 10640 5714
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10704 5030 10732 5510
rect 10796 5137 10824 7908
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10888 5166 10916 7822
rect 10980 7274 11008 8434
rect 11256 8294 11284 9114
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11072 7449 11100 7890
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11058 7440 11114 7449
rect 11058 7375 11114 7384
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10968 6928 11020 6934
rect 11072 6916 11100 7375
rect 11020 6888 11100 6916
rect 10968 6870 11020 6876
rect 11164 6662 11192 7754
rect 11244 7744 11296 7750
rect 11348 7732 11376 11863
rect 11716 11558 11744 12260
rect 11888 12242 11940 12248
rect 12084 12102 12112 12310
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12544 12209 12572 12242
rect 12530 12200 12586 12209
rect 12530 12135 12586 12144
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12162 11928 12218 11937
rect 12544 11898 12572 12135
rect 12162 11863 12218 11872
rect 12532 11892 12584 11898
rect 11888 11824 11940 11830
rect 11886 11792 11888 11801
rect 11940 11792 11942 11801
rect 11886 11727 11942 11736
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11440 11132 11468 11290
rect 11520 11144 11572 11150
rect 11440 11104 11520 11132
rect 11520 11086 11572 11092
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11532 10606 11560 10746
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11440 9178 11468 9998
rect 11532 9178 11560 10542
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11624 9926 11652 10474
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11624 9382 11652 9862
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11624 9042 11652 9318
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11532 8362 11560 8910
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11426 7848 11482 7857
rect 11426 7783 11482 7792
rect 11296 7704 11376 7732
rect 11244 7686 11296 7692
rect 11256 7274 11284 7686
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11152 6656 11204 6662
rect 11072 6616 11152 6644
rect 11072 6458 11100 6616
rect 11152 6598 11204 6604
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11060 6248 11112 6254
rect 11058 6216 11060 6225
rect 11112 6216 11114 6225
rect 11058 6151 11114 6160
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5234 11008 6054
rect 11164 5953 11192 6394
rect 11150 5944 11206 5953
rect 11150 5879 11206 5888
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10876 5160 10928 5166
rect 10782 5128 10838 5137
rect 10876 5102 10928 5108
rect 10782 5063 10838 5072
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10704 4185 10732 4694
rect 10690 4176 10746 4185
rect 10690 4111 10746 4120
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10600 3528 10652 3534
rect 10506 3496 10562 3505
rect 10600 3470 10652 3476
rect 10506 3431 10562 3440
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 10336 800 10364 2858
rect 10428 2854 10456 3130
rect 10704 3058 10732 3606
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10796 2774 10824 5063
rect 10966 4720 11022 4729
rect 10966 4655 11022 4664
rect 10980 4486 11008 4655
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10888 3777 10916 4150
rect 10966 4040 11022 4049
rect 10966 3975 11022 3984
rect 10874 3768 10930 3777
rect 10874 3703 10876 3712
rect 10928 3703 10930 3712
rect 10876 3674 10928 3680
rect 10888 3602 10916 3674
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10980 3466 11008 3975
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 10888 3233 10916 3402
rect 10874 3224 10930 3233
rect 11072 3194 11100 5714
rect 11164 4622 11192 5782
rect 11348 5778 11376 7142
rect 11440 6934 11468 7783
rect 11532 7206 11560 7958
rect 11624 7410 11652 8978
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11348 4758 11376 5510
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11440 4690 11468 6870
rect 11532 6322 11560 7142
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11518 5944 11574 5953
rect 11518 5879 11574 5888
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4146 11192 4558
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11244 4276 11296 4282
rect 11348 4264 11376 4422
rect 11296 4236 11376 4264
rect 11244 4218 11296 4224
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11440 4026 11468 4626
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11348 3998 11468 4026
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10874 3159 10930 3168
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10520 2746 10824 2774
rect 10414 2680 10470 2689
rect 10414 2615 10416 2624
rect 10468 2615 10470 2624
rect 10416 2586 10468 2592
rect 10520 1834 10548 2746
rect 11072 2514 11100 2994
rect 11164 2650 11192 3878
rect 11256 3369 11284 3946
rect 11348 3602 11376 3998
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11242 3360 11298 3369
rect 11242 3295 11298 3304
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11348 2582 11376 3538
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 10508 1828 10560 1834
rect 10508 1770 10560 1776
rect 11256 800 11284 2314
rect 11440 2310 11468 3878
rect 11532 2514 11560 5879
rect 11624 5658 11652 7346
rect 11716 6934 11744 11494
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10418 11836 11086
rect 11900 11014 11928 11222
rect 12084 11218 12112 11698
rect 12176 11558 12204 11863
rect 12532 11834 12584 11840
rect 12256 11688 12308 11694
rect 12254 11656 12256 11665
rect 12308 11656 12310 11665
rect 12254 11591 12310 11600
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12452 11354 12480 11494
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12532 11280 12584 11286
rect 12452 11228 12532 11234
rect 12452 11222 12584 11228
rect 12622 11248 12678 11257
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12452 11206 12572 11222
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11992 10606 12020 11086
rect 12084 10742 12112 11154
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11808 10390 12020 10418
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11808 8634 11836 9454
rect 11900 9382 11928 10134
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11808 6254 11836 8230
rect 11900 6254 11928 9318
rect 11992 9081 12020 10390
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12084 10033 12112 10066
rect 12256 10056 12308 10062
rect 12070 10024 12126 10033
rect 12256 9998 12308 10004
rect 12070 9959 12126 9968
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12084 9489 12112 9590
rect 12070 9480 12126 9489
rect 12070 9415 12126 9424
rect 12268 9178 12296 9998
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12072 9172 12124 9178
rect 12256 9172 12308 9178
rect 12124 9132 12204 9160
rect 12072 9114 12124 9120
rect 11978 9072 12034 9081
rect 11978 9007 12034 9016
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 6458 12020 6734
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11992 5778 12020 6258
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11624 5630 11744 5658
rect 11716 5574 11744 5630
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11900 4706 11928 5578
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11624 4690 11928 4706
rect 11612 4684 11928 4690
rect 11664 4678 11928 4684
rect 11612 4626 11664 4632
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11624 4457 11652 4490
rect 11610 4448 11666 4457
rect 11610 4383 11666 4392
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11624 3534 11652 4082
rect 11716 3738 11744 4558
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11808 3058 11836 4558
rect 11900 4010 11928 4678
rect 11992 4078 12020 4762
rect 12084 4758 12112 8298
rect 12176 6361 12204 9132
rect 12256 9114 12308 9120
rect 12360 9110 12388 9318
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12360 8838 12388 9046
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 7546 12296 8230
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12162 6352 12218 6361
rect 12162 6287 12218 6296
rect 12164 6248 12216 6254
rect 12268 6236 12296 6938
rect 12216 6208 12296 6236
rect 12164 6190 12216 6196
rect 12176 5642 12204 6190
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12360 5817 12388 6054
rect 12346 5808 12402 5817
rect 12346 5743 12402 5752
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12254 4856 12310 4865
rect 12254 4791 12256 4800
rect 12308 4791 12310 4800
rect 12256 4762 12308 4768
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12268 4622 12296 4762
rect 12360 4622 12388 4966
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11992 3942 12020 4014
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 12072 3664 12124 3670
rect 11992 3624 12072 3652
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11900 3126 11928 3538
rect 11992 3194 12020 3624
rect 12072 3606 12124 3612
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11888 3120 11940 3126
rect 12084 3097 12112 3130
rect 11888 3062 11940 3068
rect 12070 3088 12126 3097
rect 11796 3052 11848 3058
rect 12176 3058 12204 3946
rect 12070 3023 12126 3032
rect 12164 3052 12216 3058
rect 11796 2994 11848 3000
rect 12164 2994 12216 3000
rect 12268 2990 12296 4422
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12360 3602 12388 3878
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12452 3482 12480 11206
rect 12622 11183 12624 11192
rect 12676 11183 12678 11192
rect 12624 11154 12676 11160
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 9994 12664 10474
rect 12728 10266 12756 11494
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 13188 11354 13216 11494
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12530 9480 12586 9489
rect 12530 9415 12586 9424
rect 12624 9444 12676 9450
rect 12544 9178 12572 9415
rect 12624 9386 12676 9392
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12636 8922 12664 9386
rect 12728 9178 12756 10066
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9364 13032 9862
rect 13188 9738 13216 11086
rect 13280 10130 13308 12310
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13820 11824 13872 11830
rect 13450 11792 13506 11801
rect 13820 11766 13872 11772
rect 13450 11727 13506 11736
rect 13636 11756 13688 11762
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13372 11286 13400 11562
rect 13464 11558 13492 11727
rect 13636 11698 13688 11704
rect 13648 11558 13676 11698
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13372 10010 13400 11222
rect 13464 11218 13492 11494
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13648 11150 13676 11494
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10538 13584 10950
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13452 10464 13504 10470
rect 13504 10412 13584 10418
rect 13452 10406 13584 10412
rect 13464 10390 13584 10406
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13280 9982 13400 10010
rect 13280 9926 13308 9982
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13188 9710 13308 9738
rect 13004 9336 13216 9364
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13188 9178 13216 9336
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12544 8906 12664 8922
rect 12532 8900 12664 8906
rect 12584 8894 12664 8900
rect 12532 8842 12584 8848
rect 12544 8090 12572 8842
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12636 7818 12664 8434
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12728 7546 12756 8298
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 13188 8090 13216 8230
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12532 7472 12584 7478
rect 12584 7432 12664 7460
rect 12532 7414 12584 7420
rect 12636 7313 12664 7432
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12622 7304 12678 7313
rect 12622 7239 12624 7248
rect 12676 7239 12678 7248
rect 12624 7210 12676 7216
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12636 5846 12664 6870
rect 12728 6798 12756 7346
rect 13280 7206 13308 9710
rect 13372 9178 13400 9862
rect 13464 9722 13492 10134
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13556 9489 13584 10390
rect 13740 10062 13768 11018
rect 13832 11014 13860 11766
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13818 10160 13874 10169
rect 13818 10095 13874 10104
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9722 13768 9998
rect 13832 9722 13860 10095
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13542 9480 13598 9489
rect 13542 9415 13598 9424
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13452 9376 13504 9382
rect 13450 9344 13452 9353
rect 13504 9344 13506 9353
rect 13450 9279 13506 9288
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13464 8974 13492 9279
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13634 9072 13690 9081
rect 13634 9007 13690 9016
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 13004 6458 13032 6802
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13188 6186 13216 7142
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12544 5030 12572 5782
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4826 12664 4966
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 13188 3738 13216 6122
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 12452 3454 12664 3482
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 11900 2650 11928 2858
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11716 2514 11744 2586
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 12176 800 12204 2858
rect 12360 2854 12388 3334
rect 12636 2990 12664 3454
rect 13188 3126 13216 3674
rect 13280 3505 13308 3878
rect 13266 3496 13322 3505
rect 13266 3431 13322 3440
rect 13280 3126 13308 3431
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12820 2922 12848 3062
rect 13188 2990 13216 3062
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2650 12480 2790
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 13372 2514 13400 8230
rect 13464 7750 13492 8910
rect 13648 8906 13676 9007
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13740 8498 13768 9114
rect 13832 9042 13860 9386
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13818 8936 13874 8945
rect 13924 8922 13952 12038
rect 14016 11937 14044 12650
rect 14096 12640 14148 12646
rect 14280 12640 14332 12646
rect 14148 12600 14228 12628
rect 14096 12582 14148 12588
rect 14200 12238 14228 12600
rect 14280 12582 14332 12588
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14002 11928 14058 11937
rect 14002 11863 14058 11872
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14016 11121 14044 11494
rect 14108 11354 14136 11766
rect 14200 11354 14228 12174
rect 14292 11898 14320 12582
rect 14384 12434 14412 13466
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14384 12406 14504 12434
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14278 11656 14334 11665
rect 14278 11591 14334 11600
rect 14292 11558 14320 11591
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14002 11112 14058 11121
rect 14002 11047 14058 11056
rect 14108 10962 14136 11290
rect 13874 8894 13952 8922
rect 14016 10934 14136 10962
rect 13818 8871 13874 8880
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13556 8294 13584 8366
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13544 8016 13596 8022
rect 13648 8004 13676 8230
rect 13596 7976 13676 8004
rect 13544 7958 13596 7964
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13556 7342 13584 7822
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 7002 13584 7142
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13556 6322 13584 6666
rect 13648 6458 13676 7346
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5914 13584 6258
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13450 5128 13506 5137
rect 13450 5063 13452 5072
rect 13504 5063 13506 5072
rect 13452 5034 13504 5040
rect 13648 2990 13676 5510
rect 13740 4010 13768 7686
rect 13832 7342 13860 8871
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13924 7546 13952 7822
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13818 6896 13874 6905
rect 13874 6840 13952 6848
rect 13818 6831 13820 6840
rect 13872 6820 13952 6840
rect 13820 6802 13872 6808
rect 13818 6352 13874 6361
rect 13818 6287 13874 6296
rect 13832 5914 13860 6287
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13818 5808 13874 5817
rect 13818 5743 13874 5752
rect 13832 5574 13860 5743
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13832 4622 13860 5170
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13924 4282 13952 6820
rect 14016 5778 14044 10934
rect 14292 9674 14320 11494
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 10266 14412 11086
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14108 9646 14320 9674
rect 14108 8945 14136 9646
rect 14094 8936 14150 8945
rect 14476 8922 14504 12406
rect 14568 12374 14596 13194
rect 14752 12986 14780 13330
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14844 12986 14872 13194
rect 15028 13190 15056 13738
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13530 15332 13670
rect 15764 13530 15792 13926
rect 16040 13802 16068 13926
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 15856 13530 15884 13738
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14922 12880 14978 12889
rect 14922 12815 14978 12824
rect 14936 12646 14964 12815
rect 15120 12714 15148 13466
rect 15200 13456 15252 13462
rect 15304 13433 15332 13466
rect 15200 13398 15252 13404
rect 15290 13424 15346 13433
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14568 12170 14596 12310
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14830 12200 14886 12209
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14568 11694 14596 11766
rect 14752 11694 14780 12174
rect 14830 12135 14886 12144
rect 14844 11898 14872 12135
rect 14936 12102 14964 12582
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 15120 11354 15148 12038
rect 15212 11540 15240 13398
rect 15290 13359 15346 13368
rect 15566 13424 15622 13433
rect 15566 13359 15622 13368
rect 15382 13288 15438 13297
rect 15292 13252 15344 13258
rect 15382 13223 15384 13232
rect 15292 13194 15344 13200
rect 15436 13223 15438 13232
rect 15384 13194 15436 13200
rect 15304 12866 15332 13194
rect 15304 12838 15424 12866
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15304 11762 15332 12310
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15212 11512 15332 11540
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14740 11008 14792 11014
rect 14792 10968 14872 10996
rect 14740 10950 14792 10956
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9926 14780 10406
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14094 8871 14150 8880
rect 14292 8894 14504 8922
rect 14556 8900 14608 8906
rect 14108 8838 14136 8871
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14108 7206 14136 8774
rect 14292 8412 14320 8894
rect 14556 8842 14608 8848
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8566 14412 8774
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14292 8384 14412 8412
rect 14384 7313 14412 8384
rect 14476 8022 14504 8434
rect 14568 8294 14596 8842
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14476 7818 14504 7958
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14370 7304 14426 7313
rect 14370 7239 14426 7248
rect 14096 7200 14148 7206
rect 14148 7160 14228 7188
rect 14096 7142 14148 7148
rect 14200 6866 14228 7160
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14108 5574 14136 5714
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 4729 14136 5510
rect 14094 4720 14150 4729
rect 14094 4655 14150 4664
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13832 3670 13860 4082
rect 14016 4078 14044 4422
rect 14004 4072 14056 4078
rect 13910 4040 13966 4049
rect 14004 4014 14056 4020
rect 13910 3975 13966 3984
rect 13924 3738 13952 3975
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13728 3392 13780 3398
rect 13780 3340 13860 3346
rect 13728 3334 13860 3340
rect 13740 3318 13860 3334
rect 13832 3194 13860 3318
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 14200 3097 14228 6802
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6225 14412 6598
rect 14370 6216 14426 6225
rect 14476 6186 14504 7414
rect 14370 6151 14426 6160
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14292 4622 14320 5850
rect 14476 5710 14504 6122
rect 14568 6118 14596 8230
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14384 5166 14412 5510
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14476 5098 14504 5510
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14384 3534 14412 4966
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14476 4282 14504 4626
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14186 3088 14242 3097
rect 14186 3023 14242 3032
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 14660 2514 14688 9862
rect 14752 9518 14780 9862
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14844 9042 14872 10968
rect 15028 10742 15056 11154
rect 15120 11150 15148 11290
rect 15108 11144 15160 11150
rect 15160 11104 15240 11132
rect 15108 11086 15160 11092
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15028 10062 15056 10678
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14844 8401 14872 8978
rect 15028 8974 15056 9862
rect 15212 9450 15240 11104
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 14924 8968 14976 8974
rect 14922 8936 14924 8945
rect 15016 8968 15068 8974
rect 14976 8936 14978 8945
rect 15016 8910 15068 8916
rect 14922 8871 14978 8880
rect 14830 8392 14886 8401
rect 14830 8327 14886 8336
rect 14844 6905 14872 8327
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14830 6896 14886 6905
rect 14830 6831 14886 6840
rect 14844 6662 14872 6831
rect 15028 6798 15056 7686
rect 15212 7546 15240 7890
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 15120 6440 15148 6666
rect 14936 6412 15148 6440
rect 14936 6254 14964 6412
rect 14924 6248 14976 6254
rect 15200 6248 15252 6254
rect 14924 6190 14976 6196
rect 15028 6208 15200 6236
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14752 5030 14780 6054
rect 14844 5914 14872 6122
rect 14936 6118 14964 6190
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14832 5772 14884 5778
rect 15028 5760 15056 6208
rect 15200 6190 15252 6196
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 14884 5732 15056 5760
rect 14832 5714 14884 5720
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14844 4826 14872 5578
rect 15120 5098 15148 5646
rect 15212 5137 15240 5850
rect 15198 5128 15254 5137
rect 15108 5092 15160 5098
rect 15198 5063 15254 5072
rect 15108 5034 15160 5040
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14844 3194 14872 4762
rect 15120 4622 15148 5034
rect 15198 4992 15254 5001
rect 15198 4927 15254 4936
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15120 4146 15148 4558
rect 15212 4146 15240 4927
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15120 3738 15148 4082
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12452 2310 12480 2382
rect 15304 2378 15332 11512
rect 15396 2514 15424 12838
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15488 11898 15516 12650
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15580 11778 15608 13359
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15672 12986 15700 13262
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15672 12374 15700 12718
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15488 11750 15608 11778
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 15488 9042 15516 11750
rect 16040 11218 16068 11766
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16040 10062 16068 10406
rect 15660 10056 15712 10062
rect 15566 10024 15622 10033
rect 15660 9998 15712 10004
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15566 9959 15622 9968
rect 15580 9466 15608 9959
rect 15672 9722 15700 9998
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15580 9438 15700 9466
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15488 8430 15516 8978
rect 15580 8498 15608 9318
rect 15672 9178 15700 9438
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15672 8514 15700 9114
rect 16040 9042 16068 9386
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 15672 8498 15792 8514
rect 15568 8492 15620 8498
rect 15672 8492 15804 8498
rect 15672 8486 15752 8492
rect 15568 8434 15620 8440
rect 15752 8434 15804 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15580 7970 15608 8434
rect 15488 7954 15608 7970
rect 15476 7948 15608 7954
rect 15528 7942 15608 7948
rect 15660 7948 15712 7954
rect 15476 7890 15528 7896
rect 15660 7890 15712 7896
rect 15488 7410 15516 7890
rect 15672 7834 15700 7890
rect 15580 7806 15700 7834
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15580 6730 15608 7806
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 16132 7528 16160 14350
rect 16224 13394 16252 14486
rect 16500 14006 16528 16759
rect 16578 16400 16634 17200
rect 17774 16416 17830 16425
rect 16592 14618 16620 16400
rect 18786 16400 18842 17200
rect 17774 16351 17830 16360
rect 17682 15192 17738 15201
rect 17682 15127 17738 15136
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 17236 14482 17264 14758
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16224 12889 16252 12922
rect 16210 12880 16266 12889
rect 16210 12815 16266 12824
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 10674 16252 12038
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16224 9450 16252 10610
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 15672 7500 16160 7528
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5817 15516 6054
rect 15474 5808 15530 5817
rect 15474 5743 15530 5752
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15580 5234 15608 5714
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15488 4282 15516 4422
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15566 3360 15622 3369
rect 15566 3295 15622 3304
rect 15580 3194 15608 3295
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15580 2582 15608 3130
rect 15672 2650 15700 7500
rect 15934 7440 15990 7449
rect 15934 7375 15990 7384
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 7002 15792 7142
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15948 6730 15976 7375
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 16132 4826 16160 6598
rect 16224 5302 16252 8366
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16316 2990 16344 13874
rect 16408 13530 16436 13942
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16394 13424 16450 13433
rect 16394 13359 16450 13368
rect 16408 13326 16436 13359
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16592 12782 16620 13466
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16500 11694 16528 12582
rect 16578 12472 16634 12481
rect 16578 12407 16634 12416
rect 16592 12374 16620 12407
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16592 12170 16620 12310
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16684 11898 16712 14282
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16776 12850 16804 13466
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16868 12238 16896 12310
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16488 11688 16540 11694
rect 16580 11688 16632 11694
rect 16488 11630 16540 11636
rect 16578 11656 16580 11665
rect 16632 11656 16634 11665
rect 16578 11591 16634 11600
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 11218 16528 11494
rect 16776 11354 16804 11698
rect 16960 11642 16988 13806
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 17052 11898 17080 13398
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12481 17172 13262
rect 17130 12472 17186 12481
rect 17130 12407 17186 12416
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17038 11792 17094 11801
rect 17038 11727 17094 11736
rect 16868 11614 16988 11642
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16868 11234 16896 11614
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16776 11206 16896 11234
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16486 10840 16542 10849
rect 16486 10775 16542 10784
rect 16500 10674 16528 10775
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16394 9752 16450 9761
rect 16394 9687 16396 9696
rect 16448 9687 16450 9696
rect 16396 9658 16448 9664
rect 16500 9518 16528 10202
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16396 9376 16448 9382
rect 16394 9344 16396 9353
rect 16448 9344 16450 9353
rect 16394 9279 16450 9288
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16408 4706 16436 8502
rect 16500 8362 16528 9454
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16500 7274 16528 8026
rect 16592 7410 16620 10950
rect 16776 10713 16804 11206
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16868 10810 16896 11018
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16762 10704 16818 10713
rect 16762 10639 16818 10648
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16684 9722 16712 9930
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 7478 16712 8230
rect 16776 8090 16804 10639
rect 16960 10198 16988 11494
rect 17052 11286 17080 11727
rect 17130 11384 17186 11393
rect 17130 11319 17186 11328
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 17144 11132 17172 11319
rect 17052 11104 17172 11132
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16948 8832 17000 8838
rect 16868 8792 16948 8820
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16500 5234 16528 6666
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16408 4678 16528 4706
rect 16394 4176 16450 4185
rect 16394 4111 16450 4120
rect 16408 3670 16436 4111
rect 16396 3664 16448 3670
rect 16500 3641 16528 4678
rect 16592 4078 16620 5306
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16396 3606 16448 3612
rect 16486 3632 16542 3641
rect 16486 3567 16542 3576
rect 16684 3534 16712 3878
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16776 3466 16804 5714
rect 16868 4010 16896 8792
rect 16948 8774 17000 8780
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 6458 16988 8366
rect 17052 7857 17080 11104
rect 17130 9752 17186 9761
rect 17130 9687 17132 9696
rect 17184 9687 17186 9696
rect 17132 9658 17184 9664
rect 17144 8430 17172 9658
rect 17236 9194 17264 14282
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17328 12374 17356 13874
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17328 11898 17356 12310
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17420 11665 17448 14486
rect 17696 14482 17724 15127
rect 17788 14958 17816 16351
rect 17866 16008 17922 16017
rect 17866 15943 17922 15952
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17684 14476 17736 14482
rect 17512 14436 17684 14464
rect 17512 12850 17540 14436
rect 17684 14418 17736 14424
rect 17788 13938 17816 14894
rect 17880 13954 17908 15943
rect 18050 14784 18106 14793
rect 18050 14719 18106 14728
rect 18064 14550 18092 14719
rect 18052 14544 18104 14550
rect 17972 14504 18052 14532
rect 17972 14074 18000 14504
rect 18052 14486 18104 14492
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17776 13932 17828 13938
rect 17880 13926 18000 13954
rect 17776 13874 17828 13880
rect 17972 13870 18000 13926
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17604 13530 17632 13738
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17696 13297 17724 13330
rect 17682 13288 17738 13297
rect 17682 13223 17738 13232
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17604 11898 17632 13126
rect 17696 12617 17724 13223
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17682 12608 17738 12617
rect 17682 12543 17738 12552
rect 17788 12306 17816 12786
rect 17880 12442 17908 13806
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17972 12322 18000 13262
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17880 12294 18000 12322
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17406 11656 17462 11665
rect 17406 11591 17462 11600
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17328 11354 17356 11494
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17420 10266 17448 11494
rect 17512 11150 17540 11834
rect 17788 11762 17816 12242
rect 17592 11756 17644 11762
rect 17776 11756 17828 11762
rect 17592 11698 17644 11704
rect 17696 11716 17776 11744
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17604 10810 17632 11698
rect 17696 11286 17724 11716
rect 17776 11698 17828 11704
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17604 10470 17632 10746
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17604 9722 17632 10066
rect 17788 9994 17816 10474
rect 17880 10266 17908 12294
rect 18064 12209 18092 14282
rect 18144 14272 18196 14278
rect 18432 14249 18460 14418
rect 18800 14414 18828 16400
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18144 14214 18196 14220
rect 18418 14240 18474 14249
rect 18156 12434 18184 14214
rect 18418 14175 18474 14184
rect 18420 13864 18472 13870
rect 18418 13832 18420 13841
rect 18472 13832 18474 13841
rect 18418 13767 18474 13776
rect 18418 13424 18474 13433
rect 18418 13359 18420 13368
rect 18472 13359 18474 13368
rect 18420 13330 18472 13336
rect 18432 12442 18460 13330
rect 18510 13016 18566 13025
rect 18510 12951 18566 12960
rect 18524 12782 18552 12951
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18972 12504 19024 12510
rect 18972 12446 19024 12452
rect 18420 12436 18472 12442
rect 18156 12406 18276 12434
rect 18050 12200 18106 12209
rect 18050 12135 18106 12144
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17880 10062 17908 10202
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17236 9166 17356 9194
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17038 7848 17094 7857
rect 17038 7783 17094 7792
rect 17144 7546 17172 8366
rect 17236 8090 17264 9046
rect 17328 8514 17356 9166
rect 17420 8906 17448 9386
rect 17788 9382 17816 9930
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9489 17908 9862
rect 17866 9480 17922 9489
rect 17866 9415 17922 9424
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17512 9178 17540 9318
rect 17880 9178 17908 9415
rect 17972 9178 18000 11154
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17328 8486 17448 8514
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17236 7342 17264 7890
rect 17328 7546 17356 8298
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17236 7002 17264 7278
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17420 5930 17448 8486
rect 17604 8378 17632 9114
rect 17868 8424 17920 8430
rect 17512 8350 17632 8378
rect 17866 8392 17868 8401
rect 17920 8392 17922 8401
rect 17512 7002 17540 8350
rect 17866 8327 17922 8336
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17592 8288 17644 8294
rect 17972 8265 18000 8298
rect 17592 8230 17644 8236
rect 17958 8256 18014 8265
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17328 5914 17448 5930
rect 17316 5908 17448 5914
rect 17368 5902 17448 5908
rect 17316 5850 17368 5856
rect 17604 4758 17632 8230
rect 17958 8191 18014 8200
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7546 17908 7958
rect 17958 7848 18014 7857
rect 17958 7783 17960 7792
rect 18012 7783 18014 7792
rect 17960 7754 18012 7760
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17868 7336 17920 7342
rect 17866 7304 17868 7313
rect 17920 7304 17922 7313
rect 18064 7290 18092 11834
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 8430 18184 11494
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18156 7478 18184 7686
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 17866 7239 17922 7248
rect 17972 7262 18092 7290
rect 17880 7002 17908 7239
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17972 6730 18000 7262
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 6934 18092 7142
rect 18142 7032 18198 7041
rect 18142 6967 18198 6976
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18156 6866 18184 6967
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18064 5846 18092 6054
rect 18052 5840 18104 5846
rect 18052 5782 18104 5788
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18064 5166 18092 5510
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4758 18092 4966
rect 18142 4856 18198 4865
rect 18142 4791 18198 4800
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 17420 4078 17448 4694
rect 18156 4690 18184 4791
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 18142 4040 18198 4049
rect 16856 4004 16908 4010
rect 18142 3975 18144 3984
rect 16856 3946 16908 3952
rect 18196 3975 18198 3984
rect 18144 3946 18196 3952
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16868 3398 16896 3946
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3670 17816 3878
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16868 3126 16896 3334
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 17038 3088 17094 3097
rect 17328 3058 17356 3334
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17038 3023 17094 3032
rect 17316 3052 17368 3058
rect 17052 2990 17080 3023
rect 17316 2994 17368 3000
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 16304 2984 16356 2990
rect 16118 2952 16174 2961
rect 15844 2916 15896 2922
rect 16304 2926 16356 2932
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 16118 2887 16174 2896
rect 15844 2858 15896 2864
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15660 2508 15712 2514
rect 15764 2496 15792 2790
rect 15856 2514 15884 2858
rect 16132 2854 16160 2887
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16316 2774 16344 2926
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16316 2746 16620 2774
rect 16592 2514 16620 2746
rect 16960 2582 16988 2790
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 17052 2514 17080 2926
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 15712 2468 15792 2496
rect 15844 2508 15896 2514
rect 15660 2450 15712 2456
rect 15844 2450 15896 2456
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 13096 800 13124 2314
rect 13924 800 13952 2314
rect 14844 800 14872 2314
rect 15672 1986 15700 2450
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 15672 1958 15792 1986
rect 15764 800 15792 1958
rect 16592 1057 16620 2314
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16578 1048 16634 1057
rect 16578 983 16634 992
rect 16684 800 16712 2246
rect 17236 1562 17264 2790
rect 17420 2582 17448 2790
rect 17512 2650 17540 2858
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17224 1556 17276 1562
rect 17224 1498 17276 1504
rect 3330 232 3386 241
rect 3330 167 3386 176
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17512 649 17540 2246
rect 17604 1873 17632 2790
rect 17590 1864 17646 1873
rect 17590 1799 17646 1808
rect 17592 1556 17644 1562
rect 17592 1498 17644 1504
rect 17604 800 17632 1498
rect 17696 1465 17724 2994
rect 17788 2689 17816 3062
rect 17774 2680 17830 2689
rect 17774 2615 17830 2624
rect 17776 2304 17828 2310
rect 17880 2281 17908 3470
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18156 3233 18184 3402
rect 18142 3224 18198 3233
rect 18142 3159 18198 3168
rect 18248 2582 18276 12406
rect 18420 12378 18472 12384
rect 18984 12209 19012 12446
rect 18970 12200 19026 12209
rect 18970 12135 19026 12144
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 6984 18368 12038
rect 18972 11280 19024 11286
rect 18970 11248 18972 11257
rect 19024 11248 19026 11257
rect 18970 11183 19026 11192
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18432 10062 18460 11086
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10441 18552 11018
rect 18604 10464 18656 10470
rect 18510 10432 18566 10441
rect 18604 10406 18656 10412
rect 18510 10367 18566 10376
rect 18616 10198 18644 10406
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18524 9382 18552 10066
rect 18616 10033 18644 10134
rect 18602 10024 18658 10033
rect 18602 9959 18658 9968
rect 18602 9616 18658 9625
rect 18602 9551 18658 9560
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 9217 18552 9318
rect 18510 9208 18566 9217
rect 18510 9143 18566 9152
rect 18418 8800 18474 8809
rect 18418 8735 18474 8744
rect 18432 8634 18460 8735
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18432 8430 18460 8570
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18616 8022 18644 9551
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18510 7440 18566 7449
rect 18510 7375 18512 7384
rect 18564 7375 18566 7384
rect 18512 7346 18564 7352
rect 18340 6956 18460 6984
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18340 6458 18368 6802
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18432 6254 18460 6956
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18524 6633 18552 6666
rect 18510 6624 18566 6633
rect 18510 6559 18566 6568
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18510 6216 18566 6225
rect 18510 6151 18512 6160
rect 18564 6151 18566 6160
rect 18512 6122 18564 6128
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18432 5914 18460 6054
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18510 5672 18566 5681
rect 18510 5607 18512 5616
rect 18564 5607 18566 5616
rect 18512 5578 18564 5584
rect 18510 5264 18566 5273
rect 18510 5199 18512 5208
rect 18564 5199 18566 5208
rect 18512 5170 18564 5176
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18524 4457 18552 4490
rect 18510 4448 18566 4457
rect 18510 4383 18566 4392
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18524 3641 18552 3946
rect 18510 3632 18566 3641
rect 18510 3567 18566 3576
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 2990 18368 3334
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18236 2576 18288 2582
rect 18236 2518 18288 2524
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 17776 2246 17828 2252
rect 17866 2272 17922 2281
rect 17682 1456 17738 1465
rect 17682 1391 17738 1400
rect 17498 640 17554 649
rect 17498 575 17554 584
rect 17590 0 17646 800
rect 17788 241 17816 2246
rect 17866 2207 17922 2216
rect 18524 800 18552 2314
rect 19432 1760 19484 1766
rect 19432 1702 19484 1708
rect 19444 800 19472 1702
rect 17774 232 17830 241
rect 17774 167 17830 176
rect 18510 0 18566 800
rect 19430 0 19486 800
<< via2 >>
rect 3054 16360 3110 16416
rect 3514 16768 3570 16824
rect 2962 15952 3018 16008
rect 2502 15544 2558 15600
rect 2226 15136 2282 15192
rect 1858 14728 1914 14784
rect 2226 14492 2228 14512
rect 2228 14492 2280 14512
rect 2280 14492 2282 14512
rect 2226 14456 2282 14492
rect 1490 14320 1546 14376
rect 1490 13912 1546 13968
rect 1674 13912 1730 13968
rect 1858 13504 1914 13560
rect 1490 13096 1546 13152
rect 1858 12708 1914 12744
rect 1858 12688 1860 12708
rect 1860 12688 1912 12708
rect 1912 12688 1914 12708
rect 1490 12280 1546 12336
rect 1398 11328 1454 11384
rect 2226 11872 2282 11928
rect 1674 10648 1730 10704
rect 2042 10920 2098 10976
rect 1858 10412 1860 10432
rect 1860 10412 1912 10432
rect 1912 10412 1914 10432
rect 1858 10376 1914 10412
rect 1766 10104 1822 10160
rect 16486 16768 16542 16824
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 3606 14492 3608 14512
rect 3608 14492 3660 14512
rect 3660 14492 3662 14512
rect 3606 14456 3662 14492
rect 2870 10512 2926 10568
rect 3054 10512 3110 10568
rect 2318 9968 2374 10024
rect 1490 8880 1546 8936
rect 1490 7248 1546 7304
rect 1766 6860 1822 6896
rect 1766 6840 1768 6860
rect 1768 6840 1820 6860
rect 1820 6840 1822 6860
rect 1490 6432 1546 6488
rect 1858 6060 1860 6080
rect 1860 6060 1912 6080
rect 1912 6060 1914 6080
rect 1858 6024 1914 6060
rect 1490 5480 1546 5536
rect 1858 5072 1914 5128
rect 1398 4700 1400 4720
rect 1400 4700 1452 4720
rect 1452 4700 1454 4720
rect 1398 4664 1454 4700
rect 2042 6996 2098 7032
rect 2042 6976 2044 6996
rect 2044 6976 2096 6996
rect 2096 6976 2098 6996
rect 2134 6196 2136 6216
rect 2136 6196 2188 6216
rect 2188 6196 2190 6216
rect 2134 6160 2190 6196
rect 1766 3168 1822 3224
rect 1582 2932 1584 2952
rect 1584 2932 1636 2952
rect 1636 2932 1638 2952
rect 1582 2896 1638 2932
rect 1490 2216 1546 2272
rect 1398 992 1454 1048
rect 3146 9288 3202 9344
rect 3054 8472 3110 8528
rect 2870 7656 2926 7712
rect 3330 9696 3386 9752
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 5630 13932 5686 13968
rect 5630 13912 5632 13932
rect 5632 13912 5684 13932
rect 5684 13912 5686 13932
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3882 12180 3884 12200
rect 3884 12180 3936 12200
rect 3936 12180 3938 12200
rect 3882 12144 3938 12180
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3606 10240 3662 10296
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 4066 10124 4122 10160
rect 4066 10104 4068 10124
rect 4068 10104 4120 10124
rect 4120 10104 4122 10124
rect 3698 9968 3754 10024
rect 4158 9988 4214 10024
rect 4158 9968 4160 9988
rect 4160 9968 4212 9988
rect 4212 9968 4214 9988
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 3422 8064 3478 8120
rect 3514 7656 3570 7712
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3882 8492 3938 8528
rect 3882 8472 3884 8492
rect 3884 8472 3936 8492
rect 3936 8472 3938 8492
rect 3882 7792 3938 7848
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3698 7384 3754 7440
rect 3422 7248 3478 7304
rect 3146 6704 3202 6760
rect 2686 4528 2742 4584
rect 2594 3712 2650 3768
rect 2870 3848 2926 3904
rect 3238 5616 3294 5672
rect 4066 6840 4122 6896
rect 4618 12144 4674 12200
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 4618 10376 4674 10432
rect 4710 8880 4766 8936
rect 4618 7948 4674 7984
rect 4618 7928 4620 7948
rect 4620 7928 4672 7948
rect 4672 7928 4674 7948
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 4434 6160 4490 6216
rect 4158 5752 4214 5808
rect 3330 4256 3386 4312
rect 2502 3476 2504 3496
rect 2504 3476 2556 3496
rect 2556 3476 2558 3496
rect 2502 3440 2558 3476
rect 2226 3032 2282 3088
rect 1858 1808 1914 1864
rect 2318 2760 2374 2816
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3882 4684 3938 4720
rect 3882 4664 3884 4684
rect 3884 4664 3936 4684
rect 3936 4664 3938 4684
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3698 3848 3754 3904
rect 5722 10648 5778 10704
rect 5630 10240 5686 10296
rect 5814 10240 5870 10296
rect 4894 9560 4950 9616
rect 6182 12164 6238 12200
rect 6182 12144 6184 12164
rect 6184 12144 6236 12164
rect 6236 12144 6238 12164
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6734 12144 6790 12200
rect 6550 11600 6606 11656
rect 6458 11092 6460 11112
rect 6460 11092 6512 11112
rect 6512 11092 6514 11112
rect 6458 11056 6514 11092
rect 6274 10648 6330 10704
rect 4986 9288 5042 9344
rect 4802 5208 4858 5264
rect 4618 4528 4674 4584
rect 4342 3848 4398 3904
rect 3698 3168 3754 3224
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 4434 3440 4490 3496
rect 2778 2624 2834 2680
rect 2226 1400 2282 1456
rect 1766 584 1822 640
rect 5446 6976 5502 7032
rect 5906 9424 5962 9480
rect 6274 9288 6330 9344
rect 6458 9016 6514 9072
rect 6090 8880 6146 8936
rect 6458 8916 6460 8936
rect 6460 8916 6512 8936
rect 6512 8916 6514 8936
rect 6458 8880 6514 8916
rect 6182 8336 6238 8392
rect 6090 7520 6146 7576
rect 4986 4528 5042 4584
rect 5170 4664 5226 4720
rect 5538 4564 5540 4584
rect 5540 4564 5592 4584
rect 5592 4564 5594 4584
rect 5538 4528 5594 4564
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 5538 4020 5540 4040
rect 5540 4020 5592 4040
rect 5592 4020 5594 4040
rect 5538 3984 5594 4020
rect 5354 3440 5410 3496
rect 5722 3576 5778 3632
rect 5814 3032 5870 3088
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 7746 11872 7802 11928
rect 8114 11328 8170 11384
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 6826 8336 6882 8392
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6826 7928 6882 7984
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6090 3848 6146 3904
rect 6182 3576 6238 3632
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 7378 8744 7434 8800
rect 7378 7384 7434 7440
rect 7654 7268 7710 7304
rect 7654 7248 7656 7268
rect 7656 7248 7708 7268
rect 7708 7248 7710 7268
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6734 3712 6790 3768
rect 6734 2760 6790 2816
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 8390 10104 8446 10160
rect 8298 9424 8354 9480
rect 7930 8472 7986 8528
rect 8206 9016 8262 9072
rect 8482 8780 8484 8800
rect 8484 8780 8536 8800
rect 8536 8780 8538 8800
rect 8114 8064 8170 8120
rect 8482 8744 8538 8780
rect 8114 5788 8116 5808
rect 8116 5788 8168 5808
rect 8168 5788 8170 5808
rect 8114 5752 8170 5788
rect 8298 7248 8354 7304
rect 8482 7520 8538 7576
rect 8942 11892 8998 11928
rect 8942 11872 8944 11892
rect 8944 11872 8996 11892
rect 8996 11872 8998 11892
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 8390 6840 8446 6896
rect 8482 5616 8538 5672
rect 8390 5208 8446 5264
rect 8482 4564 8484 4584
rect 8484 4564 8536 4584
rect 8536 4564 8538 4584
rect 8482 4528 8538 4564
rect 9126 8064 9182 8120
rect 9586 12164 9642 12200
rect 9586 12144 9588 12164
rect 9588 12144 9640 12164
rect 9640 12144 9642 12164
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10230 11872 10286 11928
rect 9402 10648 9458 10704
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10322 10140 10324 10160
rect 10324 10140 10376 10160
rect 10376 10140 10378 10160
rect 10322 10104 10378 10140
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9954 9424 10010 9480
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9310 5208 9366 5264
rect 9034 3732 9090 3768
rect 9034 3712 9036 3732
rect 9036 3712 9088 3732
rect 9088 3712 9090 3732
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9586 3576 9642 3632
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10874 12144 10930 12200
rect 10690 11464 10746 11520
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 16394 15544 16450 15600
rect 15198 14340 15254 14376
rect 15198 14320 15200 14340
rect 15200 14320 15252 14340
rect 15252 14320 15254 14340
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 11334 11872 11390 11928
rect 11242 11500 11244 11520
rect 11244 11500 11296 11520
rect 11296 11500 11298 11520
rect 11242 11464 11298 11500
rect 11242 11192 11298 11248
rect 11058 10548 11060 10568
rect 11060 10548 11112 10568
rect 11112 10548 11114 10568
rect 11058 10512 11114 10548
rect 11058 9596 11060 9616
rect 11060 9596 11112 9616
rect 11112 9596 11114 9616
rect 11058 9560 11114 9596
rect 11150 8880 11206 8936
rect 11058 7384 11114 7440
rect 12530 12144 12586 12200
rect 12162 11872 12218 11928
rect 11886 11772 11888 11792
rect 11888 11772 11940 11792
rect 11940 11772 11942 11792
rect 11886 11736 11942 11772
rect 11426 7792 11482 7848
rect 11058 6196 11060 6216
rect 11060 6196 11112 6216
rect 11112 6196 11114 6216
rect 11058 6160 11114 6196
rect 11150 5888 11206 5944
rect 10782 5072 10838 5128
rect 10690 4120 10746 4176
rect 10506 3440 10562 3496
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10966 4664 11022 4720
rect 10966 3984 11022 4040
rect 10874 3732 10930 3768
rect 10874 3712 10876 3732
rect 10876 3712 10928 3732
rect 10928 3712 10930 3732
rect 10874 3168 10930 3224
rect 11518 5888 11574 5944
rect 10414 2644 10470 2680
rect 10414 2624 10416 2644
rect 10416 2624 10468 2644
rect 10468 2624 10470 2644
rect 11242 3304 11298 3360
rect 12254 11636 12256 11656
rect 12256 11636 12308 11656
rect 12308 11636 12310 11656
rect 12254 11600 12310 11636
rect 12622 11212 12678 11248
rect 12070 9968 12126 10024
rect 12070 9424 12126 9480
rect 11978 9016 12034 9072
rect 11610 4392 11666 4448
rect 12162 6296 12218 6352
rect 12346 5752 12402 5808
rect 12254 4820 12310 4856
rect 12254 4800 12256 4820
rect 12256 4800 12308 4820
rect 12308 4800 12310 4820
rect 12070 3032 12126 3088
rect 12622 11192 12624 11212
rect 12624 11192 12676 11212
rect 12676 11192 12678 11212
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12530 9424 12586 9480
rect 13450 11736 13506 11792
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12622 7268 12678 7304
rect 12622 7248 12624 7268
rect 12624 7248 12676 7268
rect 12676 7248 12678 7268
rect 13818 10104 13874 10160
rect 13542 9424 13598 9480
rect 13450 9324 13452 9344
rect 13452 9324 13504 9344
rect 13504 9324 13506 9344
rect 13450 9288 13506 9324
rect 13634 9016 13690 9072
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 13266 3440 13322 3496
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 13818 8880 13874 8936
rect 14002 11872 14058 11928
rect 14278 11600 14334 11656
rect 14002 11056 14058 11112
rect 13450 5092 13506 5128
rect 13450 5072 13452 5092
rect 13452 5072 13504 5092
rect 13504 5072 13506 5092
rect 13818 6860 13874 6896
rect 13818 6840 13820 6860
rect 13820 6840 13872 6860
rect 13872 6840 13874 6860
rect 13818 6296 13874 6352
rect 13818 5752 13874 5808
rect 14094 8880 14150 8936
rect 14922 12824 14978 12880
rect 14830 12144 14886 12200
rect 15290 13368 15346 13424
rect 15566 13368 15622 13424
rect 15382 13252 15438 13288
rect 15382 13232 15384 13252
rect 15384 13232 15436 13252
rect 15436 13232 15438 13252
rect 14370 7248 14426 7304
rect 14094 4664 14150 4720
rect 13910 3984 13966 4040
rect 14370 6160 14426 6216
rect 14186 3032 14242 3088
rect 14922 8916 14924 8936
rect 14924 8916 14976 8936
rect 14976 8916 14978 8936
rect 14922 8880 14978 8916
rect 14830 8336 14886 8392
rect 14830 6840 14886 6896
rect 15198 5072 15254 5128
rect 15198 4936 15254 4992
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15566 9968 15622 10024
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 17774 16360 17830 16416
rect 17682 15136 17738 15192
rect 16210 12824 16266 12880
rect 15474 5752 15530 5808
rect 15566 3304 15622 3360
rect 15934 7384 15990 7440
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 16394 13368 16450 13424
rect 16578 12416 16634 12472
rect 16578 11636 16580 11656
rect 16580 11636 16632 11656
rect 16632 11636 16634 11656
rect 16578 11600 16634 11636
rect 17130 12416 17186 12472
rect 17038 11736 17094 11792
rect 16486 10784 16542 10840
rect 16394 9716 16450 9752
rect 16394 9696 16396 9716
rect 16396 9696 16448 9716
rect 16448 9696 16450 9716
rect 16394 9324 16396 9344
rect 16396 9324 16448 9344
rect 16448 9324 16450 9344
rect 16394 9288 16450 9324
rect 16762 10648 16818 10704
rect 17130 11328 17186 11384
rect 16394 4120 16450 4176
rect 16486 3576 16542 3632
rect 17130 9716 17186 9752
rect 17130 9696 17132 9716
rect 17132 9696 17184 9716
rect 17184 9696 17186 9716
rect 17866 15952 17922 16008
rect 18050 14728 18106 14784
rect 17682 13232 17738 13288
rect 17682 12552 17738 12608
rect 17406 11600 17462 11656
rect 18418 14184 18474 14240
rect 18418 13812 18420 13832
rect 18420 13812 18472 13832
rect 18472 13812 18474 13832
rect 18418 13776 18474 13812
rect 18418 13388 18474 13424
rect 18418 13368 18420 13388
rect 18420 13368 18472 13388
rect 18472 13368 18474 13388
rect 18510 12960 18566 13016
rect 18050 12144 18106 12200
rect 17038 7792 17094 7848
rect 17866 9424 17922 9480
rect 17866 8372 17868 8392
rect 17868 8372 17920 8392
rect 17920 8372 17922 8392
rect 17866 8336 17922 8372
rect 17958 8200 18014 8256
rect 17958 7812 18014 7848
rect 17958 7792 17960 7812
rect 17960 7792 18012 7812
rect 18012 7792 18014 7812
rect 17866 7284 17868 7304
rect 17868 7284 17920 7304
rect 17920 7284 17922 7304
rect 17866 7248 17922 7284
rect 18142 6976 18198 7032
rect 18142 4800 18198 4856
rect 18142 4004 18198 4040
rect 18142 3984 18144 4004
rect 18144 3984 18196 4004
rect 18196 3984 18198 4004
rect 17038 3032 17094 3088
rect 16118 2896 16174 2952
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16578 992 16634 1048
rect 3330 176 3386 232
rect 17590 1808 17646 1864
rect 17774 2624 17830 2680
rect 18142 3168 18198 3224
rect 18970 12144 19026 12200
rect 18970 11228 18972 11248
rect 18972 11228 19024 11248
rect 19024 11228 19026 11248
rect 18970 11192 19026 11228
rect 18510 10376 18566 10432
rect 18602 9968 18658 10024
rect 18602 9560 18658 9616
rect 18510 9152 18566 9208
rect 18418 8744 18474 8800
rect 18510 7404 18566 7440
rect 18510 7384 18512 7404
rect 18512 7384 18564 7404
rect 18564 7384 18566 7404
rect 18510 6568 18566 6624
rect 18510 6180 18566 6216
rect 18510 6160 18512 6180
rect 18512 6160 18564 6180
rect 18564 6160 18566 6180
rect 18510 5636 18566 5672
rect 18510 5616 18512 5636
rect 18512 5616 18564 5636
rect 18564 5616 18566 5636
rect 18510 5228 18566 5264
rect 18510 5208 18512 5228
rect 18512 5208 18564 5228
rect 18564 5208 18566 5228
rect 18510 4392 18566 4448
rect 18510 3576 18566 3632
rect 17682 1400 17738 1456
rect 17498 584 17554 640
rect 17866 2216 17922 2272
rect 17774 176 17830 232
<< metal3 >>
rect 0 16826 800 16856
rect 3509 16826 3575 16829
rect 0 16824 3575 16826
rect 0 16768 3514 16824
rect 3570 16768 3575 16824
rect 0 16766 3575 16768
rect 0 16736 800 16766
rect 3509 16763 3575 16766
rect 16481 16826 16547 16829
rect 19200 16826 20000 16856
rect 16481 16824 20000 16826
rect 16481 16768 16486 16824
rect 16542 16768 20000 16824
rect 16481 16766 20000 16768
rect 16481 16763 16547 16766
rect 19200 16736 20000 16766
rect 0 16418 800 16448
rect 3049 16418 3115 16421
rect 0 16416 3115 16418
rect 0 16360 3054 16416
rect 3110 16360 3115 16416
rect 0 16358 3115 16360
rect 0 16328 800 16358
rect 3049 16355 3115 16358
rect 17769 16418 17835 16421
rect 19200 16418 20000 16448
rect 17769 16416 20000 16418
rect 17769 16360 17774 16416
rect 17830 16360 20000 16416
rect 17769 16358 20000 16360
rect 17769 16355 17835 16358
rect 19200 16328 20000 16358
rect 0 16010 800 16040
rect 2957 16010 3023 16013
rect 0 16008 3023 16010
rect 0 15952 2962 16008
rect 3018 15952 3023 16008
rect 0 15950 3023 15952
rect 0 15920 800 15950
rect 2957 15947 3023 15950
rect 17861 16010 17927 16013
rect 19200 16010 20000 16040
rect 17861 16008 20000 16010
rect 17861 15952 17866 16008
rect 17922 15952 20000 16008
rect 17861 15950 20000 15952
rect 17861 15947 17927 15950
rect 19200 15920 20000 15950
rect 0 15602 800 15632
rect 2497 15602 2563 15605
rect 0 15600 2563 15602
rect 0 15544 2502 15600
rect 2558 15544 2563 15600
rect 0 15542 2563 15544
rect 0 15512 800 15542
rect 2497 15539 2563 15542
rect 16389 15602 16455 15605
rect 19200 15602 20000 15632
rect 16389 15600 20000 15602
rect 16389 15544 16394 15600
rect 16450 15544 20000 15600
rect 16389 15542 20000 15544
rect 16389 15539 16455 15542
rect 19200 15512 20000 15542
rect 0 15194 800 15224
rect 2221 15194 2287 15197
rect 0 15192 2287 15194
rect 0 15136 2226 15192
rect 2282 15136 2287 15192
rect 0 15134 2287 15136
rect 0 15104 800 15134
rect 2221 15131 2287 15134
rect 17677 15194 17743 15197
rect 19200 15194 20000 15224
rect 17677 15192 20000 15194
rect 17677 15136 17682 15192
rect 17738 15136 20000 15192
rect 17677 15134 20000 15136
rect 17677 15131 17743 15134
rect 19200 15104 20000 15134
rect 0 14786 800 14816
rect 1853 14786 1919 14789
rect 0 14784 1919 14786
rect 0 14728 1858 14784
rect 1914 14728 1919 14784
rect 0 14726 1919 14728
rect 0 14696 800 14726
rect 1853 14723 1919 14726
rect 18045 14786 18111 14789
rect 19200 14786 20000 14816
rect 18045 14784 20000 14786
rect 18045 14728 18050 14784
rect 18106 14728 20000 14784
rect 18045 14726 20000 14728
rect 18045 14723 18111 14726
rect 6874 14720 7194 14721
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 19200 14696 20000 14726
rect 12805 14655 13125 14656
rect 2221 14514 2287 14517
rect 3601 14514 3667 14517
rect 2221 14512 3667 14514
rect 2221 14456 2226 14512
rect 2282 14456 3606 14512
rect 3662 14456 3667 14512
rect 2221 14454 3667 14456
rect 2221 14451 2287 14454
rect 3601 14451 3667 14454
rect 0 14378 800 14408
rect 1485 14378 1551 14381
rect 0 14376 1551 14378
rect 0 14320 1490 14376
rect 1546 14320 1551 14376
rect 0 14318 1551 14320
rect 0 14288 800 14318
rect 1485 14315 1551 14318
rect 15193 14378 15259 14381
rect 15193 14376 17418 14378
rect 15193 14320 15198 14376
rect 15254 14320 17418 14376
rect 15193 14318 17418 14320
rect 15193 14315 15259 14318
rect 17358 14242 17418 14318
rect 18413 14242 18479 14245
rect 19200 14242 20000 14272
rect 17358 14240 20000 14242
rect 17358 14184 18418 14240
rect 18474 14184 20000 14240
rect 17358 14182 20000 14184
rect 18413 14179 18479 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13970 800 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 800 13910
rect 1485 13907 1551 13910
rect 1669 13970 1735 13973
rect 5625 13970 5691 13973
rect 1669 13968 5691 13970
rect 1669 13912 1674 13968
rect 1730 13912 5630 13968
rect 5686 13912 5691 13968
rect 1669 13910 5691 13912
rect 1669 13907 1735 13910
rect 5625 13907 5691 13910
rect 18413 13834 18479 13837
rect 19200 13834 20000 13864
rect 18413 13832 20000 13834
rect 18413 13776 18418 13832
rect 18474 13776 20000 13832
rect 18413 13774 20000 13776
rect 18413 13771 18479 13774
rect 19200 13744 20000 13774
rect 6874 13632 7194 13633
rect 0 13562 800 13592
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 1853 13562 1919 13565
rect 0 13560 1919 13562
rect 0 13504 1858 13560
rect 1914 13504 1919 13560
rect 0 13502 1919 13504
rect 0 13472 800 13502
rect 1853 13499 1919 13502
rect 15285 13426 15351 13429
rect 15561 13426 15627 13429
rect 16389 13426 16455 13429
rect 15285 13424 16455 13426
rect 15285 13368 15290 13424
rect 15346 13368 15566 13424
rect 15622 13368 16394 13424
rect 16450 13368 16455 13424
rect 15285 13366 16455 13368
rect 15285 13363 15351 13366
rect 15561 13363 15627 13366
rect 16389 13363 16455 13366
rect 18413 13426 18479 13429
rect 19200 13426 20000 13456
rect 18413 13424 20000 13426
rect 18413 13368 18418 13424
rect 18474 13368 20000 13424
rect 18413 13366 20000 13368
rect 18413 13363 18479 13366
rect 19200 13336 20000 13366
rect 15377 13290 15443 13293
rect 17677 13290 17743 13293
rect 15377 13288 17743 13290
rect 15377 13232 15382 13288
rect 15438 13232 17682 13288
rect 17738 13232 17743 13288
rect 15377 13230 17743 13232
rect 15377 13227 15443 13230
rect 17677 13227 17743 13230
rect 0 13154 800 13184
rect 1485 13154 1551 13157
rect 0 13152 1551 13154
rect 0 13096 1490 13152
rect 1546 13096 1551 13152
rect 0 13094 1551 13096
rect 0 13064 800 13094
rect 1485 13091 1551 13094
rect 3909 13088 4229 13089
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 18505 13018 18571 13021
rect 19200 13018 20000 13048
rect 18505 13016 20000 13018
rect 18505 12960 18510 13016
rect 18566 12960 20000 13016
rect 18505 12958 20000 12960
rect 18505 12955 18571 12958
rect 19200 12928 20000 12958
rect 14917 12882 14983 12885
rect 16205 12882 16271 12885
rect 14917 12880 16271 12882
rect 14917 12824 14922 12880
rect 14978 12824 16210 12880
rect 16266 12824 16271 12880
rect 14917 12822 16271 12824
rect 14917 12819 14983 12822
rect 16205 12819 16271 12822
rect 0 12746 800 12776
rect 1853 12746 1919 12749
rect 0 12744 1919 12746
rect 0 12688 1858 12744
rect 1914 12688 1919 12744
rect 0 12686 1919 12688
rect 0 12656 800 12686
rect 1853 12683 1919 12686
rect 17677 12610 17743 12613
rect 19200 12610 20000 12640
rect 17677 12608 20000 12610
rect 17677 12552 17682 12608
rect 17738 12552 20000 12608
rect 17677 12550 20000 12552
rect 17677 12547 17743 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 19200 12520 20000 12550
rect 12805 12479 13125 12480
rect 16573 12474 16639 12477
rect 17125 12474 17191 12477
rect 16573 12472 17191 12474
rect 16573 12416 16578 12472
rect 16634 12416 17130 12472
rect 17186 12416 17191 12472
rect 16573 12414 17191 12416
rect 16573 12411 16639 12414
rect 17125 12411 17191 12414
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 3877 12202 3943 12205
rect 4613 12202 4679 12205
rect 6177 12202 6243 12205
rect 3877 12200 6243 12202
rect 3877 12144 3882 12200
rect 3938 12144 4618 12200
rect 4674 12144 6182 12200
rect 6238 12144 6243 12200
rect 3877 12142 6243 12144
rect 3877 12139 3943 12142
rect 4613 12139 4679 12142
rect 6177 12139 6243 12142
rect 6729 12202 6795 12205
rect 9581 12202 9647 12205
rect 6729 12200 9647 12202
rect 6729 12144 6734 12200
rect 6790 12144 9586 12200
rect 9642 12144 9647 12200
rect 6729 12142 9647 12144
rect 6729 12139 6795 12142
rect 9581 12139 9647 12142
rect 10869 12202 10935 12205
rect 12525 12202 12591 12205
rect 10869 12200 12591 12202
rect 10869 12144 10874 12200
rect 10930 12144 12530 12200
rect 12586 12144 12591 12200
rect 10869 12142 12591 12144
rect 10869 12139 10935 12142
rect 12525 12139 12591 12142
rect 14825 12202 14891 12205
rect 18045 12202 18111 12205
rect 14825 12200 18111 12202
rect 14825 12144 14830 12200
rect 14886 12144 18050 12200
rect 18106 12144 18111 12200
rect 14825 12142 18111 12144
rect 14825 12139 14891 12142
rect 18045 12139 18111 12142
rect 18965 12202 19031 12205
rect 19200 12202 20000 12232
rect 18965 12200 20000 12202
rect 18965 12144 18970 12200
rect 19026 12144 20000 12200
rect 18965 12142 20000 12144
rect 18965 12139 19031 12142
rect 19200 12112 20000 12142
rect 3909 12000 4229 12001
rect 0 11930 800 11960
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 2221 11930 2287 11933
rect 0 11928 2287 11930
rect 0 11872 2226 11928
rect 2282 11872 2287 11928
rect 0 11870 2287 11872
rect 0 11840 800 11870
rect 2221 11867 2287 11870
rect 7741 11930 7807 11933
rect 8937 11930 9003 11933
rect 7741 11928 9003 11930
rect 7741 11872 7746 11928
rect 7802 11872 8942 11928
rect 8998 11872 9003 11928
rect 7741 11870 9003 11872
rect 7741 11867 7807 11870
rect 8937 11867 9003 11870
rect 10225 11930 10291 11933
rect 11329 11930 11395 11933
rect 12157 11930 12223 11933
rect 13997 11930 14063 11933
rect 10225 11928 14063 11930
rect 10225 11872 10230 11928
rect 10286 11872 11334 11928
rect 11390 11872 12162 11928
rect 12218 11872 14002 11928
rect 14058 11872 14063 11928
rect 10225 11870 14063 11872
rect 10225 11867 10291 11870
rect 11329 11867 11395 11870
rect 12157 11867 12223 11870
rect 13997 11867 14063 11870
rect 11881 11794 11947 11797
rect 13445 11794 13511 11797
rect 11881 11792 13511 11794
rect 11881 11736 11886 11792
rect 11942 11736 13450 11792
rect 13506 11736 13511 11792
rect 11881 11734 13511 11736
rect 11881 11731 11947 11734
rect 13445 11731 13511 11734
rect 17033 11794 17099 11797
rect 19200 11794 20000 11824
rect 17033 11792 20000 11794
rect 17033 11736 17038 11792
rect 17094 11736 20000 11792
rect 17033 11734 20000 11736
rect 17033 11731 17099 11734
rect 19200 11704 20000 11734
rect 6545 11658 6611 11661
rect 12249 11658 12315 11661
rect 14273 11658 14339 11661
rect 16573 11658 16639 11661
rect 17401 11658 17467 11661
rect 6545 11656 12315 11658
rect 6545 11600 6550 11656
rect 6606 11600 12254 11656
rect 12310 11600 12315 11656
rect 6545 11598 12315 11600
rect 6545 11595 6611 11598
rect 12249 11595 12315 11598
rect 12620 11656 16639 11658
rect 12620 11600 14278 11656
rect 14334 11600 16578 11656
rect 16634 11600 16639 11656
rect 12620 11598 16639 11600
rect 10685 11522 10751 11525
rect 11237 11522 11303 11525
rect 12620 11522 12680 11598
rect 14273 11595 14339 11598
rect 16573 11595 16639 11598
rect 17174 11656 17467 11658
rect 17174 11600 17406 11656
rect 17462 11600 17467 11656
rect 17174 11598 17467 11600
rect 9630 11520 12680 11522
rect 9630 11464 10690 11520
rect 10746 11464 11242 11520
rect 11298 11464 12680 11520
rect 9630 11462 12680 11464
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 1393 11386 1459 11389
rect 0 11384 1459 11386
rect 0 11328 1398 11384
rect 1454 11328 1459 11384
rect 0 11326 1459 11328
rect 0 11296 800 11326
rect 1393 11323 1459 11326
rect 8109 11386 8175 11389
rect 9630 11386 9690 11462
rect 10685 11459 10751 11462
rect 11237 11459 11303 11462
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 17174 11389 17234 11598
rect 17401 11595 17467 11598
rect 8109 11384 9690 11386
rect 8109 11328 8114 11384
rect 8170 11328 9690 11384
rect 8109 11326 9690 11328
rect 17125 11384 17234 11389
rect 17125 11328 17130 11384
rect 17186 11328 17234 11384
rect 17125 11326 17234 11328
rect 8109 11323 8175 11326
rect 17125 11323 17191 11326
rect 11237 11250 11303 11253
rect 12617 11250 12683 11253
rect 11237 11248 12683 11250
rect 11237 11192 11242 11248
rect 11298 11192 12622 11248
rect 12678 11192 12683 11248
rect 11237 11190 12683 11192
rect 11237 11187 11303 11190
rect 12617 11187 12683 11190
rect 18965 11250 19031 11253
rect 19200 11250 20000 11280
rect 18965 11248 20000 11250
rect 18965 11192 18970 11248
rect 19026 11192 20000 11248
rect 18965 11190 20000 11192
rect 18965 11187 19031 11190
rect 19200 11160 20000 11190
rect 6453 11114 6519 11117
rect 13997 11114 14063 11117
rect 6453 11112 14063 11114
rect 6453 11056 6458 11112
rect 6514 11056 14002 11112
rect 14058 11056 14063 11112
rect 6453 11054 14063 11056
rect 6453 11051 6519 11054
rect 13997 11051 14063 11054
rect 0 10978 800 11008
rect 2037 10978 2103 10981
rect 0 10976 2103 10978
rect 0 10920 2042 10976
rect 2098 10920 2103 10976
rect 0 10918 2103 10920
rect 0 10888 800 10918
rect 2037 10915 2103 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 16481 10842 16547 10845
rect 19200 10842 20000 10872
rect 16481 10840 20000 10842
rect 16481 10784 16486 10840
rect 16542 10784 20000 10840
rect 16481 10782 20000 10784
rect 16481 10779 16547 10782
rect 19200 10752 20000 10782
rect 1669 10706 1735 10709
rect 5717 10706 5783 10709
rect 6269 10706 6335 10709
rect 1669 10704 6335 10706
rect 1669 10648 1674 10704
rect 1730 10648 5722 10704
rect 5778 10648 6274 10704
rect 6330 10648 6335 10704
rect 1669 10646 6335 10648
rect 1669 10643 1735 10646
rect 5717 10643 5783 10646
rect 6269 10643 6335 10646
rect 9397 10706 9463 10709
rect 16757 10706 16823 10709
rect 9397 10704 16823 10706
rect 9397 10648 9402 10704
rect 9458 10648 16762 10704
rect 16818 10648 16823 10704
rect 9397 10646 16823 10648
rect 9397 10643 9463 10646
rect 16757 10643 16823 10646
rect 0 10570 800 10600
rect 2865 10570 2931 10573
rect 0 10568 2931 10570
rect 0 10512 2870 10568
rect 2926 10512 2931 10568
rect 0 10510 2931 10512
rect 0 10480 800 10510
rect 2865 10507 2931 10510
rect 3049 10570 3115 10573
rect 11053 10570 11119 10573
rect 3049 10568 11119 10570
rect 3049 10512 3054 10568
rect 3110 10512 11058 10568
rect 11114 10512 11119 10568
rect 3049 10510 11119 10512
rect 3049 10507 3115 10510
rect 11053 10507 11119 10510
rect 1853 10434 1919 10437
rect 4613 10434 4679 10437
rect 1853 10432 4679 10434
rect 1853 10376 1858 10432
rect 1914 10376 4618 10432
rect 4674 10376 4679 10432
rect 1853 10374 4679 10376
rect 1853 10371 1919 10374
rect 4613 10371 4679 10374
rect 18505 10434 18571 10437
rect 19200 10434 20000 10464
rect 18505 10432 20000 10434
rect 18505 10376 18510 10432
rect 18566 10376 20000 10432
rect 18505 10374 20000 10376
rect 18505 10371 18571 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 3601 10298 3667 10301
rect 5625 10298 5691 10301
rect 5809 10298 5875 10301
rect 3601 10296 5691 10298
rect 3601 10240 3606 10296
rect 3662 10240 5630 10296
rect 5686 10240 5691 10296
rect 3601 10238 5691 10240
rect 3601 10235 3667 10238
rect 5625 10235 5691 10238
rect 5766 10296 5875 10298
rect 5766 10240 5814 10296
rect 5870 10240 5875 10296
rect 5766 10235 5875 10240
rect 0 10162 800 10192
rect 1761 10162 1827 10165
rect 0 10160 1827 10162
rect 0 10104 1766 10160
rect 1822 10104 1827 10160
rect 0 10102 1827 10104
rect 0 10072 800 10102
rect 1761 10099 1827 10102
rect 4061 10162 4127 10165
rect 5766 10162 5826 10235
rect 8385 10162 8451 10165
rect 4061 10160 8451 10162
rect 4061 10104 4066 10160
rect 4122 10104 8390 10160
rect 8446 10104 8451 10160
rect 4061 10102 8451 10104
rect 4061 10099 4127 10102
rect 8385 10099 8451 10102
rect 10317 10162 10383 10165
rect 13813 10162 13879 10165
rect 10317 10160 13879 10162
rect 10317 10104 10322 10160
rect 10378 10104 13818 10160
rect 13874 10104 13879 10160
rect 10317 10102 13879 10104
rect 10317 10099 10383 10102
rect 13813 10099 13879 10102
rect 2313 10026 2379 10029
rect 3693 10026 3759 10029
rect 4153 10026 4219 10029
rect 2313 10024 4219 10026
rect 2313 9968 2318 10024
rect 2374 9968 3698 10024
rect 3754 9968 4158 10024
rect 4214 9968 4219 10024
rect 2313 9966 4219 9968
rect 2313 9963 2379 9966
rect 3693 9963 3759 9966
rect 4153 9963 4219 9966
rect 12065 10026 12131 10029
rect 15561 10026 15627 10029
rect 12065 10024 15627 10026
rect 12065 9968 12070 10024
rect 12126 9968 15566 10024
rect 15622 9968 15627 10024
rect 12065 9966 15627 9968
rect 12065 9963 12131 9966
rect 15561 9963 15627 9966
rect 18597 10026 18663 10029
rect 19200 10026 20000 10056
rect 18597 10024 20000 10026
rect 18597 9968 18602 10024
rect 18658 9968 20000 10024
rect 18597 9966 20000 9968
rect 18597 9963 18663 9966
rect 19200 9936 20000 9966
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 9759 16090 9760
rect 3325 9754 3391 9757
rect 0 9752 3391 9754
rect 0 9696 3330 9752
rect 3386 9696 3391 9752
rect 0 9694 3391 9696
rect 0 9664 800 9694
rect 3325 9691 3391 9694
rect 16389 9754 16455 9757
rect 17125 9754 17191 9757
rect 16389 9752 17191 9754
rect 16389 9696 16394 9752
rect 16450 9696 17130 9752
rect 17186 9696 17191 9752
rect 16389 9694 17191 9696
rect 16389 9691 16455 9694
rect 17125 9691 17191 9694
rect 4889 9618 4955 9621
rect 11053 9618 11119 9621
rect 4889 9616 11119 9618
rect 4889 9560 4894 9616
rect 4950 9560 11058 9616
rect 11114 9560 11119 9616
rect 4889 9558 11119 9560
rect 4889 9555 4955 9558
rect 11053 9555 11119 9558
rect 18597 9618 18663 9621
rect 19200 9618 20000 9648
rect 18597 9616 20000 9618
rect 18597 9560 18602 9616
rect 18658 9560 20000 9616
rect 18597 9558 20000 9560
rect 18597 9555 18663 9558
rect 19200 9528 20000 9558
rect 5901 9482 5967 9485
rect 8293 9482 8359 9485
rect 5901 9480 8359 9482
rect 5901 9424 5906 9480
rect 5962 9424 8298 9480
rect 8354 9424 8359 9480
rect 5901 9422 8359 9424
rect 5901 9419 5967 9422
rect 8293 9419 8359 9422
rect 9949 9482 10015 9485
rect 12065 9482 12131 9485
rect 12198 9482 12204 9484
rect 9949 9480 12204 9482
rect 9949 9424 9954 9480
rect 10010 9424 12070 9480
rect 12126 9424 12204 9480
rect 9949 9422 12204 9424
rect 9949 9419 10015 9422
rect 12065 9419 12131 9422
rect 12198 9420 12204 9422
rect 12268 9482 12274 9484
rect 12525 9482 12591 9485
rect 13537 9482 13603 9485
rect 17861 9482 17927 9485
rect 12268 9480 17927 9482
rect 12268 9424 12530 9480
rect 12586 9424 13542 9480
rect 13598 9424 17866 9480
rect 17922 9424 17927 9480
rect 12268 9422 17927 9424
rect 12268 9420 12274 9422
rect 12525 9419 12591 9422
rect 13537 9419 13603 9422
rect 17861 9419 17927 9422
rect 0 9346 800 9376
rect 3141 9346 3207 9349
rect 0 9344 3207 9346
rect 0 9288 3146 9344
rect 3202 9288 3207 9344
rect 0 9286 3207 9288
rect 0 9256 800 9286
rect 3141 9283 3207 9286
rect 4981 9346 5047 9349
rect 6269 9346 6335 9349
rect 4981 9344 6335 9346
rect 4981 9288 4986 9344
rect 5042 9288 6274 9344
rect 6330 9288 6335 9344
rect 4981 9286 6335 9288
rect 4981 9283 5047 9286
rect 6269 9283 6335 9286
rect 13445 9346 13511 9349
rect 16389 9346 16455 9349
rect 13445 9344 16455 9346
rect 13445 9288 13450 9344
rect 13506 9288 16394 9344
rect 16450 9288 16455 9344
rect 13445 9286 16455 9288
rect 13445 9283 13511 9286
rect 16389 9283 16455 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 18505 9210 18571 9213
rect 19200 9210 20000 9240
rect 18505 9208 20000 9210
rect 18505 9152 18510 9208
rect 18566 9152 20000 9208
rect 18505 9150 20000 9152
rect 18505 9147 18571 9150
rect 19200 9120 20000 9150
rect 6453 9074 6519 9077
rect 8201 9074 8267 9077
rect 6453 9072 8267 9074
rect 6453 9016 6458 9072
rect 6514 9016 8206 9072
rect 8262 9016 8267 9072
rect 6453 9014 8267 9016
rect 6453 9011 6519 9014
rect 8201 9011 8267 9014
rect 11973 9074 12039 9077
rect 13629 9074 13695 9077
rect 11973 9072 13695 9074
rect 11973 9016 11978 9072
rect 12034 9016 13634 9072
rect 13690 9016 13695 9072
rect 11973 9014 13695 9016
rect 11973 9011 12039 9014
rect 13629 9011 13695 9014
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 4705 8938 4771 8941
rect 6085 8938 6151 8941
rect 6453 8938 6519 8941
rect 4705 8936 6519 8938
rect 4705 8880 4710 8936
rect 4766 8880 6090 8936
rect 6146 8880 6458 8936
rect 6514 8880 6519 8936
rect 4705 8878 6519 8880
rect 4705 8875 4771 8878
rect 6085 8875 6151 8878
rect 6453 8875 6519 8878
rect 11145 8938 11211 8941
rect 13813 8938 13879 8941
rect 11145 8936 13879 8938
rect 11145 8880 11150 8936
rect 11206 8880 13818 8936
rect 13874 8880 13879 8936
rect 11145 8878 13879 8880
rect 11145 8875 11211 8878
rect 13813 8875 13879 8878
rect 14089 8938 14155 8941
rect 14917 8938 14983 8941
rect 14089 8936 14983 8938
rect 14089 8880 14094 8936
rect 14150 8880 14922 8936
rect 14978 8880 14983 8936
rect 14089 8878 14983 8880
rect 14089 8875 14155 8878
rect 14917 8875 14983 8878
rect 7373 8802 7439 8805
rect 8477 8802 8543 8805
rect 7373 8800 8543 8802
rect 7373 8744 7378 8800
rect 7434 8744 8482 8800
rect 8538 8744 8543 8800
rect 7373 8742 8543 8744
rect 7373 8739 7439 8742
rect 8477 8739 8543 8742
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 18413 8739 18479 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 19200 8712 20000 8742
rect 15770 8671 16090 8672
rect 0 8530 800 8560
rect 3049 8530 3115 8533
rect 0 8528 3115 8530
rect 0 8472 3054 8528
rect 3110 8472 3115 8528
rect 0 8470 3115 8472
rect 0 8440 800 8470
rect 3049 8467 3115 8470
rect 3877 8530 3943 8533
rect 7925 8530 7991 8533
rect 3877 8528 7991 8530
rect 3877 8472 3882 8528
rect 3938 8472 7930 8528
rect 7986 8472 7991 8528
rect 3877 8470 7991 8472
rect 3877 8467 3943 8470
rect 7925 8467 7991 8470
rect 6177 8394 6243 8397
rect 6821 8394 6887 8397
rect 6177 8392 6887 8394
rect 6177 8336 6182 8392
rect 6238 8336 6826 8392
rect 6882 8336 6887 8392
rect 6177 8334 6887 8336
rect 6177 8331 6243 8334
rect 6821 8331 6887 8334
rect 14825 8394 14891 8397
rect 17861 8394 17927 8397
rect 14825 8392 17927 8394
rect 14825 8336 14830 8392
rect 14886 8336 17866 8392
rect 17922 8336 17927 8392
rect 14825 8334 17927 8336
rect 14825 8331 14891 8334
rect 17861 8331 17927 8334
rect 17953 8258 18019 8261
rect 19200 8258 20000 8288
rect 17953 8256 20000 8258
rect 17953 8200 17958 8256
rect 18014 8200 20000 8256
rect 17953 8198 20000 8200
rect 17953 8195 18019 8198
rect 6874 8192 7194 8193
rect 0 8122 800 8152
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19200 8168 20000 8198
rect 12805 8127 13125 8128
rect 3417 8122 3483 8125
rect 0 8120 3483 8122
rect 0 8064 3422 8120
rect 3478 8064 3483 8120
rect 0 8062 3483 8064
rect 0 8032 800 8062
rect 3417 8059 3483 8062
rect 8109 8122 8175 8125
rect 9121 8122 9187 8125
rect 8109 8120 9187 8122
rect 8109 8064 8114 8120
rect 8170 8064 9126 8120
rect 9182 8064 9187 8120
rect 8109 8062 9187 8064
rect 8109 8059 8175 8062
rect 9121 8059 9187 8062
rect 4613 7986 4679 7989
rect 6821 7986 6887 7989
rect 4613 7984 6887 7986
rect 4613 7928 4618 7984
rect 4674 7928 6826 7984
rect 6882 7928 6887 7984
rect 4613 7926 6887 7928
rect 4613 7923 4679 7926
rect 6821 7923 6887 7926
rect 3877 7850 3943 7853
rect 3558 7848 3943 7850
rect 3558 7792 3882 7848
rect 3938 7792 3943 7848
rect 3558 7790 3943 7792
rect 0 7714 800 7744
rect 3558 7717 3618 7790
rect 3877 7787 3943 7790
rect 11421 7850 11487 7853
rect 17033 7850 17099 7853
rect 11421 7848 17099 7850
rect 11421 7792 11426 7848
rect 11482 7792 17038 7848
rect 17094 7792 17099 7848
rect 11421 7790 17099 7792
rect 11421 7787 11487 7790
rect 17033 7787 17099 7790
rect 17953 7850 18019 7853
rect 19200 7850 20000 7880
rect 17953 7848 20000 7850
rect 17953 7792 17958 7848
rect 18014 7792 20000 7848
rect 17953 7790 20000 7792
rect 17953 7787 18019 7790
rect 19200 7760 20000 7790
rect 2865 7714 2931 7717
rect 3509 7716 3618 7717
rect 3509 7714 3556 7716
rect 0 7712 2931 7714
rect 0 7656 2870 7712
rect 2926 7656 2931 7712
rect 0 7654 2931 7656
rect 3428 7712 3556 7714
rect 3428 7656 3514 7712
rect 3428 7654 3556 7656
rect 0 7624 800 7654
rect 2865 7651 2931 7654
rect 3509 7652 3556 7654
rect 3620 7652 3626 7716
rect 3509 7651 3575 7652
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 6085 7578 6151 7581
rect 8477 7578 8543 7581
rect 6085 7576 8543 7578
rect 6085 7520 6090 7576
rect 6146 7520 8482 7576
rect 8538 7520 8543 7576
rect 6085 7518 8543 7520
rect 6085 7515 6151 7518
rect 8477 7515 8543 7518
rect 3693 7442 3759 7445
rect 7373 7442 7439 7445
rect 3693 7440 7439 7442
rect 3693 7384 3698 7440
rect 3754 7384 7378 7440
rect 7434 7384 7439 7440
rect 3693 7382 7439 7384
rect 3693 7379 3759 7382
rect 7373 7379 7439 7382
rect 11053 7442 11119 7445
rect 15929 7442 15995 7445
rect 11053 7440 15995 7442
rect 11053 7384 11058 7440
rect 11114 7384 15934 7440
rect 15990 7384 15995 7440
rect 11053 7382 15995 7384
rect 11053 7379 11119 7382
rect 15929 7379 15995 7382
rect 18505 7442 18571 7445
rect 19200 7442 20000 7472
rect 18505 7440 20000 7442
rect 18505 7384 18510 7440
rect 18566 7384 20000 7440
rect 18505 7382 20000 7384
rect 18505 7379 18571 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 1485 7306 1551 7309
rect 0 7304 1551 7306
rect 0 7248 1490 7304
rect 1546 7248 1551 7304
rect 0 7246 1551 7248
rect 0 7216 800 7246
rect 1485 7243 1551 7246
rect 3417 7306 3483 7309
rect 7649 7306 7715 7309
rect 8293 7306 8359 7309
rect 3417 7304 8359 7306
rect 3417 7248 3422 7304
rect 3478 7248 7654 7304
rect 7710 7248 8298 7304
rect 8354 7248 8359 7304
rect 3417 7246 8359 7248
rect 3417 7243 3483 7246
rect 7649 7243 7715 7246
rect 8293 7243 8359 7246
rect 12617 7306 12683 7309
rect 14365 7306 14431 7309
rect 17861 7306 17927 7309
rect 12617 7304 17927 7306
rect 12617 7248 12622 7304
rect 12678 7248 14370 7304
rect 14426 7248 17866 7304
rect 17922 7248 17927 7304
rect 12617 7246 17927 7248
rect 12617 7243 12683 7246
rect 14365 7243 14431 7246
rect 17861 7243 17927 7246
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 2037 7034 2103 7037
rect 5441 7034 5507 7037
rect 2037 7032 5507 7034
rect 2037 6976 2042 7032
rect 2098 6976 5446 7032
rect 5502 6976 5507 7032
rect 2037 6974 5507 6976
rect 2037 6971 2103 6974
rect 5441 6971 5507 6974
rect 18137 7034 18203 7037
rect 19200 7034 20000 7064
rect 18137 7032 20000 7034
rect 18137 6976 18142 7032
rect 18198 6976 20000 7032
rect 18137 6974 20000 6976
rect 18137 6971 18203 6974
rect 19200 6944 20000 6974
rect 0 6898 800 6928
rect 1761 6898 1827 6901
rect 4061 6898 4127 6901
rect 8385 6898 8451 6901
rect 0 6896 1827 6898
rect 0 6840 1766 6896
rect 1822 6840 1827 6896
rect 0 6838 1827 6840
rect 0 6808 800 6838
rect 1761 6835 1827 6838
rect 3144 6896 8451 6898
rect 3144 6840 4066 6896
rect 4122 6840 8390 6896
rect 8446 6840 8451 6896
rect 3144 6838 8451 6840
rect 3144 6765 3204 6838
rect 4061 6835 4127 6838
rect 8385 6835 8451 6838
rect 13813 6898 13879 6901
rect 14825 6898 14891 6901
rect 13813 6896 14891 6898
rect 13813 6840 13818 6896
rect 13874 6840 14830 6896
rect 14886 6840 14891 6896
rect 13813 6838 14891 6840
rect 13813 6835 13879 6838
rect 14825 6835 14891 6838
rect 3141 6760 3207 6765
rect 3141 6704 3146 6760
rect 3202 6704 3207 6760
rect 3141 6699 3207 6704
rect 18505 6626 18571 6629
rect 19200 6626 20000 6656
rect 18505 6624 20000 6626
rect 18505 6568 18510 6624
rect 18566 6568 20000 6624
rect 18505 6566 20000 6568
rect 18505 6563 18571 6566
rect 3909 6560 4229 6561
rect 0 6490 800 6520
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 19200 6536 20000 6566
rect 15770 6495 16090 6496
rect 1485 6490 1551 6493
rect 0 6488 1551 6490
rect 0 6432 1490 6488
rect 1546 6432 1551 6488
rect 0 6430 1551 6432
rect 0 6400 800 6430
rect 1485 6427 1551 6430
rect 12157 6354 12223 6357
rect 13813 6354 13879 6357
rect 12157 6352 13879 6354
rect 12157 6296 12162 6352
rect 12218 6296 13818 6352
rect 13874 6296 13879 6352
rect 12157 6294 13879 6296
rect 12157 6291 12223 6294
rect 13813 6291 13879 6294
rect 2129 6218 2195 6221
rect 4429 6218 4495 6221
rect 2129 6216 4495 6218
rect 2129 6160 2134 6216
rect 2190 6160 4434 6216
rect 4490 6160 4495 6216
rect 2129 6158 4495 6160
rect 2129 6155 2195 6158
rect 4429 6155 4495 6158
rect 11053 6218 11119 6221
rect 14365 6218 14431 6221
rect 11053 6216 14431 6218
rect 11053 6160 11058 6216
rect 11114 6160 14370 6216
rect 14426 6160 14431 6216
rect 11053 6158 14431 6160
rect 11053 6155 11119 6158
rect 14365 6155 14431 6158
rect 18505 6218 18571 6221
rect 19200 6218 20000 6248
rect 18505 6216 20000 6218
rect 18505 6160 18510 6216
rect 18566 6160 20000 6216
rect 18505 6158 20000 6160
rect 18505 6155 18571 6158
rect 19200 6128 20000 6158
rect 0 6082 800 6112
rect 1853 6082 1919 6085
rect 0 6080 1919 6082
rect 0 6024 1858 6080
rect 1914 6024 1919 6080
rect 0 6022 1919 6024
rect 0 5992 800 6022
rect 1853 6019 1919 6022
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 11145 5946 11211 5949
rect 11513 5946 11579 5949
rect 11145 5944 11579 5946
rect 11145 5888 11150 5944
rect 11206 5888 11518 5944
rect 11574 5888 11579 5944
rect 11145 5886 11579 5888
rect 11145 5883 11211 5886
rect 11513 5883 11579 5886
rect 4153 5810 4219 5813
rect 8109 5810 8175 5813
rect 4153 5808 8175 5810
rect 4153 5752 4158 5808
rect 4214 5752 8114 5808
rect 8170 5752 8175 5808
rect 4153 5750 8175 5752
rect 4153 5747 4219 5750
rect 8109 5747 8175 5750
rect 12341 5810 12407 5813
rect 13813 5810 13879 5813
rect 15469 5810 15535 5813
rect 12341 5808 15535 5810
rect 12341 5752 12346 5808
rect 12402 5752 13818 5808
rect 13874 5752 15474 5808
rect 15530 5752 15535 5808
rect 12341 5750 15535 5752
rect 12341 5747 12407 5750
rect 13813 5747 13879 5750
rect 15469 5747 15535 5750
rect 3233 5674 3299 5677
rect 8477 5674 8543 5677
rect 3233 5672 8543 5674
rect 3233 5616 3238 5672
rect 3294 5616 8482 5672
rect 8538 5616 8543 5672
rect 3233 5614 8543 5616
rect 3233 5611 3299 5614
rect 8477 5611 8543 5614
rect 18505 5674 18571 5677
rect 19200 5674 20000 5704
rect 18505 5672 20000 5674
rect 18505 5616 18510 5672
rect 18566 5616 20000 5672
rect 18505 5614 20000 5616
rect 18505 5611 18571 5614
rect 19200 5584 20000 5614
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 4797 5266 4863 5269
rect 8385 5266 8451 5269
rect 9305 5266 9371 5269
rect 4797 5264 9371 5266
rect 4797 5208 4802 5264
rect 4858 5208 8390 5264
rect 8446 5208 9310 5264
rect 9366 5208 9371 5264
rect 4797 5206 9371 5208
rect 4797 5203 4863 5206
rect 8385 5203 8451 5206
rect 9305 5203 9371 5206
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 1853 5130 1919 5133
rect 0 5128 1919 5130
rect 0 5072 1858 5128
rect 1914 5072 1919 5128
rect 0 5070 1919 5072
rect 0 5040 800 5070
rect 1853 5067 1919 5070
rect 10777 5130 10843 5133
rect 13445 5130 13511 5133
rect 15193 5130 15259 5133
rect 10777 5128 13370 5130
rect 10777 5072 10782 5128
rect 10838 5072 13370 5128
rect 10777 5070 13370 5072
rect 10777 5067 10843 5070
rect 13310 4994 13370 5070
rect 13445 5128 15259 5130
rect 13445 5072 13450 5128
rect 13506 5072 15198 5128
rect 15254 5072 15259 5128
rect 13445 5070 15259 5072
rect 13445 5067 13511 5070
rect 15193 5067 15259 5070
rect 15193 4994 15259 4997
rect 13310 4992 15259 4994
rect 13310 4936 15198 4992
rect 15254 4936 15259 4992
rect 13310 4934 15259 4936
rect 15193 4931 15259 4934
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 12249 4860 12315 4861
rect 12198 4796 12204 4860
rect 12268 4858 12315 4860
rect 18137 4858 18203 4861
rect 19200 4858 20000 4888
rect 12268 4856 12360 4858
rect 12310 4800 12360 4856
rect 12268 4798 12360 4800
rect 18137 4856 20000 4858
rect 18137 4800 18142 4856
rect 18198 4800 20000 4856
rect 18137 4798 20000 4800
rect 12268 4796 12315 4798
rect 12249 4795 12315 4796
rect 18137 4795 18203 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 1393 4722 1459 4725
rect 0 4720 1459 4722
rect 0 4664 1398 4720
rect 1454 4664 1459 4720
rect 0 4662 1459 4664
rect 0 4632 800 4662
rect 1393 4659 1459 4662
rect 3877 4722 3943 4725
rect 5165 4722 5231 4725
rect 3877 4720 5231 4722
rect 3877 4664 3882 4720
rect 3938 4664 5170 4720
rect 5226 4664 5231 4720
rect 3877 4662 5231 4664
rect 3877 4659 3943 4662
rect 5165 4659 5231 4662
rect 10961 4722 11027 4725
rect 14089 4722 14155 4725
rect 10961 4720 14155 4722
rect 10961 4664 10966 4720
rect 11022 4664 14094 4720
rect 14150 4664 14155 4720
rect 10961 4662 14155 4664
rect 10961 4659 11027 4662
rect 14089 4659 14155 4662
rect 2681 4586 2747 4589
rect 4613 4586 4679 4589
rect 2681 4584 4679 4586
rect 2681 4528 2686 4584
rect 2742 4528 4618 4584
rect 4674 4528 4679 4584
rect 2681 4526 4679 4528
rect 2681 4523 2747 4526
rect 4613 4523 4679 4526
rect 4981 4586 5047 4589
rect 5533 4586 5599 4589
rect 8477 4586 8543 4589
rect 4981 4584 8543 4586
rect 4981 4528 4986 4584
rect 5042 4528 5538 4584
rect 5594 4528 8482 4584
rect 8538 4528 8543 4584
rect 4981 4526 8543 4528
rect 4981 4523 5047 4526
rect 5533 4523 5599 4526
rect 8477 4523 8543 4526
rect 11462 4388 11468 4452
rect 11532 4450 11538 4452
rect 11605 4450 11671 4453
rect 11532 4448 11671 4450
rect 11532 4392 11610 4448
rect 11666 4392 11671 4448
rect 11532 4390 11671 4392
rect 11532 4388 11538 4390
rect 11605 4387 11671 4390
rect 18505 4450 18571 4453
rect 19200 4450 20000 4480
rect 18505 4448 20000 4450
rect 18505 4392 18510 4448
rect 18566 4392 20000 4448
rect 18505 4390 20000 4392
rect 18505 4387 18571 4390
rect 3909 4384 4229 4385
rect 0 4314 800 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19200 4360 20000 4390
rect 15770 4319 16090 4320
rect 3325 4314 3391 4317
rect 0 4312 3391 4314
rect 0 4256 3330 4312
rect 3386 4256 3391 4312
rect 0 4254 3391 4256
rect 0 4224 800 4254
rect 3325 4251 3391 4254
rect 10685 4178 10751 4181
rect 16389 4178 16455 4181
rect 10685 4176 16455 4178
rect 10685 4120 10690 4176
rect 10746 4120 16394 4176
rect 16450 4120 16455 4176
rect 10685 4118 16455 4120
rect 10685 4115 10751 4118
rect 16389 4115 16455 4118
rect 5533 4042 5599 4045
rect 10961 4042 11027 4045
rect 13905 4042 13971 4045
rect 5533 4040 11027 4042
rect 5533 3984 5538 4040
rect 5594 3984 10966 4040
rect 11022 3984 11027 4040
rect 5533 3982 11027 3984
rect 5533 3979 5599 3982
rect 10961 3979 11027 3982
rect 12390 4040 13971 4042
rect 12390 3984 13910 4040
rect 13966 3984 13971 4040
rect 12390 3982 13971 3984
rect 0 3906 800 3936
rect 2865 3906 2931 3909
rect 0 3904 2931 3906
rect 0 3848 2870 3904
rect 2926 3848 2931 3904
rect 0 3846 2931 3848
rect 0 3816 800 3846
rect 2865 3843 2931 3846
rect 3550 3844 3556 3908
rect 3620 3906 3626 3908
rect 3693 3906 3759 3909
rect 3620 3904 3759 3906
rect 3620 3848 3698 3904
rect 3754 3848 3759 3904
rect 3620 3846 3759 3848
rect 3620 3844 3626 3846
rect 3693 3843 3759 3846
rect 4337 3906 4403 3909
rect 6085 3906 6151 3909
rect 12390 3906 12450 3982
rect 13905 3979 13971 3982
rect 18137 4042 18203 4045
rect 19200 4042 20000 4072
rect 18137 4040 20000 4042
rect 18137 3984 18142 4040
rect 18198 3984 20000 4040
rect 18137 3982 20000 3984
rect 18137 3979 18203 3982
rect 19200 3952 20000 3982
rect 4337 3904 6151 3906
rect 4337 3848 4342 3904
rect 4398 3848 6090 3904
rect 6146 3848 6151 3904
rect 4337 3846 6151 3848
rect 4337 3843 4403 3846
rect 6085 3843 6151 3846
rect 7422 3846 12450 3906
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 2589 3770 2655 3773
rect 6729 3770 6795 3773
rect 2589 3768 6795 3770
rect 2589 3712 2594 3768
rect 2650 3712 6734 3768
rect 6790 3712 6795 3768
rect 2589 3710 6795 3712
rect 2589 3707 2655 3710
rect 6729 3707 6795 3710
rect 5717 3634 5783 3637
rect 6177 3634 6243 3637
rect 7422 3634 7482 3846
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 9029 3770 9095 3773
rect 10869 3770 10935 3773
rect 9029 3768 10935 3770
rect 9029 3712 9034 3768
rect 9090 3712 10874 3768
rect 10930 3712 10935 3768
rect 9029 3710 10935 3712
rect 9029 3707 9095 3710
rect 10869 3707 10935 3710
rect 5717 3632 7482 3634
rect 5717 3576 5722 3632
rect 5778 3576 6182 3632
rect 6238 3576 7482 3632
rect 5717 3574 7482 3576
rect 9581 3634 9647 3637
rect 16481 3634 16547 3637
rect 9581 3632 16547 3634
rect 9581 3576 9586 3632
rect 9642 3576 16486 3632
rect 16542 3576 16547 3632
rect 9581 3574 16547 3576
rect 5717 3571 5783 3574
rect 6177 3571 6243 3574
rect 9581 3571 9647 3574
rect 16481 3571 16547 3574
rect 18505 3634 18571 3637
rect 19200 3634 20000 3664
rect 18505 3632 20000 3634
rect 18505 3576 18510 3632
rect 18566 3576 20000 3632
rect 18505 3574 20000 3576
rect 18505 3571 18571 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 2497 3498 2563 3501
rect 0 3496 2563 3498
rect 0 3440 2502 3496
rect 2558 3440 2563 3496
rect 0 3438 2563 3440
rect 0 3408 800 3438
rect 2497 3435 2563 3438
rect 4429 3498 4495 3501
rect 5349 3498 5415 3501
rect 4429 3496 5415 3498
rect 4429 3440 4434 3496
rect 4490 3440 5354 3496
rect 5410 3440 5415 3496
rect 4429 3438 5415 3440
rect 4429 3435 4495 3438
rect 5349 3435 5415 3438
rect 10501 3498 10567 3501
rect 13261 3498 13327 3501
rect 10501 3496 13327 3498
rect 10501 3440 10506 3496
rect 10562 3440 13266 3496
rect 13322 3440 13327 3496
rect 10501 3438 13327 3440
rect 10501 3435 10567 3438
rect 13261 3435 13327 3438
rect 11237 3362 11303 3365
rect 15561 3362 15627 3365
rect 11237 3360 15627 3362
rect 11237 3304 11242 3360
rect 11298 3304 15566 3360
rect 15622 3304 15627 3360
rect 11237 3302 15627 3304
rect 11237 3299 11303 3302
rect 15561 3299 15627 3302
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 1761 3226 1827 3229
rect 3693 3226 3759 3229
rect 1761 3224 3759 3226
rect 1761 3168 1766 3224
rect 1822 3168 3698 3224
rect 3754 3168 3759 3224
rect 1761 3166 3759 3168
rect 1761 3163 1827 3166
rect 3693 3163 3759 3166
rect 10869 3226 10935 3229
rect 18137 3226 18203 3229
rect 19200 3226 20000 3256
rect 10869 3224 12266 3226
rect 10869 3168 10874 3224
rect 10930 3168 12266 3224
rect 10869 3166 12266 3168
rect 10869 3163 10935 3166
rect 0 3090 800 3120
rect 2221 3090 2287 3093
rect 0 3088 2287 3090
rect 0 3032 2226 3088
rect 2282 3032 2287 3088
rect 0 3030 2287 3032
rect 0 3000 800 3030
rect 2221 3027 2287 3030
rect 5809 3090 5875 3093
rect 12065 3090 12131 3093
rect 5809 3088 12131 3090
rect 5809 3032 5814 3088
rect 5870 3032 12070 3088
rect 12126 3032 12131 3088
rect 5809 3030 12131 3032
rect 12206 3090 12266 3166
rect 18137 3224 20000 3226
rect 18137 3168 18142 3224
rect 18198 3168 20000 3224
rect 18137 3166 20000 3168
rect 18137 3163 18203 3166
rect 19200 3136 20000 3166
rect 14181 3090 14247 3093
rect 17033 3090 17099 3093
rect 12206 3088 17099 3090
rect 12206 3032 14186 3088
rect 14242 3032 17038 3088
rect 17094 3032 17099 3088
rect 12206 3030 17099 3032
rect 5809 3027 5875 3030
rect 12065 3027 12131 3030
rect 14181 3027 14247 3030
rect 17033 3027 17099 3030
rect 1577 2954 1643 2957
rect 16113 2954 16179 2957
rect 1577 2952 16179 2954
rect 1577 2896 1582 2952
rect 1638 2896 16118 2952
rect 16174 2896 16179 2952
rect 1577 2894 16179 2896
rect 1577 2891 1643 2894
rect 16113 2891 16179 2894
rect 2313 2818 2379 2821
rect 6729 2818 6795 2821
rect 2313 2816 6795 2818
rect 2313 2760 2318 2816
rect 2374 2760 6734 2816
rect 6790 2760 6795 2816
rect 2313 2758 6795 2760
rect 2313 2755 2379 2758
rect 6729 2755 6795 2758
rect 6874 2752 7194 2753
rect 0 2682 800 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 2773 2682 2839 2685
rect 0 2680 2839 2682
rect 0 2624 2778 2680
rect 2834 2624 2839 2680
rect 0 2622 2839 2624
rect 0 2592 800 2622
rect 2773 2619 2839 2622
rect 10409 2682 10475 2685
rect 11462 2682 11468 2684
rect 10409 2680 11468 2682
rect 10409 2624 10414 2680
rect 10470 2624 11468 2680
rect 10409 2622 11468 2624
rect 10409 2619 10475 2622
rect 11462 2620 11468 2622
rect 11532 2620 11538 2684
rect 17769 2682 17835 2685
rect 19200 2682 20000 2712
rect 17769 2680 20000 2682
rect 17769 2624 17774 2680
rect 17830 2624 20000 2680
rect 17769 2622 20000 2624
rect 17769 2619 17835 2622
rect 19200 2592 20000 2622
rect 0 2274 800 2304
rect 1485 2274 1551 2277
rect 0 2272 1551 2274
rect 0 2216 1490 2272
rect 1546 2216 1551 2272
rect 0 2214 1551 2216
rect 0 2184 800 2214
rect 1485 2211 1551 2214
rect 17861 2274 17927 2277
rect 19200 2274 20000 2304
rect 17861 2272 20000 2274
rect 17861 2216 17866 2272
rect 17922 2216 20000 2272
rect 17861 2214 20000 2216
rect 17861 2211 17927 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19200 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 800 1896
rect 1853 1866 1919 1869
rect 0 1864 1919 1866
rect 0 1808 1858 1864
rect 1914 1808 1919 1864
rect 0 1806 1919 1808
rect 0 1776 800 1806
rect 1853 1803 1919 1806
rect 17585 1866 17651 1869
rect 19200 1866 20000 1896
rect 17585 1864 20000 1866
rect 17585 1808 17590 1864
rect 17646 1808 20000 1864
rect 17585 1806 20000 1808
rect 17585 1803 17651 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 2221 1458 2287 1461
rect 0 1456 2287 1458
rect 0 1400 2226 1456
rect 2282 1400 2287 1456
rect 0 1398 2287 1400
rect 0 1368 800 1398
rect 2221 1395 2287 1398
rect 17677 1458 17743 1461
rect 19200 1458 20000 1488
rect 17677 1456 20000 1458
rect 17677 1400 17682 1456
rect 17738 1400 20000 1456
rect 17677 1398 20000 1400
rect 17677 1395 17743 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 1393 1050 1459 1053
rect 0 1048 1459 1050
rect 0 992 1398 1048
rect 1454 992 1459 1048
rect 0 990 1459 992
rect 0 960 800 990
rect 1393 987 1459 990
rect 16573 1050 16639 1053
rect 19200 1050 20000 1080
rect 16573 1048 20000 1050
rect 16573 992 16578 1048
rect 16634 992 20000 1048
rect 16573 990 20000 992
rect 16573 987 16639 990
rect 19200 960 20000 990
rect 0 642 800 672
rect 1761 642 1827 645
rect 0 640 1827 642
rect 0 584 1766 640
rect 1822 584 1827 640
rect 0 582 1827 584
rect 0 552 800 582
rect 1761 579 1827 582
rect 17493 642 17559 645
rect 19200 642 20000 672
rect 17493 640 20000 642
rect 17493 584 17498 640
rect 17554 584 20000 640
rect 17493 582 20000 584
rect 17493 579 17559 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 3325 234 3391 237
rect 0 232 3391 234
rect 0 176 3330 232
rect 3386 176 3391 232
rect 0 174 3391 176
rect 0 144 800 174
rect 3325 171 3391 174
rect 17769 234 17835 237
rect 19200 234 20000 264
rect 17769 232 20000 234
rect 17769 176 17774 232
rect 17830 176 20000 232
rect 17769 174 20000 176
rect 17769 171 17835 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 12204 9420 12268 9484
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3556 7712 3620 7716
rect 3556 7656 3570 7712
rect 3570 7656 3620 7712
rect 3556 7652 3620 7656
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 12204 4856 12268 4860
rect 12204 4800 12254 4856
rect 12254 4800 12268 4856
rect 12204 4796 12268 4800
rect 11468 4388 11532 4452
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 3556 3844 3620 3908
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 11468 2620 11532 2684
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3555 7716 3621 7717
rect 3555 7652 3556 7716
rect 3620 7652 3621 7716
rect 3555 7651 3621 7652
rect 3558 3909 3618 7651
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3555 3908 3621 3909
rect 3555 3844 3556 3908
rect 3620 3844 3621 3908
rect 3555 3843 3621 3844
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12203 9484 12269 9485
rect 12203 9420 12204 9484
rect 12268 9420 12269 9484
rect 12203 9419 12269 9420
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 12206 4861 12266 9419
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12203 4860 12269 4861
rect 12203 4796 12204 4860
rect 12268 4796 12269 4860
rect 12203 4795 12269 4796
rect 11467 4452 11533 4453
rect 11467 4388 11468 4452
rect 11532 4388 11533 4452
rect 11467 4387 11533 4388
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 11470 2685 11530 4387
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 11467 2684 11533 2685
rect 11467 2620 11468 2684
rect 11532 2620 11533 2684
rect 11467 2619 11533 2620
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 2128 13125 2688
rect 15770 14176 16091 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16091 14176
rect 15770 13088 16091 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16091 13088
rect 15770 12000 16091 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16091 12000
rect 15770 10912 16091 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16091 10912
rect 15770 9824 16091 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16091 9824
rect 15770 8736 16091 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16091 8736
rect 15770 7648 16091 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16091 7648
rect 15770 6560 16091 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16091 6560
rect 15770 5472 16091 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16091 5472
rect 15770 4384 16091 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16091 4384
rect 15770 3296 16091 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16091 3296
rect 15770 2208 16091 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16091 2208
rect 15770 2128 16091 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform -1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output49
timestamp 1624635492
transform -1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1624635492
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform -1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform -1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3956 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 3956 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4784 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4692 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1624635492
transform -1 0 4692 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1624635492
transform -1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1624635492
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1624635492
transform -1 0 6348 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1624635492
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1624635492
transform 1 0 5612 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1624635492
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform -1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6532 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 8280 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 8556 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform -1 0 8372 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform -1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform -1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 9016 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1624635492
transform -1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_95
timestamp 1624635492
transform 1 0 9844 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1624635492
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9844 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10120 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1624635492
transform -1 0 11500 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11776 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1624635492
transform -1 0 12512 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output50
timestamp 1624635492
transform -1 0 11316 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output52
timestamp 1624635492
transform -1 0 12880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1624635492
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform -1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output51
timestamp 1624635492
transform -1 0 13064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 13432 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 12880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1624635492
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform -1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_143 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14260 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1624635492
transform -1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1624635492
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 15180 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1624635492
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1624635492
transform 1 0 15732 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1624635492
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform 1 0 16284 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1624635492
transform -1 0 16284 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _36_
timestamp 1624635492
transform -1 0 16376 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 16560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_168
timestamp 1624635492
transform 1 0 16560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1624635492
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform -1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1624635492
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1624635492
transform -1 0 17480 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1624635492
transform -1 0 17480 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform 1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform 1 0 18216 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output47
timestamp 1624635492
transform 1 0 18216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform -1 0 3220 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1624635492
transform 1 0 4692 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1624635492
transform -1 0 4692 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform -1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1624635492
transform 1 0 4968 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 5244 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 6716 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7452 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11316 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform -1 0 10304 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1624635492
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12052 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1624635492
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1624635492
transform -1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 13892 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1624635492
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1624635492
transform -1 0 16560 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1624635492
transform 1 0 16192 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1624635492
transform -1 0 17480 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1624635492
transform -1 0 17848 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1624635492
transform -1 0 17204 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1624635492
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1624635492
transform -1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_178
timestamp 1624635492
transform 1 0 17480 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1624635492
transform -1 0 2024 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2024 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3496 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1624635492
transform -1 0 5980 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_56
timestamp 1624635492
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7728 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 7544 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9200 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1624635492
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1624635492
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1624635492
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_110
timestamp 1624635492
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14444 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14444 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_133
timestamp 1624635492
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_158 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15640 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_166
timestamp 1624635492
transform 1 0 16376 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1624635492
transform -1 0 17848 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1624635492
transform -1 0 17572 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1624635492
transform -1 0 17296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1624635492
transform 1 0 17848 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1624635492
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1624635492
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1624635492
transform -1 0 6164 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6624 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 6440 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1624635492
transform -1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11224 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9568 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 9292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1624635492
transform -1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 9568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1624635492
transform 1 0 12236 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1624635492
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 15180 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_155
timestamp 1624635492
transform 1 0 15364 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1624635492
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_167
timestamp 1624635492
transform 1 0 16468 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_175
timestamp 1624635492
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_179
timestamp 1624635492
transform 1 0 17572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1624635492
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 2852 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3956 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3128 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1624635492
transform 1 0 5612 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 6532 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  output110
timestamp 1624635492
transform -1 0 6164 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 7360 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1624635492
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 8188 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9292 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1624635492
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1624635492
transform -1 0 10304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_100
timestamp 1624635492
transform 1 0 10304 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 13156 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 15548 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13248 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_131
timestamp 1624635492
transform 1 0 13156 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1624635492
transform 1 0 15548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_162
timestamp 1624635492
transform 1 0 16008 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform -1 0 18124 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1624635492
transform 1 0 17664 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_170
timestamp 1624635492
transform 1 0 16744 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_172
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1624635492
transform 1 0 18124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 2116 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2944 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1624635492
transform 1 0 2668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1624635492
transform -1 0 2668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1624635492
transform -1 0 2392 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 1564 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1624635492
transform -1 0 3312 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1624635492
transform 1 0 3312 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1624635492
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5520 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4692 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6992 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1624635492
transform -1 0 6348 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1624635492
transform -1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8648 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1624635492
transform 1 0 7912 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 9016 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_82
timestamp 1624635492
transform 1 0 8648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9016 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9936 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1624635492
transform -1 0 9936 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 10488 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12144 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1624635492
transform 1 0 11960 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11592 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 15088 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1624635492
transform 1 0 12788 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1624635492
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_140
timestamp 1624635492
transform 1 0 13984 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1624635492
transform 1 0 15180 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_164
timestamp 1624635492
transform 1 0 16192 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1624635492
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_172
timestamp 1624635492
transform 1 0 16928 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1624635492
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1624635492
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1624635492
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1624635492
transform -1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1624635492
transform -1 0 17848 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1624635492
transform -1 0 17848 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_185
timestamp 1624635492
transform 1 0 18124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_185
timestamp 1624635492
transform 1 0 18124 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1624635492
transform -1 0 18124 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1624635492
transform -1 0 18124 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2300 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 2116 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4692 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1624635492
transform 1 0 6440 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_48
timestamp 1624635492
transform 1 0 5520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7452 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11408 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9936 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1624635492
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13432 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1624635492
transform -1 0 12604 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13432 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1624635492
transform -1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_162
timestamp 1624635492
transform 1 0 16008 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1624635492
transform -1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1624635492
transform -1 0 17388 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1624635492
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_174
timestamp 1624635492
transform 1 0 17112 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp 1624635492
transform 1 0 17388 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 1564 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1624635492
transform 1 0 4416 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 6348 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 8556 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7268 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 8372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 10120 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp 1624635492
transform 1 0 10028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1624635492
transform 1 0 12328 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1624635492
transform 1 0 12052 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13156 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1624635492
transform 1 0 14536 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1624635492
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_168
timestamp 1624635492
transform 1 0 16560 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1624635492
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_172
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1624635492
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1624635492
transform -1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1624635492
transform -1 0 17848 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1624635492
transform 1 0 18124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1624635492
transform -1 0 18124 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2576 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2576 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform -1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4876 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 3772 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1624635492
transform 1 0 6348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 6808 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1624635492
transform -1 0 7912 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1624635492
transform -1 0 8740 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1624635492
transform 1 0 8740 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1624635492
transform -1 0 10764 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1624635492
transform 1 0 10856 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_105
timestamp 1624635492
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1624635492
transform -1 0 13156 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 15824 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_127
timestamp 1624635492
transform 1 0 12788 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_133
timestamp 1624635492
transform 1 0 13340 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 15824 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1624635492
transform -1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 18584 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform 1 0 17664 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_176
timestamp 1624635492
transform 1 0 17296 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 2852 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1624635492
transform 1 0 3220 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 4324 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4324 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1624635492
transform 1 0 5152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1624635492
transform -1 0 6348 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_47
timestamp 1624635492
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1624635492
transform -1 0 8188 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9660 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 9660 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1624635492
transform 1 0 11776 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1624635492
transform -1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1624635492
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14260 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1624635492
transform 1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1624635492
transform 1 0 15088 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 15916 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1624635492
transform -1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1624635492
transform -1 0 17388 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1624635492
transform -1 0 18584 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform 1 0 17664 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1624635492
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1624635492
transform 1 0 1932 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2208 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1624635492
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6808 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1624635492
transform -1 0 6440 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_48
timestamp 1624635492
transform 1 0 5520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1624635492
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9568 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10396 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1624635492
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1624635492
transform 1 0 12144 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1624635492
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1624635492
transform 1 0 11224 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1624635492
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14444 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_138
timestamp 1624635492
transform 1 0 13800 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 16008 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_156
timestamp 1624635492
transform 1 0 15456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1624635492
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1624635492
transform 1 0 18308 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1624635492
transform 1 0 17480 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2668 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1624635492
transform -1 0 3220 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1624635492
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1624635492
transform 1 0 2852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1624635492
transform 1 0 3772 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1624635492
transform 1 0 4048 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 5336 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1624635492
transform 1 0 3220 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 4140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 5336 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp 1624635492
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7452 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1624635492
transform -1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7636 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1624635492
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1624635492
transform 1 0 8464 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11040 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10948 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_91
timestamp 1624635492
transform 1 0 9476 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1624635492
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10948 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1624635492
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 12144 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11776 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12328 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 13156 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13156 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_140
timestamp 1624635492
transform 1 0 13984 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1624635492
transform 1 0 14444 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14168 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1624635492
transform 1 0 17388 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 18584 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1624635492
transform -1 0 17388 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_172
timestamp 1624635492
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform -1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5612 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3312 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1624635492
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1624635492
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 7912 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9384 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 13156 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13340 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1624635492
transform -1 0 16836 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 18584 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3772 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform -1 0 2300 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5980 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1624635492
transform -1 0 7636 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1624635492
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1624635492
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_50
timestamp 1624635492
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1624635492
transform -1 0 8464 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1624635492
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 11960 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11960 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1624635492
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1624635492
transform 1 0 13432 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15364 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 15180 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 15364 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1624635492
transform 1 0 14628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1624635492
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform -1 0 17572 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 17204 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1624635492
transform 1 0 2576 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1624635492
transform -1 0 1932 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1624635492
transform 1 0 1932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 3036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_15
timestamp 1624635492
transform 1 0 2484 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 4692 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1624635492
transform 1 0 3588 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 7452 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9844 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1624635492
transform 1 0 8924 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_94
timestamp 1624635492
transform 1 0 9752 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1624635492
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 12236 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1624635492
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1624635492
transform 1 0 14352 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1624635492
transform -1 0 16836 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16008 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1624635492
transform 1 0 17756 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2116 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1624635492
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 4692 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6072 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1624635492
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1624635492
transform 1 0 8188 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1624635492
transform -1 0 8188 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1624635492
transform 1 0 7084 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1624635492
transform -1 0 9384 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10396 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9568 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11868 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 14260 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1624635492
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1624635492
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 16284 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 17940 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 18584 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 1624635492
transform 1 0 17940 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1624635492
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1624635492
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 2484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1624635492
transform -1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1624635492
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1624635492
transform 1 0 2852 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 2944 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_26
timestamp 1624635492
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1624635492
transform 1 0 3036 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1624635492
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 1624635492
transform 1 0 4692 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_36
timestamp 1624635492
transform 1 0 4416 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 4324 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_51
timestamp 1624635492
transform 1 0 5796 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_47
timestamp 1624635492
transform 1 0 5428 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_44
timestamp 1624635492
transform 1 0 5152 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 5428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1624635492
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_54
timestamp 1624635492
transform 1 0 6072 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 6624 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8096 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9936 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1624635492
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1624635492
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7360 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_74
timestamp 1624635492
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1624635492
transform -1 0 11500 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9476 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_96
timestamp 1624635492
transform 1 0 9936 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_89
timestamp 1624635492
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_100
timestamp 1624635492
transform 1 0 10304 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1624635492
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_118
timestamp 1624635492
transform 1 0 11960 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_112
timestamp 1624635492
transform 1 0 11408 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_115
timestamp 1624635492
transform 1 0 11684 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1624635492
transform -1 0 14720 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1624635492
transform -1 0 15180 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 13708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1624635492
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1624635492
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 15180 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 15548 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1624635492
transform 1 0 14720 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp 1624635492
transform 1 0 16192 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp 1624635492
transform 1 0 15548 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 15732 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 15916 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15824 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 16192 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _35_
timestamp 1624635492
transform -1 0 16560 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16560 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17204 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1624635492
transform 1 0 17388 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 18216 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1624635492
transform -1 0 17848 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform -1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1624635492
transform -1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1624635492
transform -1 0 18584 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform -1 0 2392 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1624635492
transform 1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_28
timestamp 1624635492
transform 1 0 3680 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_40
timestamp 1624635492
transform 1 0 4784 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1624635492
transform 1 0 5888 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1624635492
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1624635492
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1624635492
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1624635492
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1624635492
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_123
timestamp 1624635492
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 12696 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_21_133
timestamp 1624635492
transform 1 0 13340 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_145
timestamp 1624635492
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15640 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_149
timestamp 1624635492
transform 1 0 14812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1624635492
transform -1 0 18584 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1624635492
transform -1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1624635492
transform -1 0 17848 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1624635492
transform -1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1624635492
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1624635492
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1624635492
transform -1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1624635492
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 4324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_35
timestamp 1624635492
transform 1 0 4324 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 6440 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output48
timestamp 1624635492
transform -1 0 5888 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_47
timestamp 1624635492
transform 1 0 5428 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_52
timestamp 1624635492
transform 1 0 5888 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_59
timestamp 1624635492
transform 1 0 6532 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1624635492
transform 1 0 7728 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_71
timestamp 1624635492
transform 1 0 7636 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_77
timestamp 1624635492
transform 1 0 8188 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform -1 0 10304 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1624635492
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_88
timestamp 1624635492
transform 1 0 9200 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_100
timestamp 1624635492
transform 1 0 10304 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11776 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform -1 0 12512 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1624635492
transform 1 0 11408 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 1624635492
transform 1 0 11868 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_124
timestamp 1624635492
transform 1 0 12512 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_136
timestamp 1624635492
transform 1 0 13616 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15824 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1624635492
transform -1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform -1 0 14904 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform 1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 15180 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_150
timestamp 1624635492
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _34_
timestamp 1624635492
transform 1 0 17204 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 17112 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform -1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1624635492
transform -1 0 18216 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 17848 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1624635492
transform -1 0 17112 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1624635492
transform 1 0 16652 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 1122 16400 1178 17200 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 3330 16400 3386 17200 6 SC_IN_TOP
port 2 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 SC_OUT_BOT
port 3 nsew signal tristate
rlabel metal2 s 5538 16400 5594 17200 6 SC_OUT_TOP
port 4 nsew signal tristate
rlabel metal2 s 1214 0 1270 800 6 bottom_grid_pin_0_
port 5 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_10_
port 6 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 bottom_grid_pin_11_
port 7 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 bottom_grid_pin_12_
port 8 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 bottom_grid_pin_13_
port 9 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 bottom_grid_pin_14_
port 10 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 bottom_grid_pin_15_
port 11 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_1_
port 12 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 bottom_grid_pin_2_
port 13 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 bottom_grid_pin_3_
port 14 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 bottom_grid_pin_4_
port 15 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 bottom_grid_pin_5_
port 16 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 bottom_grid_pin_6_
port 17 nsew signal tristate
rlabel metal2 s 7562 0 7618 800 6 bottom_grid_pin_7_
port 18 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 bottom_grid_pin_8_
port 19 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 bottom_grid_pin_9_
port 20 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 bottom_width_0_height_0__pin_0_
port 21 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 bottom_width_0_height_0__pin_1_lower
port 22 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 bottom_width_0_height_0__pin_1_upper
port 23 nsew signal tristate
rlabel metal2 s 7746 16400 7802 17200 6 ccff_head
port 24 nsew signal input
rlabel metal2 s 9954 16400 10010 17200 6 ccff_tail
port 25 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[0]
port 26 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[10]
port 27 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_in[11]
port 28 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 chanx_left_in[12]
port 29 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 chanx_left_in[13]
port 30 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 chanx_left_in[14]
port 31 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 chanx_left_in[15]
port 32 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 chanx_left_in[16]
port 33 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 chanx_left_in[17]
port 34 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 chanx_left_in[18]
port 35 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 chanx_left_in[19]
port 36 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[1]
port 37 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[2]
port 38 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[3]
port 39 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[4]
port 40 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[5]
port 41 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[6]
port 42 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[7]
port 43 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[8]
port 44 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[9]
port 45 nsew signal input
rlabel metal3 s 0 552 800 672 6 chanx_left_out[0]
port 46 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[10]
port 47 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[11]
port 48 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[12]
port 49 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[13]
port 50 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[14]
port 51 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 chanx_left_out[15]
port 52 nsew signal tristate
rlabel metal3 s 0 7216 800 7336 6 chanx_left_out[16]
port 53 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 chanx_left_out[17]
port 54 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 chanx_left_out[18]
port 55 nsew signal tristate
rlabel metal3 s 0 8440 800 8560 6 chanx_left_out[19]
port 56 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 chanx_left_out[1]
port 57 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[2]
port 58 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[3]
port 59 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 chanx_left_out[4]
port 60 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 chanx_left_out[5]
port 61 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[6]
port 62 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[7]
port 63 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_out[8]
port 64 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 chanx_left_out[9]
port 65 nsew signal tristate
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_in[0]
port 66 nsew signal input
rlabel metal3 s 19200 12928 20000 13048 6 chanx_right_in[10]
port 67 nsew signal input
rlabel metal3 s 19200 13336 20000 13456 6 chanx_right_in[11]
port 68 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[12]
port 69 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[13]
port 70 nsew signal input
rlabel metal3 s 19200 14696 20000 14816 6 chanx_right_in[14]
port 71 nsew signal input
rlabel metal3 s 19200 15104 20000 15224 6 chanx_right_in[15]
port 72 nsew signal input
rlabel metal3 s 19200 15512 20000 15632 6 chanx_right_in[16]
port 73 nsew signal input
rlabel metal3 s 19200 15920 20000 16040 6 chanx_right_in[17]
port 74 nsew signal input
rlabel metal3 s 19200 16328 20000 16448 6 chanx_right_in[18]
port 75 nsew signal input
rlabel metal3 s 19200 16736 20000 16856 6 chanx_right_in[19]
port 76 nsew signal input
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_in[1]
port 77 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[2]
port 78 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[3]
port 79 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 80 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[5]
port 81 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[6]
port 82 nsew signal input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[7]
port 83 nsew signal input
rlabel metal3 s 19200 12112 20000 12232 6 chanx_right_in[8]
port 84 nsew signal input
rlabel metal3 s 19200 12520 20000 12640 6 chanx_right_in[9]
port 85 nsew signal input
rlabel metal3 s 19200 144 20000 264 6 chanx_right_out[0]
port 86 nsew signal tristate
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[10]
port 87 nsew signal tristate
rlabel metal3 s 19200 4768 20000 4888 6 chanx_right_out[11]
port 88 nsew signal tristate
rlabel metal3 s 19200 5176 20000 5296 6 chanx_right_out[12]
port 89 nsew signal tristate
rlabel metal3 s 19200 5584 20000 5704 6 chanx_right_out[13]
port 90 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[14]
port 91 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[15]
port 92 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[16]
port 93 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[17]
port 94 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[18]
port 95 nsew signal tristate
rlabel metal3 s 19200 8168 20000 8288 6 chanx_right_out[19]
port 96 nsew signal tristate
rlabel metal3 s 19200 552 20000 672 6 chanx_right_out[1]
port 97 nsew signal tristate
rlabel metal3 s 19200 960 20000 1080 6 chanx_right_out[2]
port 98 nsew signal tristate
rlabel metal3 s 19200 1368 20000 1488 6 chanx_right_out[3]
port 99 nsew signal tristate
rlabel metal3 s 19200 1776 20000 1896 6 chanx_right_out[4]
port 100 nsew signal tristate
rlabel metal3 s 19200 2184 20000 2304 6 chanx_right_out[5]
port 101 nsew signal tristate
rlabel metal3 s 19200 2592 20000 2712 6 chanx_right_out[6]
port 102 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[7]
port 103 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[8]
port 104 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[9]
port 105 nsew signal tristate
rlabel metal2 s 14370 16400 14426 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 106 nsew signal tristate
rlabel metal2 s 16578 16400 16634 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 107 nsew signal input
rlabel metal2 s 18786 16400 18842 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 108 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 prog_clk_0_S_in
port 109 nsew signal input
rlabel metal3 s 0 144 800 264 6 prog_clk_0_W_out
port 110 nsew signal tristate
rlabel metal2 s 12162 16400 12218 17200 6 top_grid_pin_0_
port 111 nsew signal tristate
rlabel metal4 s 15771 2128 16091 14736 6 VPWR
port 112 nsew power bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VPWR
port 113 nsew power bidirectional
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 114 nsew power bidirectional
rlabel metal4 s 12805 2128 13125 14736 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
