magic
tech sky130A
magscale 1 2
timestamp 1656973540
<< viali >>
rect 5365 22185 5399 22219
rect 13369 22185 13403 22219
rect 20913 22185 20947 22219
rect 22017 22185 22051 22219
rect 10793 22117 10827 22151
rect 19257 22117 19291 22151
rect 20821 22117 20855 22151
rect 1593 22049 1627 22083
rect 7297 22049 7331 22083
rect 8585 22049 8619 22083
rect 9505 22049 9539 22083
rect 10241 22049 10275 22083
rect 12081 22049 12115 22083
rect 12173 22049 12207 22083
rect 13553 22049 13587 22083
rect 14197 22049 14231 22083
rect 16313 22049 16347 22083
rect 16773 22049 16807 22083
rect 17601 22049 17635 22083
rect 18521 22049 18555 22083
rect 19809 22049 19843 22083
rect 20177 22049 20211 22083
rect 21465 22049 21499 22083
rect 1961 21981 1995 22015
rect 2237 21981 2271 22015
rect 2605 21981 2639 22015
rect 2881 21981 2915 22015
rect 3249 21981 3283 22015
rect 3617 21981 3651 22015
rect 4070 21981 4104 22015
rect 4261 21981 4295 22015
rect 4629 21981 4663 22015
rect 4905 21981 4939 22015
rect 5457 21981 5491 22015
rect 5733 21981 5767 22015
rect 6185 21981 6219 22015
rect 6745 21981 6779 22015
rect 9229 21981 9263 22015
rect 10885 21981 10919 22015
rect 11161 21981 11195 22015
rect 12909 21981 12943 22015
rect 13185 21981 13219 22015
rect 13645 21981 13679 22015
rect 14933 21981 14967 22015
rect 15301 21981 15335 22015
rect 15485 21981 15519 22015
rect 21833 21981 21867 22015
rect 22201 21981 22235 22015
rect 22569 21981 22603 22015
rect 23121 21981 23155 22015
rect 7021 21913 7055 21947
rect 7481 21913 7515 21947
rect 8493 21913 8527 21947
rect 9689 21913 9723 21947
rect 10517 21913 10551 21947
rect 12449 21913 12483 21947
rect 12633 21913 12667 21947
rect 12817 21913 12851 21947
rect 14565 21913 14599 21947
rect 16221 21913 16255 21947
rect 16957 21913 16991 21947
rect 17877 21913 17911 21947
rect 1777 21845 1811 21879
rect 2421 21845 2455 21879
rect 3065 21845 3099 21879
rect 3433 21845 3467 21879
rect 3893 21845 3927 21879
rect 4445 21845 4479 21879
rect 4813 21845 4847 21879
rect 5089 21845 5123 21879
rect 5641 21845 5675 21879
rect 5917 21845 5951 21879
rect 6009 21845 6043 21879
rect 6377 21845 6411 21879
rect 6561 21845 6595 21879
rect 6929 21845 6963 21879
rect 7573 21845 7607 21879
rect 7941 21845 7975 21879
rect 8033 21845 8067 21879
rect 8401 21845 8435 21879
rect 9045 21845 9079 21879
rect 9597 21845 9631 21879
rect 10057 21845 10091 21879
rect 10425 21845 10459 21879
rect 11069 21845 11103 21879
rect 11345 21845 11379 21879
rect 11621 21845 11655 21879
rect 11989 21845 12023 21879
rect 13093 21845 13127 21879
rect 13829 21845 13863 21879
rect 15209 21845 15243 21879
rect 15669 21845 15703 21879
rect 15761 21845 15795 21879
rect 16129 21845 16163 21879
rect 17049 21845 17083 21879
rect 17417 21845 17451 21879
rect 17785 21845 17819 21879
rect 18245 21845 18279 21879
rect 18613 21845 18647 21879
rect 18705 21845 18739 21879
rect 19073 21845 19107 21879
rect 19625 21845 19659 21879
rect 19717 21845 19751 21879
rect 20361 21845 20395 21879
rect 20453 21845 20487 21879
rect 21281 21845 21315 21879
rect 21373 21845 21407 21879
rect 22385 21845 22419 21879
rect 22753 21845 22787 21879
rect 22937 21845 22971 21879
rect 1501 21641 1535 21675
rect 2145 21641 2179 21675
rect 2421 21641 2455 21675
rect 2881 21641 2915 21675
rect 3525 21641 3559 21675
rect 4353 21641 4387 21675
rect 5917 21641 5951 21675
rect 8585 21641 8619 21675
rect 9413 21641 9447 21675
rect 11805 21641 11839 21675
rect 12265 21641 12299 21675
rect 14565 21641 14599 21675
rect 16037 21641 16071 21675
rect 17049 21641 17083 21675
rect 17417 21641 17451 21675
rect 18711 21641 18745 21675
rect 20545 21641 20579 21675
rect 20913 21641 20947 21675
rect 22017 21641 22051 21675
rect 22201 21641 22235 21675
rect 22661 21641 22695 21675
rect 2789 21573 2823 21607
rect 6561 21573 6595 21607
rect 9045 21573 9079 21607
rect 12633 21573 12667 21607
rect 17693 21573 17727 21607
rect 1685 21505 1719 21539
rect 2053 21505 2087 21539
rect 2329 21505 2363 21539
rect 2605 21505 2639 21539
rect 3065 21505 3099 21539
rect 3433 21505 3467 21539
rect 3709 21505 3743 21539
rect 3801 21505 3835 21539
rect 4077 21505 4111 21539
rect 4537 21505 4571 21539
rect 4629 21505 4663 21539
rect 5089 21505 5123 21539
rect 5365 21505 5399 21539
rect 5641 21505 5675 21539
rect 6837 21505 6871 21539
rect 7389 21505 7423 21539
rect 8217 21505 8251 21539
rect 10241 21505 10275 21539
rect 11897 21505 11931 21539
rect 12449 21505 12483 21539
rect 14933 21505 14967 21539
rect 15025 21505 15059 21539
rect 16957 21505 16991 21539
rect 17509 21505 17543 21539
rect 18153 21505 18187 21539
rect 21005 21505 21039 21539
rect 21373 21505 21407 21539
rect 21833 21505 21867 21539
rect 22385 21505 22419 21539
rect 22477 21505 22511 21539
rect 22845 21505 22879 21539
rect 6193 21437 6227 21471
rect 7481 21437 7515 21471
rect 7573 21437 7607 21471
rect 7941 21437 7975 21471
rect 8125 21437 8159 21471
rect 8769 21437 8803 21471
rect 8953 21437 8987 21471
rect 9505 21437 9539 21471
rect 9828 21437 9862 21471
rect 10011 21437 10045 21471
rect 11713 21437 11747 21471
rect 12725 21437 12759 21471
rect 13048 21437 13082 21471
rect 13188 21437 13222 21471
rect 13461 21437 13495 21471
rect 14749 21437 14783 21471
rect 15853 21437 15887 21471
rect 15945 21437 15979 21471
rect 16773 21437 16807 21471
rect 18245 21437 18279 21471
rect 18751 21439 18785 21473
rect 18981 21437 19015 21471
rect 20269 21437 20303 21471
rect 20453 21437 20487 21471
rect 1869 21369 1903 21403
rect 3249 21369 3283 21403
rect 4813 21369 4847 21403
rect 5181 21369 5215 21403
rect 6653 21369 6687 21403
rect 15393 21369 15427 21403
rect 17969 21369 18003 21403
rect 21557 21369 21591 21403
rect 3985 21301 4019 21335
rect 4261 21301 4295 21335
rect 4905 21301 4939 21335
rect 5457 21301 5491 21335
rect 7021 21301 7055 21335
rect 11345 21301 11379 21335
rect 15577 21301 15611 21335
rect 16405 21301 16439 21335
rect 17877 21301 17911 21335
rect 20085 21301 20119 21335
rect 21189 21301 21223 21335
rect 23029 21301 23063 21335
rect 2513 21097 2547 21131
rect 2789 21097 2823 21131
rect 3065 21097 3099 21131
rect 3341 21097 3375 21131
rect 6009 21097 6043 21131
rect 11069 21097 11103 21131
rect 20729 21097 20763 21131
rect 22661 21097 22695 21131
rect 6929 21029 6963 21063
rect 10793 21029 10827 21063
rect 13737 21029 13771 21063
rect 13921 21029 13955 21063
rect 14841 21029 14875 21063
rect 21557 21029 21591 21063
rect 2973 20961 3007 20995
rect 5457 20961 5491 20995
rect 6193 20961 6227 20995
rect 6377 20961 6411 20995
rect 8306 20961 8340 20995
rect 9416 20961 9450 20995
rect 9689 20961 9723 20995
rect 12403 20961 12437 20995
rect 13093 20961 13127 20995
rect 14197 20961 14231 20995
rect 14381 20961 14415 20995
rect 15577 20961 15611 20995
rect 16497 20961 16531 20995
rect 18337 20961 18371 20995
rect 18610 20961 18644 20995
rect 21189 20961 21223 20995
rect 21281 20961 21315 20995
rect 22109 20961 22143 20995
rect 2053 20893 2087 20927
rect 2237 20893 2271 20927
rect 3617 20893 3651 20927
rect 3893 20893 3927 20927
rect 4353 20893 4387 20927
rect 4905 20893 4939 20927
rect 5181 20893 5215 20927
rect 5641 20893 5675 20927
rect 6469 20893 6503 20927
rect 8033 20893 8067 20927
rect 8769 20893 8803 20927
rect 8953 20893 8987 20927
rect 12173 20893 12207 20927
rect 12909 20893 12943 20927
rect 15393 20893 15427 20927
rect 15945 20893 15979 20927
rect 16129 20893 16163 20927
rect 16773 20893 16807 20927
rect 19073 20893 19107 20927
rect 20637 20893 20671 20927
rect 22477 20893 22511 20927
rect 22845 20893 22879 20927
rect 2421 20825 2455 20859
rect 4629 20825 4663 20859
rect 15301 20825 15335 20859
rect 16313 20825 16347 20859
rect 16681 20825 16715 20859
rect 20370 20825 20404 20859
rect 3433 20757 3467 20791
rect 4077 20757 4111 20791
rect 4261 20757 4295 20791
rect 4721 20757 4755 20791
rect 4997 20757 5031 20791
rect 5549 20757 5583 20791
rect 6837 20757 6871 20791
rect 8302 20757 8336 20791
rect 9419 20757 9453 20791
rect 10885 20757 10919 20791
rect 12442 20757 12476 20791
rect 13277 20757 13311 20791
rect 13369 20757 13403 20791
rect 14473 20757 14507 20791
rect 14933 20757 14967 20791
rect 15761 20757 15795 20791
rect 17141 20757 17175 20791
rect 17233 20757 17267 20791
rect 18606 20757 18640 20791
rect 19257 20757 19291 20791
rect 21097 20757 21131 20791
rect 21925 20757 21959 20791
rect 22017 20757 22051 20791
rect 23029 20757 23063 20791
rect 2421 20553 2455 20587
rect 2881 20553 2915 20587
rect 3065 20553 3099 20587
rect 3985 20553 4019 20587
rect 5089 20553 5123 20587
rect 6009 20553 6043 20587
rect 8125 20553 8159 20587
rect 8953 20553 8987 20587
rect 9505 20553 9539 20587
rect 9965 20553 9999 20587
rect 11345 20553 11379 20587
rect 13461 20553 13495 20587
rect 13921 20553 13955 20587
rect 14289 20553 14323 20587
rect 15945 20553 15979 20587
rect 20177 20553 20211 20587
rect 21465 20553 21499 20587
rect 21833 20553 21867 20587
rect 22293 20553 22327 20587
rect 3249 20485 3283 20519
rect 9413 20485 9447 20519
rect 14657 20485 14691 20519
rect 17877 20485 17911 20519
rect 18604 20485 18638 20519
rect 20913 20485 20947 20519
rect 3893 20417 3927 20451
rect 4721 20417 4755 20451
rect 5641 20417 5675 20451
rect 7490 20417 7524 20451
rect 7757 20417 7791 20451
rect 8585 20417 8619 20451
rect 10241 20417 10275 20451
rect 10701 20417 10735 20451
rect 11852 20417 11886 20451
rect 13829 20417 13863 20451
rect 15577 20417 15611 20451
rect 16405 20417 16439 20451
rect 17049 20417 17083 20451
rect 20085 20417 20119 20451
rect 21005 20417 21039 20451
rect 21649 20417 21683 20451
rect 22109 20417 22143 20451
rect 22477 20417 22511 20451
rect 22845 20417 22879 20451
rect 3433 20349 3467 20383
rect 4077 20349 4111 20383
rect 4445 20349 4479 20383
rect 4629 20349 4663 20383
rect 5917 20349 5951 20383
rect 8309 20349 8343 20383
rect 8493 20349 8527 20383
rect 9597 20349 9631 20383
rect 10425 20349 10459 20383
rect 10609 20349 10643 20383
rect 11529 20349 11563 20383
rect 12035 20349 12069 20383
rect 12265 20349 12299 20383
rect 14013 20349 14047 20383
rect 14749 20349 14783 20383
rect 14933 20349 14967 20383
rect 15301 20349 15335 20383
rect 15485 20349 15519 20383
rect 17141 20349 17175 20383
rect 17233 20349 17267 20383
rect 17969 20349 18003 20383
rect 18153 20349 18187 20383
rect 18337 20349 18371 20383
rect 19901 20349 19935 20383
rect 20821 20349 20855 20383
rect 5457 20281 5491 20315
rect 9045 20281 9079 20315
rect 13369 20281 13403 20315
rect 16221 20281 16255 20315
rect 19717 20281 19751 20315
rect 20545 20281 20579 20315
rect 22661 20281 22695 20315
rect 3525 20213 3559 20247
rect 5365 20213 5399 20247
rect 6377 20213 6411 20247
rect 10057 20213 10091 20247
rect 11069 20213 11103 20247
rect 16037 20213 16071 20247
rect 16681 20213 16715 20247
rect 17509 20213 17543 20247
rect 21373 20213 21407 20247
rect 23029 20213 23063 20247
rect 4169 20009 4203 20043
rect 4353 20009 4387 20043
rect 8585 20009 8619 20043
rect 10333 20009 10367 20043
rect 12449 20009 12483 20043
rect 13921 20009 13955 20043
rect 21833 20009 21867 20043
rect 16221 19941 16255 19975
rect 4813 19873 4847 19907
rect 4997 19873 5031 19907
rect 12541 19873 12575 19907
rect 13277 19873 13311 19907
rect 13461 19873 13495 19907
rect 14105 19873 14139 19907
rect 16405 19873 16439 19907
rect 17325 19873 17359 19907
rect 20913 19873 20947 19907
rect 22109 19873 22143 19907
rect 3617 19805 3651 19839
rect 3985 19805 4019 19839
rect 4721 19805 4755 19839
rect 5549 19805 5583 19839
rect 7113 19805 7147 19839
rect 7205 19805 7239 19839
rect 8677 19805 8711 19839
rect 8953 19805 8987 19839
rect 10609 19805 10643 19839
rect 12081 19805 12115 19839
rect 12265 19805 12299 19839
rect 12909 19805 12943 19839
rect 14841 19805 14875 19839
rect 17417 19805 17451 19839
rect 17693 19805 17727 19839
rect 19257 19805 19291 19839
rect 21005 19805 21039 19839
rect 21649 19805 21683 19839
rect 22845 19805 22879 19839
rect 5365 19737 5399 19771
rect 6846 19737 6880 19771
rect 7450 19737 7484 19771
rect 9198 19737 9232 19771
rect 11836 19737 11870 19771
rect 13553 19737 13587 19771
rect 14381 19737 14415 19771
rect 15108 19737 15142 19771
rect 17960 19737 17994 19771
rect 19524 19737 19558 19771
rect 21097 19737 21131 19771
rect 3433 19669 3467 19703
rect 3801 19669 3835 19703
rect 5273 19669 5307 19703
rect 5733 19669 5767 19703
rect 10425 19669 10459 19703
rect 10701 19669 10735 19703
rect 13093 19669 13127 19703
rect 14657 19669 14691 19703
rect 16589 19669 16623 19703
rect 16681 19669 16715 19703
rect 17049 19669 17083 19703
rect 17601 19669 17635 19703
rect 19073 19669 19107 19703
rect 20637 19669 20671 19703
rect 21465 19669 21499 19703
rect 22293 19669 22327 19703
rect 22385 19669 22419 19703
rect 22753 19669 22787 19703
rect 23029 19669 23063 19703
rect 3065 19465 3099 19499
rect 3525 19465 3559 19499
rect 4353 19465 4387 19499
rect 4629 19465 4663 19499
rect 7849 19465 7883 19499
rect 9505 19465 9539 19499
rect 10977 19465 11011 19499
rect 11161 19465 11195 19499
rect 11529 19465 11563 19499
rect 13277 19465 13311 19499
rect 13553 19465 13587 19499
rect 14381 19465 14415 19499
rect 15853 19465 15887 19499
rect 16129 19465 16163 19499
rect 16681 19465 16715 19499
rect 18153 19465 18187 19499
rect 19625 19465 19659 19499
rect 21097 19465 21131 19499
rect 22293 19465 22327 19499
rect 17794 19397 17828 19431
rect 22201 19397 22235 19431
rect 3157 19329 3191 19363
rect 3893 19329 3927 19363
rect 3985 19329 4019 19363
rect 4445 19329 4479 19363
rect 5937 19329 5971 19363
rect 6193 19329 6227 19363
rect 6377 19329 6411 19363
rect 6633 19329 6667 19363
rect 8033 19329 8067 19363
rect 8125 19329 8159 19363
rect 8392 19329 8426 19363
rect 9597 19329 9631 19363
rect 9853 19329 9887 19363
rect 11345 19329 11379 19363
rect 12653 19329 12687 19363
rect 12909 19329 12943 19363
rect 13093 19329 13127 19363
rect 13369 19329 13403 19363
rect 13921 19329 13955 19363
rect 14013 19329 14047 19363
rect 14473 19329 14507 19363
rect 14740 19329 14774 19363
rect 15945 19329 15979 19363
rect 16405 19329 16439 19363
rect 18061 19329 18095 19363
rect 19277 19329 19311 19363
rect 19533 19329 19567 19363
rect 20749 19329 20783 19363
rect 21005 19329 21039 19363
rect 21281 19329 21315 19363
rect 21373 19329 21407 19363
rect 22845 19329 22879 19363
rect 2973 19261 3007 19295
rect 3801 19261 3835 19295
rect 13829 19261 13863 19295
rect 22477 19261 22511 19295
rect 22753 19261 22787 19295
rect 16221 19193 16255 19227
rect 21557 19193 21591 19227
rect 21833 19193 21867 19227
rect 2697 19125 2731 19159
rect 4813 19125 4847 19159
rect 7757 19125 7791 19159
rect 23029 19125 23063 19159
rect 3801 18921 3835 18955
rect 8769 18921 8803 18955
rect 12449 18921 12483 18955
rect 12541 18921 12575 18955
rect 15485 18921 15519 18955
rect 17049 18921 17083 18955
rect 18521 18921 18555 18955
rect 18797 18921 18831 18955
rect 3617 18853 3651 18887
rect 16957 18853 16991 18887
rect 20729 18853 20763 18887
rect 3065 18785 3099 18819
rect 5825 18785 5859 18819
rect 8953 18785 8987 18819
rect 18429 18785 18463 18819
rect 22661 18785 22695 18819
rect 22753 18785 22787 18819
rect 2789 18717 2823 18751
rect 3985 18717 4019 18751
rect 4353 18717 4387 18751
rect 5558 18717 5592 18751
rect 7297 18717 7331 18751
rect 7389 18717 7423 18751
rect 9229 18717 9263 18751
rect 9413 18717 9447 18751
rect 9597 18717 9631 18751
rect 9864 18717 9898 18751
rect 11069 18717 11103 18751
rect 11325 18717 11359 18751
rect 13921 18717 13955 18751
rect 14105 18717 14139 18751
rect 15577 18717 15611 18751
rect 18705 18717 18739 18751
rect 18981 18717 19015 18751
rect 20637 18717 20671 18751
rect 21842 18717 21876 18751
rect 22109 18717 22143 18751
rect 23029 18717 23063 18751
rect 3249 18649 3283 18683
rect 4169 18649 4203 18683
rect 7030 18649 7064 18683
rect 7656 18649 7690 18683
rect 13676 18649 13710 18683
rect 14372 18649 14406 18683
rect 15844 18649 15878 18683
rect 18162 18649 18196 18683
rect 20392 18649 20426 18683
rect 22569 18649 22603 18683
rect 2605 18581 2639 18615
rect 3157 18581 3191 18615
rect 4445 18581 4479 18615
rect 5917 18581 5951 18615
rect 10977 18581 11011 18615
rect 19257 18581 19291 18615
rect 22201 18581 22235 18615
rect 2053 18377 2087 18411
rect 3985 18377 4019 18411
rect 4445 18377 4479 18411
rect 4905 18377 4939 18411
rect 5273 18377 5307 18411
rect 7849 18377 7883 18411
rect 8125 18377 8159 18411
rect 8309 18377 8343 18411
rect 8493 18377 8527 18411
rect 11529 18377 11563 18411
rect 14657 18377 14691 18411
rect 16681 18377 16715 18411
rect 17417 18377 17451 18411
rect 21833 18377 21867 18411
rect 22293 18377 22327 18411
rect 22753 18377 22787 18411
rect 5365 18309 5399 18343
rect 9628 18309 9662 18343
rect 11980 18309 12014 18343
rect 22845 18309 22879 18343
rect 1869 18241 1903 18275
rect 2145 18241 2179 18275
rect 2789 18241 2823 18275
rect 2881 18241 2915 18275
rect 3617 18241 3651 18275
rect 5827 18241 5861 18275
rect 6633 18241 6667 18275
rect 9873 18241 9907 18275
rect 9965 18241 9999 18275
rect 10232 18241 10266 18275
rect 11713 18241 11747 18275
rect 14298 18241 14332 18275
rect 14565 18241 14599 18275
rect 15770 18241 15804 18275
rect 16129 18241 16163 18275
rect 17233 18241 17267 18275
rect 17601 18241 17635 18275
rect 18429 18241 18463 18275
rect 18797 18241 18831 18275
rect 19064 18241 19098 18275
rect 20525 18241 20559 18275
rect 22201 18241 22235 18275
rect 2973 18173 3007 18207
rect 3341 18173 3375 18207
rect 3525 18173 3559 18207
rect 4261 18173 4295 18207
rect 4353 18173 4387 18207
rect 5457 18173 5491 18207
rect 6377 18173 6411 18207
rect 16037 18173 16071 18207
rect 18245 18173 18279 18207
rect 20269 18173 20303 18207
rect 22477 18173 22511 18207
rect 2421 18105 2455 18139
rect 6009 18105 6043 18139
rect 7757 18105 7791 18139
rect 11345 18105 11379 18139
rect 13093 18105 13127 18139
rect 13185 18105 13219 18139
rect 20177 18105 20211 18139
rect 23029 18105 23063 18139
rect 2329 18037 2363 18071
rect 4813 18037 4847 18071
rect 6101 18037 6135 18071
rect 16313 18037 16347 18071
rect 16405 18037 16439 18071
rect 17693 18037 17727 18071
rect 21649 18037 21683 18071
rect 3801 17833 3835 17867
rect 5917 17833 5951 17867
rect 9689 17833 9723 17867
rect 13921 17833 13955 17867
rect 15485 17833 15519 17867
rect 17325 17833 17359 17867
rect 19073 17833 19107 17867
rect 21741 17833 21775 17867
rect 22753 17833 22787 17867
rect 19257 17765 19291 17799
rect 2789 17697 2823 17731
rect 2973 17697 3007 17731
rect 16957 17697 16991 17731
rect 20913 17697 20947 17731
rect 22017 17697 22051 17731
rect 3065 17629 3099 17663
rect 3985 17629 4019 17663
rect 4169 17629 4203 17663
rect 4445 17629 4479 17663
rect 7297 17629 7331 17663
rect 8769 17629 8803 17663
rect 9045 17629 9079 17663
rect 9229 17629 9263 17663
rect 9413 17629 9447 17663
rect 9597 17629 9631 17663
rect 11069 17629 11103 17663
rect 11253 17629 11287 17663
rect 11529 17629 11563 17663
rect 11805 17629 11839 17663
rect 11989 17629 12023 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 13737 17629 13771 17663
rect 14105 17629 14139 17663
rect 17141 17629 17175 17663
rect 17693 17629 17727 17663
rect 20637 17629 20671 17663
rect 21557 17629 21591 17663
rect 22845 17629 22879 17663
rect 4712 17561 4746 17595
rect 7030 17561 7064 17595
rect 8502 17561 8536 17595
rect 10802 17561 10836 17595
rect 12532 17561 12566 17595
rect 14372 17561 14406 17595
rect 16690 17561 16724 17595
rect 17960 17561 17994 17595
rect 20370 17561 20404 17595
rect 22109 17561 22143 17595
rect 3433 17493 3467 17527
rect 4353 17493 4387 17527
rect 5825 17493 5859 17527
rect 7389 17493 7423 17527
rect 13645 17493 13679 17527
rect 15577 17493 15611 17527
rect 17601 17493 17635 17527
rect 21005 17493 21039 17527
rect 21097 17493 21131 17527
rect 21465 17493 21499 17527
rect 22201 17493 22235 17527
rect 22569 17493 22603 17527
rect 23121 17493 23155 17527
rect 3893 17289 3927 17323
rect 6745 17289 6779 17323
rect 9045 17289 9079 17323
rect 10517 17289 10551 17323
rect 10701 17289 10735 17323
rect 10885 17289 10919 17323
rect 11069 17289 11103 17323
rect 11253 17289 11287 17323
rect 14197 17289 14231 17323
rect 16221 17289 16255 17323
rect 16681 17289 16715 17323
rect 18153 17289 18187 17323
rect 18613 17289 18647 17323
rect 18705 17289 18739 17323
rect 20545 17289 20579 17323
rect 21005 17289 21039 17323
rect 21649 17289 21683 17323
rect 23029 17289 23063 17323
rect 4169 17221 4203 17255
rect 5080 17221 5114 17255
rect 13185 17221 13219 17255
rect 13461 17221 13495 17255
rect 17794 17221 17828 17255
rect 21373 17221 21407 17255
rect 22201 17221 22235 17255
rect 3709 17153 3743 17187
rect 4353 17153 4387 17187
rect 4721 17153 4755 17187
rect 7932 17153 7966 17187
rect 9137 17153 9171 17187
rect 9393 17153 9427 17187
rect 12734 17153 12768 17187
rect 13001 17153 13035 17187
rect 13645 17153 13679 17187
rect 13921 17153 13955 17187
rect 14013 17153 14047 17187
rect 14289 17153 14323 17187
rect 14565 17153 14599 17187
rect 14821 17153 14855 17187
rect 16037 17153 16071 17187
rect 18061 17153 18095 17187
rect 18337 17153 18371 17187
rect 18429 17153 18463 17187
rect 19818 17153 19852 17187
rect 20637 17153 20671 17187
rect 22293 17153 22327 17187
rect 22753 17153 22787 17187
rect 3985 17085 4019 17119
rect 4813 17085 4847 17119
rect 6837 17085 6871 17119
rect 6929 17085 6963 17119
rect 7665 17085 7699 17119
rect 16497 17085 16531 17119
rect 20085 17085 20119 17119
rect 20453 17085 20487 17119
rect 22109 17085 22143 17119
rect 6377 17017 6411 17051
rect 11621 17017 11655 17051
rect 13737 17017 13771 17051
rect 14473 17017 14507 17051
rect 22937 17017 22971 17051
rect 4537 16949 4571 16983
rect 6193 16949 6227 16983
rect 7205 16949 7239 16983
rect 7389 16949 7423 16983
rect 15945 16949 15979 16983
rect 21281 16949 21315 16983
rect 22661 16949 22695 16983
rect 4169 16745 4203 16779
rect 4997 16745 5031 16779
rect 8033 16745 8067 16779
rect 12541 16745 12575 16779
rect 18429 16745 18463 16779
rect 20637 16745 20671 16779
rect 21557 16745 21591 16779
rect 22477 16745 22511 16779
rect 23029 16745 23063 16779
rect 5181 16677 5215 16711
rect 14105 16677 14139 16711
rect 18797 16677 18831 16711
rect 4721 16609 4755 16643
rect 6561 16609 6595 16643
rect 6653 16609 6687 16643
rect 9781 16609 9815 16643
rect 21005 16609 21039 16643
rect 22201 16609 22235 16643
rect 6294 16541 6328 16575
rect 10149 16541 10183 16575
rect 11621 16541 11655 16575
rect 11805 16541 11839 16575
rect 11989 16541 12023 16575
rect 12173 16541 12207 16575
rect 13921 16541 13955 16575
rect 15485 16541 15519 16575
rect 16690 16541 16724 16575
rect 16957 16541 16991 16575
rect 17049 16541 17083 16575
rect 17316 16541 17350 16575
rect 18613 16541 18647 16575
rect 18889 16541 18923 16575
rect 19257 16541 19291 16575
rect 19524 16541 19558 16575
rect 21097 16541 21131 16575
rect 22661 16541 22695 16575
rect 22937 16541 22971 16575
rect 6898 16473 6932 16507
rect 9597 16473 9631 16507
rect 10416 16473 10450 16507
rect 12357 16473 12391 16507
rect 13654 16473 13688 16507
rect 15218 16473 15252 16507
rect 4537 16405 4571 16439
rect 4629 16405 4663 16439
rect 8125 16405 8159 16439
rect 8309 16405 8343 16439
rect 9229 16405 9263 16439
rect 9689 16405 9723 16439
rect 11529 16405 11563 16439
rect 15577 16405 15611 16439
rect 19073 16405 19107 16439
rect 21189 16405 21223 16439
rect 21649 16405 21683 16439
rect 22017 16405 22051 16439
rect 22109 16405 22143 16439
rect 22753 16405 22787 16439
rect 3985 16201 4019 16235
rect 4353 16201 4387 16235
rect 8493 16201 8527 16235
rect 8861 16201 8895 16235
rect 16129 16201 16163 16235
rect 18061 16201 18095 16235
rect 18705 16201 18739 16235
rect 20637 16201 20671 16235
rect 21005 16201 21039 16235
rect 21373 16201 21407 16235
rect 21649 16201 21683 16235
rect 22569 16201 22603 16235
rect 10793 16133 10827 16167
rect 11805 16133 11839 16167
rect 11989 16133 12023 16167
rect 12357 16133 12391 16167
rect 12541 16133 12575 16167
rect 14197 16133 14231 16167
rect 14381 16133 14415 16167
rect 15016 16133 15050 16167
rect 16948 16133 16982 16167
rect 19840 16133 19874 16167
rect 22201 16133 22235 16167
rect 3433 16065 3467 16099
rect 3709 16065 3743 16099
rect 4445 16065 4479 16099
rect 5926 16065 5960 16099
rect 6193 16065 6227 16099
rect 7593 16065 7627 16099
rect 7849 16065 7883 16099
rect 7941 16065 7975 16099
rect 8125 16065 8159 16099
rect 9321 16065 9355 16099
rect 9577 16065 9611 16099
rect 11161 16065 11195 16099
rect 11345 16065 11379 16099
rect 11621 16065 11655 16099
rect 12725 16065 12759 16099
rect 12981 16065 13015 16099
rect 14749 16065 14783 16099
rect 16313 16065 16347 16099
rect 16681 16065 16715 16099
rect 18429 16065 18463 16099
rect 21189 16065 21223 16099
rect 21465 16065 21499 16099
rect 22845 16065 22879 16099
rect 22937 16065 22971 16099
rect 4537 15997 4571 16031
rect 8953 15997 8987 16031
rect 9045 15997 9079 16031
rect 18337 15997 18371 16031
rect 20085 15997 20119 16031
rect 20361 15997 20395 16031
rect 20545 15997 20579 16031
rect 22017 15997 22051 16031
rect 22109 15997 22143 16031
rect 3617 15929 3651 15963
rect 4813 15929 4847 15963
rect 6469 15929 6503 15963
rect 16497 15929 16531 15963
rect 3893 15861 3927 15895
rect 10701 15861 10735 15895
rect 12265 15861 12299 15895
rect 14105 15861 14139 15895
rect 14565 15861 14599 15895
rect 18613 15861 18647 15895
rect 22661 15861 22695 15895
rect 23121 15861 23155 15895
rect 4261 15657 4295 15691
rect 5089 15657 5123 15691
rect 6653 15657 6687 15691
rect 12817 15657 12851 15691
rect 13093 15657 13127 15691
rect 15945 15657 15979 15691
rect 16221 15657 16255 15691
rect 18245 15657 18279 15691
rect 20637 15657 20671 15691
rect 22385 15657 22419 15691
rect 6745 15589 6779 15623
rect 14565 15589 14599 15623
rect 16037 15589 16071 15623
rect 22477 15589 22511 15623
rect 4813 15521 4847 15555
rect 5273 15521 5307 15555
rect 8125 15521 8159 15555
rect 8309 15521 8343 15555
rect 8493 15521 8527 15555
rect 9597 15521 9631 15555
rect 15301 15521 15335 15555
rect 15485 15521 15519 15555
rect 18705 15521 18739 15555
rect 18797 15521 18831 15555
rect 19257 15521 19291 15555
rect 21005 15521 21039 15555
rect 21741 15521 21775 15555
rect 23029 15521 23063 15555
rect 1685 15453 1719 15487
rect 4721 15453 4755 15487
rect 11069 15453 11103 15487
rect 11437 15453 11471 15487
rect 11693 15453 11727 15487
rect 12909 15453 12943 15487
rect 13553 15453 13587 15487
rect 16405 15453 16439 15487
rect 16497 15453 16531 15487
rect 18153 15453 18187 15487
rect 22661 15453 22695 15487
rect 22937 15453 22971 15487
rect 5518 15385 5552 15419
rect 7858 15385 7892 15419
rect 9842 15385 9876 15419
rect 13277 15385 13311 15419
rect 13737 15385 13771 15419
rect 13921 15385 13955 15419
rect 14197 15385 14231 15419
rect 14381 15385 14415 15419
rect 14749 15385 14783 15419
rect 14933 15385 14967 15419
rect 15117 15385 15151 15419
rect 17886 15385 17920 15419
rect 18613 15385 18647 15419
rect 19524 15385 19558 15419
rect 22017 15385 22051 15419
rect 1501 15317 1535 15351
rect 4629 15317 4663 15351
rect 10977 15317 11011 15351
rect 15577 15317 15611 15351
rect 16681 15317 16715 15351
rect 16773 15317 16807 15351
rect 21097 15317 21131 15351
rect 21189 15317 21223 15351
rect 21557 15317 21591 15351
rect 21925 15317 21959 15351
rect 22753 15317 22787 15351
rect 8401 15113 8435 15147
rect 8769 15113 8803 15147
rect 12909 15113 12943 15147
rect 13185 15113 13219 15147
rect 13461 15113 13495 15147
rect 14381 15113 14415 15147
rect 21649 15113 21683 15147
rect 22477 15113 22511 15147
rect 22569 15113 22603 15147
rect 7104 15045 7138 15079
rect 8861 15045 8895 15079
rect 21281 15045 21315 15079
rect 4905 14977 4939 15011
rect 5641 14977 5675 15011
rect 6469 14977 6503 15011
rect 6837 14977 6871 15011
rect 11078 14977 11112 15011
rect 11345 14977 11379 15011
rect 11897 14977 11931 15011
rect 14289 14977 14323 15011
rect 15494 14977 15528 15011
rect 15761 14977 15795 15011
rect 15945 14977 15979 15011
rect 16313 14977 16347 15011
rect 16681 14977 16715 15011
rect 16937 14977 16971 15011
rect 18153 14977 18187 15011
rect 18420 14977 18454 15011
rect 20738 14977 20772 15011
rect 21465 14977 21499 15011
rect 21833 14977 21867 15011
rect 23121 14977 23155 15011
rect 5365 14909 5399 14943
rect 9045 14909 9079 14943
rect 11989 14909 12023 14943
rect 12173 14909 12207 14943
rect 21005 14909 21039 14943
rect 22661 14909 22695 14943
rect 9965 14841 9999 14875
rect 16405 14841 16439 14875
rect 18061 14841 18095 14875
rect 19533 14841 19567 14875
rect 5089 14773 5123 14807
rect 6561 14773 6595 14807
rect 8217 14773 8251 14807
rect 11529 14773 11563 14807
rect 12817 14773 12851 14807
rect 13277 14773 13311 14807
rect 13645 14773 13679 14807
rect 16037 14773 16071 14807
rect 19625 14773 19659 14807
rect 21097 14773 21131 14807
rect 22017 14773 22051 14807
rect 22109 14773 22143 14807
rect 22937 14773 22971 14807
rect 6929 14569 6963 14603
rect 8401 14569 8435 14603
rect 8585 14569 8619 14603
rect 11345 14569 11379 14603
rect 11437 14569 11471 14603
rect 11621 14569 11655 14603
rect 16957 14569 16991 14603
rect 18429 14569 18463 14603
rect 18797 14569 18831 14603
rect 20637 14569 20671 14603
rect 11161 14501 11195 14535
rect 16221 14501 16255 14535
rect 18889 14501 18923 14535
rect 21833 14501 21867 14535
rect 5089 14433 5123 14467
rect 5273 14433 5307 14467
rect 8309 14433 8343 14467
rect 9597 14433 9631 14467
rect 9781 14433 9815 14467
rect 13737 14433 13771 14467
rect 16129 14433 16163 14467
rect 18337 14433 18371 14467
rect 19257 14433 19291 14467
rect 21281 14433 21315 14467
rect 22477 14433 22511 14467
rect 22569 14433 22603 14467
rect 5457 14365 5491 14399
rect 12745 14365 12779 14399
rect 13001 14365 13035 14399
rect 14289 14365 14323 14399
rect 14381 14365 14415 14399
rect 14565 14365 14599 14399
rect 16773 14365 16807 14399
rect 18613 14365 18647 14399
rect 19073 14365 19107 14399
rect 19524 14365 19558 14399
rect 21557 14365 21591 14399
rect 21649 14365 21683 14399
rect 23029 14365 23063 14399
rect 4997 14297 5031 14331
rect 5724 14297 5758 14331
rect 8042 14297 8076 14331
rect 9321 14297 9355 14331
rect 10048 14297 10082 14331
rect 13645 14297 13679 14331
rect 15862 14297 15896 14331
rect 18070 14297 18104 14331
rect 4629 14229 4663 14263
rect 6837 14229 6871 14263
rect 8953 14229 8987 14263
rect 9413 14229 9447 14263
rect 13185 14229 13219 14263
rect 13553 14229 13587 14263
rect 14749 14229 14783 14263
rect 16497 14229 16531 14263
rect 16681 14229 16715 14263
rect 22017 14229 22051 14263
rect 22385 14229 22419 14263
rect 22937 14229 22971 14263
rect 1869 14025 1903 14059
rect 4721 14025 4755 14059
rect 9689 14025 9723 14059
rect 11253 14025 11287 14059
rect 11529 14025 11563 14059
rect 13185 14025 13219 14059
rect 14657 14025 14691 14059
rect 14841 14025 14875 14059
rect 15393 14025 15427 14059
rect 15945 14025 15979 14059
rect 16037 14025 16071 14059
rect 16405 14025 16439 14059
rect 17049 14025 17083 14059
rect 19625 14025 19659 14059
rect 21097 14025 21131 14059
rect 22201 14025 22235 14059
rect 22845 14025 22879 14059
rect 4813 13957 4847 13991
rect 10118 13957 10152 13991
rect 12050 13957 12084 13991
rect 15025 13957 15059 13991
rect 15577 13957 15611 13991
rect 21373 13957 21407 13991
rect 2053 13889 2087 13923
rect 4353 13889 4387 13923
rect 5641 13889 5675 13923
rect 6653 13889 6687 13923
rect 6920 13889 6954 13923
rect 8125 13889 8159 13923
rect 8392 13889 8426 13923
rect 9873 13889 9907 13923
rect 11805 13889 11839 13923
rect 13277 13889 13311 13923
rect 13544 13889 13578 13923
rect 15761 13889 15795 13923
rect 16313 13889 16347 13923
rect 18245 13889 18279 13923
rect 18512 13889 18546 13923
rect 19984 13889 20018 13923
rect 22661 13889 22695 13923
rect 23121 13889 23155 13923
rect 2145 13821 2179 13855
rect 4629 13821 4663 13855
rect 5733 13821 5767 13855
rect 5917 13821 5951 13855
rect 17141 13821 17175 13855
rect 17325 13821 17359 13855
rect 19717 13821 19751 13855
rect 21925 13821 21959 13855
rect 22109 13821 22143 13855
rect 15209 13753 15243 13787
rect 16681 13753 16715 13787
rect 17601 13753 17635 13787
rect 17693 13753 17727 13787
rect 17969 13753 18003 13787
rect 18061 13753 18095 13787
rect 21557 13753 21591 13787
rect 22937 13753 22971 13787
rect 4169 13685 4203 13719
rect 5181 13685 5215 13719
rect 5273 13685 5307 13719
rect 8033 13685 8067 13719
rect 9505 13685 9539 13719
rect 21281 13685 21315 13719
rect 22569 13685 22603 13719
rect 3801 13481 3835 13515
rect 4629 13481 4663 13515
rect 6561 13481 6595 13515
rect 8125 13481 8159 13515
rect 10885 13481 10919 13515
rect 14197 13481 14231 13515
rect 15301 13481 15335 13515
rect 15393 13481 15427 13515
rect 17233 13481 17267 13515
rect 21557 13481 21591 13515
rect 15117 13413 15151 13447
rect 22385 13413 22419 13447
rect 4353 13345 4387 13379
rect 5181 13345 5215 13379
rect 6193 13345 6227 13379
rect 6285 13345 6319 13379
rect 7941 13345 7975 13379
rect 15761 13345 15795 13379
rect 18613 13345 18647 13379
rect 20913 13345 20947 13379
rect 22017 13345 22051 13379
rect 22109 13345 22143 13379
rect 22845 13345 22879 13379
rect 22937 13345 22971 13379
rect 3433 13277 3467 13311
rect 5089 13277 5123 13311
rect 6101 13277 6135 13311
rect 10526 13277 10560 13311
rect 10793 13277 10827 13311
rect 12265 13277 12299 13311
rect 13185 13277 13219 13311
rect 15669 13277 15703 13311
rect 18889 13277 18923 13311
rect 20637 13277 20671 13311
rect 4169 13209 4203 13243
rect 4997 13209 5031 13243
rect 7696 13209 7730 13243
rect 8401 13209 8435 13243
rect 9045 13209 9079 13243
rect 11998 13209 12032 13243
rect 16028 13209 16062 13243
rect 18346 13209 18380 13243
rect 18797 13209 18831 13243
rect 20392 13209 20426 13243
rect 21097 13209 21131 13243
rect 21925 13209 21959 13243
rect 3617 13141 3651 13175
rect 4261 13141 4295 13175
rect 5733 13141 5767 13175
rect 9413 13141 9447 13175
rect 12449 13141 12483 13175
rect 13829 13141 13863 13175
rect 17141 13141 17175 13175
rect 19073 13141 19107 13175
rect 19257 13141 19291 13175
rect 21005 13141 21039 13175
rect 21465 13141 21499 13175
rect 22753 13141 22787 13175
rect 3617 12937 3651 12971
rect 4077 12937 4111 12971
rect 4445 12937 4479 12971
rect 4813 12937 4847 12971
rect 5825 12937 5859 12971
rect 6837 12937 6871 12971
rect 10609 12937 10643 12971
rect 12633 12937 12667 12971
rect 13093 12937 13127 12971
rect 16221 12937 16255 12971
rect 16405 12937 16439 12971
rect 18337 12937 18371 12971
rect 20177 12937 20211 12971
rect 22201 12937 22235 12971
rect 22661 12937 22695 12971
rect 4905 12869 4939 12903
rect 7297 12869 7331 12903
rect 17794 12869 17828 12903
rect 18972 12869 19006 12903
rect 3985 12801 4019 12835
rect 6745 12801 6779 12835
rect 8502 12801 8536 12835
rect 8769 12801 8803 12835
rect 9974 12801 10008 12835
rect 10241 12801 10275 12835
rect 10701 12801 10735 12835
rect 12725 12801 12759 12835
rect 13185 12801 13219 12835
rect 13452 12801 13486 12835
rect 14657 12801 14691 12835
rect 14924 12801 14958 12835
rect 18153 12801 18187 12835
rect 18429 12801 18463 12835
rect 21290 12801 21324 12835
rect 21557 12801 21591 12835
rect 23121 12801 23155 12835
rect 4261 12733 4295 12767
rect 5089 12733 5123 12767
rect 5917 12733 5951 12767
rect 6101 12733 6135 12767
rect 6929 12733 6963 12767
rect 10517 12733 10551 12767
rect 12541 12733 12575 12767
rect 18061 12733 18095 12767
rect 18705 12733 18739 12767
rect 22293 12733 22327 12767
rect 22385 12733 22419 12767
rect 8861 12665 8895 12699
rect 11069 12665 11103 12699
rect 11253 12665 11287 12699
rect 16037 12665 16071 12699
rect 20085 12665 20119 12699
rect 5457 12597 5491 12631
rect 6377 12597 6411 12631
rect 7389 12597 7423 12631
rect 11621 12597 11655 12631
rect 14565 12597 14599 12631
rect 16681 12597 16715 12631
rect 18613 12597 18647 12631
rect 21833 12597 21867 12631
rect 22937 12597 22971 12631
rect 8493 12393 8527 12427
rect 10609 12393 10643 12427
rect 12173 12393 12207 12427
rect 13277 12393 13311 12427
rect 16589 12393 16623 12427
rect 21465 12393 21499 12427
rect 9689 12325 9723 12359
rect 14473 12325 14507 12359
rect 14657 12325 14691 12359
rect 16497 12325 16531 12359
rect 4445 12257 4479 12291
rect 4629 12257 4663 12291
rect 5457 12257 5491 12291
rect 9137 12257 9171 12291
rect 10333 12257 10367 12291
rect 11989 12257 12023 12291
rect 12725 12257 12759 12291
rect 17141 12257 17175 12291
rect 17601 12257 17635 12291
rect 20913 12257 20947 12291
rect 22201 12257 22235 12291
rect 23029 12257 23063 12291
rect 5181 12189 5215 12223
rect 7021 12189 7055 12223
rect 7113 12189 7147 12223
rect 9321 12189 9355 12223
rect 12909 12189 12943 12223
rect 15117 12189 15151 12223
rect 16957 12189 16991 12223
rect 18521 12189 18555 12223
rect 18613 12189 18647 12223
rect 18889 12189 18923 12223
rect 19257 12189 19291 12223
rect 21005 12189 21039 12223
rect 21925 12189 21959 12223
rect 22845 12189 22879 12223
rect 4353 12121 4387 12155
rect 6754 12121 6788 12155
rect 7358 12121 7392 12155
rect 8585 12121 8619 12155
rect 9229 12121 9263 12155
rect 10149 12121 10183 12155
rect 11722 12121 11756 12155
rect 15384 12121 15418 12155
rect 17785 12121 17819 12155
rect 19524 12121 19558 12155
rect 21097 12121 21131 12155
rect 3985 12053 4019 12087
rect 4813 12053 4847 12087
rect 5273 12053 5307 12087
rect 5641 12053 5675 12087
rect 9781 12053 9815 12087
rect 10241 12053 10275 12087
rect 12817 12053 12851 12087
rect 15025 12053 15059 12087
rect 17049 12053 17083 12087
rect 17693 12053 17727 12087
rect 18153 12053 18187 12087
rect 18337 12053 18371 12087
rect 18797 12053 18831 12087
rect 19073 12053 19107 12087
rect 20637 12053 20671 12087
rect 21557 12053 21591 12087
rect 22017 12053 22051 12087
rect 22385 12053 22419 12087
rect 22753 12053 22787 12087
rect 3341 11849 3375 11883
rect 3617 11849 3651 11883
rect 4445 11849 4479 11883
rect 4905 11849 4939 11883
rect 4997 11849 5031 11883
rect 5457 11849 5491 11883
rect 5825 11849 5859 11883
rect 6837 11849 6871 11883
rect 9689 11849 9723 11883
rect 12909 11849 12943 11883
rect 13921 11849 13955 11883
rect 14289 11849 14323 11883
rect 14933 11849 14967 11883
rect 15393 11849 15427 11883
rect 16037 11849 16071 11883
rect 16497 11849 16531 11883
rect 16957 11849 16991 11883
rect 17417 11849 17451 11883
rect 18337 11849 18371 11883
rect 20085 11849 20119 11883
rect 5917 11781 5951 11815
rect 7950 11781 7984 11815
rect 10824 11781 10858 11815
rect 14473 11781 14507 11815
rect 14565 11781 14599 11815
rect 14749 11781 14783 11815
rect 15301 11781 15335 11815
rect 17693 11781 17727 11815
rect 22201 11781 22235 11815
rect 22661 11781 22695 11815
rect 22845 11781 22879 11815
rect 3157 11713 3191 11747
rect 3433 11713 3467 11747
rect 3985 11713 4019 11747
rect 4077 11713 4111 11747
rect 11785 11713 11819 11747
rect 13369 11713 13403 11747
rect 16129 11713 16163 11747
rect 17049 11713 17083 11747
rect 17877 11713 17911 11747
rect 18153 11713 18187 11747
rect 18429 11713 18463 11747
rect 18705 11713 18739 11747
rect 18972 11713 19006 11747
rect 21290 11713 21324 11747
rect 21557 11713 21591 11747
rect 23029 11713 23063 11747
rect 3893 11645 3927 11679
rect 5089 11645 5123 11679
rect 6101 11645 6135 11679
rect 8217 11645 8251 11679
rect 11069 11645 11103 11679
rect 11253 11645 11287 11679
rect 11529 11645 11563 11679
rect 13461 11645 13495 11679
rect 13553 11645 13587 11679
rect 15485 11645 15519 11679
rect 15945 11645 15979 11679
rect 16865 11645 16899 11679
rect 22293 11645 22327 11679
rect 22385 11645 22419 11679
rect 4537 11577 4571 11611
rect 17509 11577 17543 11611
rect 8309 11509 8343 11543
rect 13001 11509 13035 11543
rect 18061 11509 18095 11543
rect 18613 11509 18647 11543
rect 20177 11509 20211 11543
rect 21833 11509 21867 11543
rect 7205 11305 7239 11339
rect 10425 11305 10459 11339
rect 11989 11305 12023 11339
rect 13553 11305 13587 11339
rect 13645 11305 13679 11339
rect 15669 11305 15703 11339
rect 19257 11305 19291 11339
rect 21465 11305 21499 11339
rect 5733 11237 5767 11271
rect 10333 11237 10367 11271
rect 15485 11237 15519 11271
rect 22293 11237 22327 11271
rect 4169 11169 4203 11203
rect 4813 11169 4847 11203
rect 13369 11169 13403 11203
rect 14105 11169 14139 11203
rect 17049 11169 17083 11203
rect 17693 11169 17727 11203
rect 20913 11169 20947 11203
rect 21741 11169 21775 11203
rect 22845 11169 22879 11203
rect 23029 11169 23063 11203
rect 5089 11101 5123 11135
rect 7113 11101 7147 11135
rect 8585 11101 8619 11135
rect 8677 11101 8711 11135
rect 8953 11101 8987 11135
rect 9220 11101 9254 11135
rect 11805 11101 11839 11135
rect 14372 11101 14406 11135
rect 17141 11101 17175 11135
rect 20370 11101 20404 11135
rect 20637 11101 20671 11135
rect 21097 11101 21131 11135
rect 22753 11101 22787 11135
rect 4261 11033 4295 11067
rect 6846 11033 6880 11067
rect 8318 11033 8352 11067
rect 11560 11033 11594 11067
rect 13102 11033 13136 11067
rect 13921 11033 13955 11067
rect 16782 11033 16816 11067
rect 17601 11033 17635 11067
rect 17960 11033 17994 11067
rect 21005 11033 21039 11067
rect 21925 11033 21959 11067
rect 4353 10965 4387 10999
rect 4721 10965 4755 10999
rect 17325 10965 17359 10999
rect 19073 10965 19107 10999
rect 21833 10965 21867 10999
rect 22385 10965 22419 10999
rect 4629 10761 4663 10795
rect 4997 10761 5031 10795
rect 5457 10761 5491 10795
rect 12909 10761 12943 10795
rect 13277 10761 13311 10795
rect 15025 10761 15059 10795
rect 22569 10761 22603 10795
rect 5089 10693 5123 10727
rect 5917 10693 5951 10727
rect 7950 10693 7984 10727
rect 9106 10693 9140 10727
rect 11796 10693 11830 10727
rect 14666 10693 14700 10727
rect 18245 10693 18279 10727
rect 21557 10693 21591 10727
rect 22109 10693 22143 10727
rect 23029 10693 23063 10727
rect 4537 10625 4571 10659
rect 5825 10625 5859 10659
rect 10517 10625 10551 10659
rect 10701 10625 10735 10659
rect 11529 10625 11563 10659
rect 13369 10625 13403 10659
rect 14933 10625 14967 10659
rect 16138 10625 16172 10659
rect 16405 10625 16439 10659
rect 16681 10625 16715 10659
rect 16948 10625 16982 10659
rect 18337 10625 18371 10659
rect 18613 10625 18647 10659
rect 18880 10625 18914 10659
rect 20352 10625 20386 10659
rect 22201 10625 22235 10659
rect 22845 10625 22879 10659
rect 5181 10557 5215 10591
rect 6009 10557 6043 10591
rect 8217 10557 8251 10591
rect 8861 10557 8895 10591
rect 13093 10557 13127 10591
rect 20085 10557 20119 10591
rect 21925 10557 21959 10591
rect 22661 10557 22695 10591
rect 4353 10489 4387 10523
rect 6837 10489 6871 10523
rect 10241 10489 10275 10523
rect 18061 10489 18095 10523
rect 6653 10421 6687 10455
rect 8309 10421 8343 10455
rect 13553 10421 13587 10455
rect 18521 10421 18555 10455
rect 19993 10421 20027 10455
rect 21465 10421 21499 10455
rect 3617 10217 3651 10251
rect 4537 10217 4571 10251
rect 7297 10217 7331 10251
rect 10517 10217 10551 10251
rect 10609 10217 10643 10251
rect 12909 10217 12943 10251
rect 13829 10149 13863 10183
rect 15485 10149 15519 10183
rect 15669 10149 15703 10183
rect 15761 10149 15795 10183
rect 15945 10149 15979 10183
rect 20729 10149 20763 10183
rect 3985 10081 4019 10115
rect 5641 10081 5675 10115
rect 5917 10081 5951 10115
rect 11713 10081 11747 10115
rect 13553 10081 13587 10115
rect 16589 10081 16623 10115
rect 18797 10081 18831 10115
rect 22753 10081 22787 10115
rect 3433 10013 3467 10047
rect 4905 10013 4939 10047
rect 5549 10013 5583 10047
rect 8769 10013 8803 10047
rect 10333 10013 10367 10047
rect 11989 10013 12023 10047
rect 14105 10013 14139 10047
rect 14361 10013 14395 10047
rect 16773 10013 16807 10047
rect 18429 10013 18463 10047
rect 19073 10013 19107 10047
rect 19257 10013 19291 10047
rect 19524 10013 19558 10047
rect 21842 10013 21876 10047
rect 22109 10013 22143 10047
rect 22661 10013 22695 10047
rect 4169 9945 4203 9979
rect 4721 9945 4755 9979
rect 6184 9945 6218 9979
rect 8502 9945 8536 9979
rect 10066 9945 10100 9979
rect 11897 9945 11931 9979
rect 12725 9945 12759 9979
rect 18184 9945 18218 9979
rect 23029 9945 23063 9979
rect 4077 9877 4111 9911
rect 5089 9877 5123 9911
rect 5457 9877 5491 9911
rect 7389 9877 7423 9911
rect 8953 9877 8987 9911
rect 12357 9877 12391 9911
rect 13001 9877 13035 9911
rect 13369 9877 13403 9911
rect 13461 9877 13495 9911
rect 16957 9877 16991 9911
rect 17049 9877 17083 9911
rect 20637 9877 20671 9911
rect 22201 9877 22235 9911
rect 22569 9877 22603 9911
rect 3525 9673 3559 9707
rect 3801 9673 3835 9707
rect 6837 9673 6871 9707
rect 9873 9673 9907 9707
rect 11713 9673 11747 9707
rect 13277 9673 13311 9707
rect 13461 9673 13495 9707
rect 16405 9673 16439 9707
rect 16681 9673 16715 9707
rect 5089 9605 5123 9639
rect 9422 9605 9456 9639
rect 11621 9605 11655 9639
rect 22845 9605 22879 9639
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 3341 9537 3375 9571
rect 3617 9537 3651 9571
rect 4261 9537 4295 9571
rect 4353 9537 4387 9571
rect 5181 9537 5215 9571
rect 7950 9537 7984 9571
rect 9689 9537 9723 9571
rect 10609 9537 10643 9571
rect 11253 9537 11287 9571
rect 12837 9537 12871 9571
rect 13093 9537 13127 9571
rect 14574 9537 14608 9571
rect 14841 9537 14875 9571
rect 14933 9537 14967 9571
rect 15200 9537 15234 9571
rect 16865 9537 16899 9571
rect 17141 9537 17175 9571
rect 18541 9537 18575 9571
rect 18797 9537 18831 9571
rect 20002 9537 20036 9571
rect 20361 9537 20395 9571
rect 21465 9537 21499 9571
rect 22201 9537 22235 9571
rect 4445 9469 4479 9503
rect 5365 9469 5399 9503
rect 8217 9469 8251 9503
rect 10701 9469 10735 9503
rect 10885 9469 10919 9503
rect 20269 9469 20303 9503
rect 20729 9469 20763 9503
rect 21925 9469 21959 9503
rect 22109 9469 22143 9503
rect 22661 9469 22695 9503
rect 8309 9401 8343 9435
rect 16313 9401 16347 9435
rect 17049 9401 17083 9435
rect 21649 9401 21683 9435
rect 1593 9333 1627 9367
rect 3893 9333 3927 9367
rect 4721 9333 4755 9367
rect 6653 9333 6687 9367
rect 10241 9333 10275 9367
rect 11161 9333 11195 9367
rect 17325 9333 17359 9367
rect 17417 9333 17451 9367
rect 18889 9333 18923 9367
rect 22569 9333 22603 9367
rect 23029 9333 23063 9367
rect 3617 9129 3651 9163
rect 6285 9129 6319 9163
rect 12909 9129 12943 9163
rect 13829 9129 13863 9163
rect 14197 9129 14231 9163
rect 14381 9129 14415 9163
rect 15945 9129 15979 9163
rect 3985 9061 4019 9095
rect 19073 9061 19107 9095
rect 22201 9061 22235 9095
rect 2973 8993 3007 9027
rect 3157 8993 3191 9027
rect 4445 8993 4479 9027
rect 4629 8993 4663 9027
rect 5273 8993 5307 9027
rect 5365 8993 5399 9027
rect 12817 8993 12851 9027
rect 13553 8993 13587 9027
rect 14565 8993 14599 9027
rect 22661 8993 22695 9027
rect 22753 8993 22787 9027
rect 4353 8925 4387 8959
rect 5181 8925 5215 8959
rect 7665 8925 7699 8959
rect 8401 8925 8435 8959
rect 8585 8925 8619 8959
rect 9965 8925 9999 8959
rect 10232 8925 10266 8959
rect 13369 8925 13403 8959
rect 14832 8925 14866 8959
rect 17417 8925 17451 8959
rect 17509 8925 17543 8959
rect 20370 8925 20404 8959
rect 20637 8925 20671 8959
rect 22109 8925 22143 8959
rect 7398 8857 7432 8891
rect 12572 8857 12606 8891
rect 13277 8857 13311 8891
rect 17172 8857 17206 8891
rect 17776 8857 17810 8891
rect 21842 8857 21876 8891
rect 22569 8857 22603 8891
rect 3249 8789 3283 8823
rect 4813 8789 4847 8823
rect 7849 8789 7883 8823
rect 11345 8789 11379 8823
rect 11437 8789 11471 8823
rect 16037 8789 16071 8823
rect 18889 8789 18923 8823
rect 19257 8789 19291 8823
rect 20729 8789 20763 8823
rect 23029 8789 23063 8823
rect 3525 8585 3559 8619
rect 6193 8585 6227 8619
rect 8309 8585 8343 8619
rect 9965 8585 9999 8619
rect 16313 8585 16347 8619
rect 18061 8585 18095 8619
rect 19533 8585 19567 8619
rect 3157 8517 3191 8551
rect 3985 8517 4019 8551
rect 9873 8517 9907 8551
rect 16937 8517 16971 8551
rect 22845 8517 22879 8551
rect 4813 8449 4847 8483
rect 5069 8449 5103 8483
rect 7104 8449 7138 8483
rect 9422 8449 9456 8483
rect 9689 8449 9723 8483
rect 11078 8449 11112 8483
rect 11345 8449 11379 8483
rect 12642 8449 12676 8483
rect 14832 8449 14866 8483
rect 18420 8449 18454 8483
rect 19881 8449 19915 8483
rect 21189 8449 21223 8483
rect 21373 8449 21407 8483
rect 22201 8449 22235 8483
rect 23121 8449 23155 8483
rect 2973 8381 3007 8415
rect 3065 8381 3099 8415
rect 4077 8381 4111 8415
rect 4169 8381 4203 8415
rect 6837 8381 6871 8415
rect 12909 8381 12943 8415
rect 14565 8381 14599 8415
rect 16681 8381 16715 8415
rect 18153 8381 18187 8415
rect 19625 8381 19659 8415
rect 22293 8381 22327 8415
rect 22385 8381 22419 8415
rect 3617 8313 3651 8347
rect 8217 8313 8251 8347
rect 11529 8313 11563 8347
rect 15945 8313 15979 8347
rect 16129 8313 16163 8347
rect 16405 8313 16439 8347
rect 21557 8313 21591 8347
rect 21833 8313 21867 8347
rect 6469 8245 6503 8279
rect 13093 8245 13127 8279
rect 13369 8245 13403 8279
rect 13553 8245 13587 8279
rect 13737 8245 13771 8279
rect 13921 8245 13955 8279
rect 14105 8245 14139 8279
rect 14289 8245 14323 8279
rect 14473 8245 14507 8279
rect 21005 8245 21039 8279
rect 7389 8041 7423 8075
rect 18797 7973 18831 8007
rect 9781 7905 9815 7939
rect 11805 7905 11839 7939
rect 21281 7905 21315 7939
rect 21744 7905 21778 7939
rect 4445 7837 4479 7871
rect 7297 7837 7331 7871
rect 8769 7837 8803 7871
rect 10048 7837 10082 7871
rect 12173 7837 12207 7871
rect 12357 7837 12391 7871
rect 12541 7837 12575 7871
rect 14105 7837 14139 7871
rect 15577 7837 15611 7871
rect 18173 7837 18207 7871
rect 18429 7837 18463 7871
rect 18613 7837 18647 7871
rect 19073 7837 19107 7871
rect 20637 7837 20671 7871
rect 21604 7837 21638 7871
rect 22017 7837 22051 7871
rect 4712 7769 4746 7803
rect 7052 7769 7086 7803
rect 8502 7769 8536 7803
rect 11713 7769 11747 7803
rect 12808 7769 12842 7803
rect 14350 7769 14384 7803
rect 15844 7769 15878 7803
rect 20370 7769 20404 7803
rect 20913 7769 20947 7803
rect 21097 7769 21131 7803
rect 5825 7701 5859 7735
rect 5917 7701 5951 7735
rect 8953 7701 8987 7735
rect 9137 7701 9171 7735
rect 9597 7701 9631 7735
rect 11161 7701 11195 7735
rect 11253 7701 11287 7735
rect 11621 7701 11655 7735
rect 13921 7701 13955 7735
rect 15485 7701 15519 7735
rect 16957 7701 16991 7735
rect 17049 7701 17083 7735
rect 19257 7701 19291 7735
rect 20729 7701 20763 7735
rect 23121 7701 23155 7735
rect 3985 7497 4019 7531
rect 4353 7497 4387 7531
rect 6193 7497 6227 7531
rect 11345 7497 11379 7531
rect 13093 7497 13127 7531
rect 18061 7497 18095 7531
rect 21465 7497 21499 7531
rect 22109 7497 22143 7531
rect 22569 7497 22603 7531
rect 6469 7429 6503 7463
rect 6653 7429 6687 7463
rect 6837 7429 6871 7463
rect 14298 7429 14332 7463
rect 19266 7429 19300 7463
rect 19870 7429 19904 7463
rect 21281 7429 21315 7463
rect 22845 7429 22879 7463
rect 4445 7361 4479 7395
rect 4813 7361 4847 7395
rect 5080 7361 5114 7395
rect 6929 7361 6963 7395
rect 7185 7361 7219 7395
rect 8493 7361 8527 7395
rect 8760 7361 8794 7395
rect 9965 7361 9999 7395
rect 10232 7361 10266 7395
rect 11621 7361 11655 7395
rect 11713 7361 11747 7395
rect 11980 7361 12014 7395
rect 15781 7361 15815 7395
rect 16948 7361 16982 7395
rect 21649 7361 21683 7395
rect 22201 7361 22235 7395
rect 4537 7293 4571 7327
rect 14565 7293 14599 7327
rect 16037 7293 16071 7327
rect 16681 7293 16715 7327
rect 19533 7293 19567 7327
rect 19625 7293 19659 7327
rect 21925 7293 21959 7327
rect 18153 7225 18187 7259
rect 22661 7225 22695 7259
rect 8309 7157 8343 7191
rect 9873 7157 9907 7191
rect 13185 7157 13219 7191
rect 14657 7157 14691 7191
rect 16221 7157 16255 7191
rect 16405 7157 16439 7191
rect 21005 7157 21039 7191
rect 23029 7157 23063 7191
rect 5641 6953 5675 6987
rect 8493 6953 8527 6987
rect 12173 6953 12207 6987
rect 13829 6953 13863 6987
rect 14197 6953 14231 6987
rect 14381 6953 14415 6987
rect 14749 6953 14783 6987
rect 19073 6885 19107 6919
rect 20637 6885 20671 6919
rect 12265 6817 12299 6851
rect 18521 6817 18555 6851
rect 21189 6817 21223 6851
rect 21652 6817 21686 6851
rect 21925 6817 21959 6851
rect 1961 6749 1995 6783
rect 7021 6749 7055 6783
rect 7113 6749 7147 6783
rect 8677 6749 8711 6783
rect 9045 6749 9079 6783
rect 9321 6749 9355 6783
rect 10793 6749 10827 6783
rect 15954 6749 15988 6783
rect 16221 6749 16255 6783
rect 17693 6749 17727 6783
rect 17969 6749 18003 6783
rect 19257 6749 19291 6783
rect 20913 6749 20947 6783
rect 6754 6681 6788 6715
rect 7358 6681 7392 6715
rect 9588 6681 9622 6715
rect 11060 6681 11094 6715
rect 12510 6681 12544 6715
rect 17426 6681 17460 6715
rect 18613 6681 18647 6715
rect 19524 6681 19558 6715
rect 20729 6681 20763 6715
rect 2145 6613 2179 6647
rect 10701 6613 10735 6647
rect 13645 6613 13679 6647
rect 14473 6613 14507 6647
rect 14841 6613 14875 6647
rect 16313 6613 16347 6647
rect 17785 6613 17819 6647
rect 18153 6613 18187 6647
rect 18705 6613 18739 6647
rect 21097 6613 21131 6647
rect 21655 6613 21689 6647
rect 23029 6613 23063 6647
rect 8401 6409 8435 6443
rect 8861 6409 8895 6443
rect 10517 6409 10551 6443
rect 13737 6409 13771 6443
rect 13921 6409 13955 6443
rect 14473 6409 14507 6443
rect 20913 6409 20947 6443
rect 21281 6409 21315 6443
rect 22753 6409 22787 6443
rect 7674 6341 7708 6375
rect 8953 6341 8987 6375
rect 9781 6341 9815 6375
rect 10609 6341 10643 6375
rect 13286 6341 13320 6375
rect 15577 6341 15611 6375
rect 20116 6341 20150 6375
rect 22201 6341 22235 6375
rect 22293 6341 22327 6375
rect 7941 6273 7975 6307
rect 8217 6273 8251 6307
rect 9689 6273 9723 6307
rect 11161 6273 11195 6307
rect 11529 6273 11563 6307
rect 11989 6273 12023 6307
rect 13553 6273 13587 6307
rect 14381 6273 14415 6307
rect 15025 6273 15059 6307
rect 15485 6273 15519 6307
rect 15945 6273 15979 6307
rect 16221 6273 16255 6307
rect 16773 6273 16807 6307
rect 17509 6273 17543 6307
rect 17776 6273 17810 6307
rect 20637 6273 20671 6307
rect 22845 6273 22879 6307
rect 9137 6205 9171 6239
rect 9965 6205 9999 6239
rect 10793 6205 10827 6239
rect 14565 6205 14599 6239
rect 15669 6205 15703 6239
rect 17141 6205 17175 6239
rect 17417 6205 17451 6239
rect 20361 6205 20395 6239
rect 21373 6205 21407 6239
rect 21465 6205 21499 6239
rect 22385 6205 22419 6239
rect 10149 6137 10183 6171
rect 11713 6137 11747 6171
rect 15117 6137 15151 6171
rect 20821 6137 20855 6171
rect 23029 6137 23063 6171
rect 6561 6069 6595 6103
rect 8033 6069 8067 6103
rect 8493 6069 8527 6103
rect 9321 6069 9355 6103
rect 11069 6069 11103 6103
rect 11805 6069 11839 6103
rect 12173 6069 12207 6103
rect 14013 6069 14047 6103
rect 14841 6069 14875 6103
rect 16405 6069 16439 6103
rect 18889 6069 18923 6103
rect 18981 6069 19015 6103
rect 20453 6069 20487 6103
rect 21833 6069 21867 6103
rect 7481 5865 7515 5899
rect 11621 5865 11655 5899
rect 11897 5865 11931 5899
rect 12357 5865 12391 5899
rect 23029 5865 23063 5899
rect 9045 5797 9079 5831
rect 9965 5797 9999 5831
rect 10977 5797 11011 5831
rect 11437 5797 11471 5831
rect 13921 5797 13955 5831
rect 19073 5797 19107 5831
rect 20637 5797 20671 5831
rect 5181 5729 5215 5763
rect 5365 5729 5399 5763
rect 5917 5729 5951 5763
rect 8401 5729 8435 5763
rect 9505 5729 9539 5763
rect 9689 5729 9723 5763
rect 10885 5729 10919 5763
rect 13277 5729 13311 5763
rect 13461 5729 13495 5763
rect 14105 5729 14139 5763
rect 14568 5727 14602 5761
rect 14841 5729 14875 5763
rect 16129 5729 16163 5763
rect 17696 5729 17730 5763
rect 19809 5729 19843 5763
rect 22014 5729 22048 5763
rect 22477 5729 22511 5763
rect 5457 5661 5491 5695
rect 6184 5661 6218 5695
rect 8125 5661 8159 5695
rect 9413 5661 9447 5695
rect 11253 5661 11287 5695
rect 11805 5661 11839 5695
rect 16405 5661 16439 5695
rect 17233 5661 17267 5695
rect 17969 5661 18003 5695
rect 19625 5661 19659 5695
rect 20085 5661 20119 5695
rect 21741 5661 21775 5695
rect 22753 5661 22787 5695
rect 22845 5661 22879 5695
rect 8217 5593 8251 5627
rect 16957 5593 16991 5627
rect 20361 5593 20395 5627
rect 5825 5525 5859 5559
rect 7297 5525 7331 5559
rect 7757 5525 7791 5559
rect 13553 5525 13587 5559
rect 14571 5525 14605 5559
rect 15945 5525 15979 5559
rect 16313 5525 16347 5559
rect 16773 5525 16807 5559
rect 17049 5525 17083 5559
rect 17699 5525 17733 5559
rect 19257 5525 19291 5559
rect 19717 5525 19751 5559
rect 20269 5525 20303 5559
rect 22010 5525 22044 5559
rect 22569 5525 22603 5559
rect 5825 5321 5859 5355
rect 6745 5321 6779 5355
rect 7113 5321 7147 5355
rect 7205 5321 7239 5355
rect 8585 5321 8619 5355
rect 10977 5321 11011 5355
rect 13553 5321 13587 5355
rect 14013 5321 14047 5355
rect 15031 5321 15065 5355
rect 16681 5321 16715 5355
rect 17509 5321 17543 5355
rect 17969 5321 18003 5355
rect 20637 5321 20671 5355
rect 21005 5321 21039 5355
rect 21925 5321 21959 5355
rect 22293 5321 22327 5355
rect 22385 5321 22419 5355
rect 22937 5321 22971 5355
rect 5733 5253 5767 5287
rect 8125 5253 8159 5287
rect 13921 5253 13955 5287
rect 14197 5253 14231 5287
rect 14381 5253 14415 5287
rect 20545 5253 20579 5287
rect 6561 5185 6595 5219
rect 8033 5185 8067 5219
rect 9965 5185 9999 5219
rect 10701 5185 10735 5219
rect 15301 5185 15335 5219
rect 17049 5185 17083 5219
rect 17141 5185 17175 5219
rect 17877 5185 17911 5219
rect 18337 5185 18371 5219
rect 19829 5185 19863 5219
rect 21557 5185 21591 5219
rect 22753 5185 22787 5219
rect 5641 5117 5675 5151
rect 6929 5117 6963 5151
rect 8309 5117 8343 5151
rect 10241 5117 10275 5151
rect 14565 5117 14599 5151
rect 15071 5117 15105 5151
rect 17233 5117 17267 5151
rect 18061 5117 18095 5151
rect 20085 5117 20119 5151
rect 20729 5117 20763 5151
rect 22477 5117 22511 5151
rect 7573 5049 7607 5083
rect 10885 5049 10919 5083
rect 6193 4981 6227 5015
rect 7665 4981 7699 5015
rect 8769 4981 8803 5015
rect 16405 4981 16439 5015
rect 18705 4981 18739 5015
rect 20177 4981 20211 5015
rect 7113 4777 7147 4811
rect 17417 4777 17451 4811
rect 19257 4777 19291 4811
rect 21281 4777 21315 4811
rect 7205 4709 7239 4743
rect 8401 4709 8435 4743
rect 6561 4641 6595 4675
rect 6653 4641 6687 4675
rect 8033 4641 8067 4675
rect 8217 4641 8251 4675
rect 9781 4641 9815 4675
rect 9965 4641 9999 4675
rect 15577 4641 15611 4675
rect 16056 4641 16090 4675
rect 16313 4641 16347 4675
rect 18153 4641 18187 4675
rect 18889 4641 18923 4675
rect 21741 4641 21775 4675
rect 21925 4641 21959 4675
rect 22661 4641 22695 4675
rect 6101 4573 6135 4607
rect 7389 4573 7423 4607
rect 7941 4573 7975 4607
rect 10057 4573 10091 4607
rect 17877 4573 17911 4607
rect 20637 4573 20671 4607
rect 20913 4573 20947 4607
rect 21189 4573 21223 4607
rect 22477 4573 22511 4607
rect 22569 4573 22603 4607
rect 6745 4505 6779 4539
rect 18797 4505 18831 4539
rect 20370 4505 20404 4539
rect 21649 4505 21683 4539
rect 22937 4505 22971 4539
rect 6285 4437 6319 4471
rect 7573 4437 7607 4471
rect 10425 4437 10459 4471
rect 16043 4437 16077 4471
rect 17509 4437 17543 4471
rect 17969 4437 18003 4471
rect 18337 4437 18371 4471
rect 18705 4437 18739 4471
rect 20729 4437 20763 4471
rect 21005 4437 21039 4471
rect 22109 4437 22143 4471
rect 7205 4233 7239 4267
rect 17877 4233 17911 4267
rect 19165 4233 19199 4267
rect 19809 4233 19843 4267
rect 20729 4233 20763 4267
rect 22109 4233 22143 4267
rect 16129 4165 16163 4199
rect 16497 4165 16531 4199
rect 17049 4165 17083 4199
rect 22201 4165 22235 4199
rect 10425 4097 10459 4131
rect 10885 4097 10919 4131
rect 15945 4097 15979 4131
rect 16957 4097 16991 4131
rect 17785 4097 17819 4131
rect 18705 4097 18739 4131
rect 19349 4097 19383 4131
rect 19717 4097 19751 4131
rect 20637 4097 20671 4131
rect 21281 4097 21315 4131
rect 21373 4097 21407 4131
rect 22845 4097 22879 4131
rect 16773 4029 16807 4063
rect 17601 4029 17635 4063
rect 18429 4029 18463 4063
rect 18613 4029 18647 4063
rect 19533 4029 19567 4063
rect 20913 4029 20947 4063
rect 22017 4029 22051 4063
rect 20177 3961 20211 3995
rect 21097 3961 21131 3995
rect 23029 3961 23063 3995
rect 10609 3893 10643 3927
rect 11069 3893 11103 3927
rect 17417 3893 17451 3927
rect 18245 3893 18279 3927
rect 19073 3893 19107 3927
rect 20269 3893 20303 3927
rect 21557 3893 21591 3927
rect 22569 3893 22603 3927
rect 22661 3893 22695 3927
rect 17233 3689 17267 3723
rect 19349 3689 19383 3723
rect 19625 3689 19659 3723
rect 20637 3689 20671 3723
rect 22569 3689 22603 3723
rect 23029 3689 23063 3723
rect 12357 3553 12391 3587
rect 12541 3553 12575 3587
rect 15856 3553 15890 3587
rect 16129 3553 16163 3587
rect 17877 3553 17911 3587
rect 18061 3553 18095 3587
rect 19993 3553 20027 3587
rect 21465 3553 21499 3587
rect 22293 3553 22327 3587
rect 1593 3485 1627 3519
rect 12633 3485 12667 3519
rect 15393 3485 15427 3519
rect 17601 3485 17635 3519
rect 18981 3485 19015 3519
rect 19533 3485 19567 3519
rect 19809 3485 19843 3519
rect 20729 3485 20763 3519
rect 21281 3485 21315 3519
rect 22201 3485 22235 3519
rect 22753 3485 22787 3519
rect 22845 3485 22879 3519
rect 18153 3417 18187 3451
rect 18613 3417 18647 3451
rect 1409 3349 1443 3383
rect 13001 3349 13035 3383
rect 15859 3349 15893 3383
rect 17325 3349 17359 3383
rect 18521 3349 18555 3383
rect 20177 3349 20211 3383
rect 20269 3349 20303 3383
rect 20913 3349 20947 3383
rect 21373 3349 21407 3383
rect 21741 3349 21775 3383
rect 22109 3349 22143 3383
rect 16957 3145 16991 3179
rect 17049 3145 17083 3179
rect 17417 3145 17451 3179
rect 18337 3145 18371 3179
rect 18797 3145 18831 3179
rect 21373 3145 21407 3179
rect 23029 3145 23063 3179
rect 17877 3077 17911 3111
rect 19809 3077 19843 3111
rect 20545 3077 20579 3111
rect 21833 3077 21867 3111
rect 6561 3009 6595 3043
rect 18153 3009 18187 3043
rect 19257 3009 19291 3043
rect 20637 3009 20671 3043
rect 21281 3009 21315 3043
rect 22661 3009 22695 3043
rect 22845 3009 22879 3043
rect 16773 2941 16807 2975
rect 19073 2941 19107 2975
rect 19717 2941 19751 2975
rect 20085 2941 20119 2975
rect 20729 2941 20763 2975
rect 22385 2941 22419 2975
rect 19533 2873 19567 2907
rect 6377 2805 6411 2839
rect 6745 2805 6779 2839
rect 20177 2805 20211 2839
rect 21097 2805 21131 2839
rect 19349 2601 19383 2635
rect 20177 2601 20211 2635
rect 20361 2601 20395 2635
rect 20545 2601 20579 2635
rect 23029 2601 23063 2635
rect 19809 2533 19843 2567
rect 20729 2533 20763 2567
rect 20913 2533 20947 2567
rect 21097 2533 21131 2567
rect 21557 2533 21591 2567
rect 19533 2465 19567 2499
rect 22109 2465 22143 2499
rect 2513 2397 2547 2431
rect 6377 2397 6411 2431
rect 10609 2397 10643 2431
rect 10793 2397 10827 2431
rect 20085 2397 20119 2431
rect 21373 2397 21407 2431
rect 22201 2397 22235 2431
rect 22477 2397 22511 2431
rect 22845 2397 22879 2431
rect 2329 2261 2363 2295
rect 10425 2261 10459 2295
rect 19625 2261 19659 2295
rect 22385 2261 22419 2295
rect 22661 2261 22695 2295
<< metal1 >>
rect 4062 22720 4068 22772
rect 4120 22760 4126 22772
rect 5442 22760 5448 22772
rect 4120 22732 5448 22760
rect 4120 22720 4126 22732
rect 5442 22720 5448 22732
rect 5500 22720 5506 22772
rect 6178 22720 6184 22772
rect 6236 22760 6242 22772
rect 9306 22760 9312 22772
rect 6236 22732 9312 22760
rect 6236 22720 6242 22732
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 11422 22720 11428 22772
rect 11480 22760 11486 22772
rect 11882 22760 11888 22772
rect 11480 22732 11888 22760
rect 11480 22720 11486 22732
rect 11882 22720 11888 22732
rect 11940 22720 11946 22772
rect 3602 22652 3608 22704
rect 3660 22692 3666 22704
rect 12158 22692 12164 22704
rect 3660 22664 12164 22692
rect 3660 22652 3666 22664
rect 12158 22652 12164 22664
rect 12216 22652 12222 22704
rect 4982 22584 4988 22636
rect 5040 22624 5046 22636
rect 14366 22624 14372 22636
rect 5040 22596 14372 22624
rect 5040 22584 5046 22596
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 19610 22584 19616 22636
rect 19668 22624 19674 22636
rect 22002 22624 22008 22636
rect 19668 22596 22008 22624
rect 19668 22584 19674 22596
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 4614 22516 4620 22568
rect 4672 22556 4678 22568
rect 6730 22556 6736 22568
rect 4672 22528 6736 22556
rect 4672 22516 4678 22528
rect 6730 22516 6736 22528
rect 6788 22516 6794 22568
rect 7190 22516 7196 22568
rect 7248 22556 7254 22568
rect 7248 22528 19334 22556
rect 7248 22516 7254 22528
rect 5534 22448 5540 22500
rect 5592 22488 5598 22500
rect 8662 22488 8668 22500
rect 5592 22460 8668 22488
rect 5592 22448 5598 22460
rect 8662 22448 8668 22460
rect 8720 22448 8726 22500
rect 10870 22448 10876 22500
rect 10928 22488 10934 22500
rect 11514 22488 11520 22500
rect 10928 22460 11520 22488
rect 10928 22448 10934 22460
rect 11514 22448 11520 22460
rect 11572 22488 11578 22500
rect 12526 22488 12532 22500
rect 11572 22460 12532 22488
rect 11572 22448 11578 22460
rect 12526 22448 12532 22460
rect 12584 22448 12590 22500
rect 12710 22448 12716 22500
rect 12768 22488 12774 22500
rect 18322 22488 18328 22500
rect 12768 22460 18328 22488
rect 12768 22448 12774 22460
rect 18322 22448 18328 22460
rect 18380 22448 18386 22500
rect 19306 22488 19334 22528
rect 21450 22488 21456 22500
rect 19306 22460 21456 22488
rect 21450 22448 21456 22460
rect 21508 22448 21514 22500
rect 5442 22380 5448 22432
rect 5500 22420 5506 22432
rect 8018 22420 8024 22432
rect 5500 22392 8024 22420
rect 5500 22380 5506 22392
rect 8018 22380 8024 22392
rect 8076 22380 8082 22432
rect 12158 22380 12164 22432
rect 12216 22420 12222 22432
rect 13998 22420 14004 22432
rect 12216 22392 14004 22420
rect 12216 22380 12222 22392
rect 13998 22380 14004 22392
rect 14056 22380 14062 22432
rect 14090 22380 14096 22432
rect 14148 22420 14154 22432
rect 18138 22420 18144 22432
rect 14148 22392 18144 22420
rect 14148 22380 14154 22392
rect 18138 22380 18144 22392
rect 18196 22380 18202 22432
rect 1104 22330 23460 22352
rect 1104 22278 3749 22330
rect 3801 22278 3813 22330
rect 3865 22278 3877 22330
rect 3929 22278 3941 22330
rect 3993 22278 4005 22330
rect 4057 22278 9347 22330
rect 9399 22278 9411 22330
rect 9463 22278 9475 22330
rect 9527 22278 9539 22330
rect 9591 22278 9603 22330
rect 9655 22278 14945 22330
rect 14997 22278 15009 22330
rect 15061 22278 15073 22330
rect 15125 22278 15137 22330
rect 15189 22278 15201 22330
rect 15253 22278 20543 22330
rect 20595 22278 20607 22330
rect 20659 22278 20671 22330
rect 20723 22278 20735 22330
rect 20787 22278 20799 22330
rect 20851 22278 23460 22330
rect 1104 22256 23460 22278
rect 5350 22216 5356 22228
rect 5311 22188 5356 22216
rect 5350 22176 5356 22188
rect 5408 22176 5414 22228
rect 10962 22216 10968 22228
rect 9646 22188 10968 22216
rect 5166 22148 5172 22160
rect 2792 22120 5172 22148
rect 1581 22083 1639 22089
rect 1581 22049 1593 22083
rect 1627 22080 1639 22083
rect 2314 22080 2320 22092
rect 1627 22052 2320 22080
rect 1627 22049 1639 22052
rect 1581 22043 1639 22049
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 2792 22080 2820 22120
rect 5166 22108 5172 22120
rect 5224 22108 5230 22160
rect 5258 22108 5264 22160
rect 5316 22148 5322 22160
rect 9030 22148 9036 22160
rect 5316 22120 6316 22148
rect 5316 22108 5322 22120
rect 2424 22052 2820 22080
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 21981 2007 22015
rect 1949 21975 2007 21981
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 22012 2283 22015
rect 2424 22012 2452 22052
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 6288 22080 6316 22120
rect 8588 22120 9036 22148
rect 8588 22089 8616 22120
rect 9030 22108 9036 22120
rect 9088 22108 9094 22160
rect 7285 22083 7343 22089
rect 7285 22080 7297 22083
rect 3200 22052 6132 22080
rect 6288 22052 7297 22080
rect 3200 22040 3206 22052
rect 2590 22012 2596 22024
rect 2271 21984 2452 22012
rect 2551 21984 2596 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 1964 21944 1992 21975
rect 2590 21972 2596 21984
rect 2648 21972 2654 22024
rect 2869 22015 2927 22021
rect 2869 21981 2881 22015
rect 2915 22012 2927 22015
rect 3050 22012 3056 22024
rect 2915 21984 3056 22012
rect 2915 21981 2927 21984
rect 2869 21975 2927 21981
rect 3050 21972 3056 21984
rect 3108 21972 3114 22024
rect 3234 22012 3240 22024
rect 3195 21984 3240 22012
rect 3234 21972 3240 21984
rect 3292 21972 3298 22024
rect 3602 22012 3608 22024
rect 3563 21984 3608 22012
rect 3602 21972 3608 21984
rect 3660 21972 3666 22024
rect 4062 22021 4068 22024
rect 4058 21975 4068 22021
rect 4120 22012 4126 22024
rect 4249 22015 4307 22021
rect 4120 21984 4158 22012
rect 4062 21972 4068 21975
rect 4120 21972 4126 21984
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4338 22012 4344 22024
rect 4295 21984 4344 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 4338 21972 4344 21984
rect 4396 21972 4402 22024
rect 4614 22012 4620 22024
rect 4575 21984 4620 22012
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 4798 21972 4804 22024
rect 4856 22012 4862 22024
rect 4893 22015 4951 22021
rect 4893 22012 4905 22015
rect 4856 21984 4905 22012
rect 4856 21972 4862 21984
rect 4893 21981 4905 21984
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 5166 21972 5172 22024
rect 5224 22012 5230 22024
rect 5442 22012 5448 22024
rect 5224 21984 5448 22012
rect 5224 21972 5230 21984
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 5718 22012 5724 22024
rect 5679 21984 5724 22012
rect 5718 21972 5724 21984
rect 5776 21972 5782 22024
rect 6104 22008 6132 22052
rect 7285 22049 7297 22052
rect 7331 22049 7343 22083
rect 7285 22043 7343 22049
rect 8573 22083 8631 22089
rect 8573 22049 8585 22083
rect 8619 22080 8631 22083
rect 8619 22052 8653 22080
rect 8619 22049 8631 22052
rect 8573 22043 8631 22049
rect 8754 22040 8760 22092
rect 8812 22080 8818 22092
rect 9493 22083 9551 22089
rect 8812 22052 9352 22080
rect 8812 22040 8818 22052
rect 6178 22021 6184 22024
rect 6173 22008 6184 22021
rect 6104 21980 6184 22008
rect 6236 22012 6242 22024
rect 6236 21984 6273 22012
rect 6173 21975 6184 21980
rect 6178 21972 6184 21975
rect 6236 21972 6242 21984
rect 6362 21972 6368 22024
rect 6420 22012 6426 22024
rect 6730 22012 6736 22024
rect 6420 21984 6736 22012
rect 6420 21972 6426 21984
rect 6730 21972 6736 21984
rect 6788 21972 6794 22024
rect 7392 21984 8156 22012
rect 7392 21956 7420 21984
rect 2682 21944 2688 21956
rect 1964 21916 2688 21944
rect 2682 21904 2688 21916
rect 2740 21904 2746 21956
rect 7009 21947 7067 21953
rect 7009 21944 7021 21947
rect 5920 21916 7021 21944
rect 1578 21836 1584 21888
rect 1636 21876 1642 21888
rect 1765 21879 1823 21885
rect 1765 21876 1777 21879
rect 1636 21848 1777 21876
rect 1636 21836 1642 21848
rect 1765 21845 1777 21848
rect 1811 21845 1823 21879
rect 1765 21839 1823 21845
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 2409 21879 2467 21885
rect 2409 21876 2421 21879
rect 2280 21848 2421 21876
rect 2280 21836 2286 21848
rect 2409 21845 2421 21848
rect 2455 21845 2467 21879
rect 2409 21839 2467 21845
rect 2866 21836 2872 21888
rect 2924 21876 2930 21888
rect 3053 21879 3111 21885
rect 3053 21876 3065 21879
rect 2924 21848 3065 21876
rect 2924 21836 2930 21848
rect 3053 21845 3065 21848
rect 3099 21845 3111 21879
rect 3418 21876 3424 21888
rect 3379 21848 3424 21876
rect 3053 21839 3111 21845
rect 3418 21836 3424 21848
rect 3476 21836 3482 21888
rect 3602 21836 3608 21888
rect 3660 21876 3666 21888
rect 3881 21879 3939 21885
rect 3881 21876 3893 21879
rect 3660 21848 3893 21876
rect 3660 21836 3666 21848
rect 3881 21845 3893 21848
rect 3927 21845 3939 21879
rect 3881 21839 3939 21845
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4433 21879 4491 21885
rect 4433 21876 4445 21879
rect 4212 21848 4445 21876
rect 4212 21836 4218 21848
rect 4433 21845 4445 21848
rect 4479 21845 4491 21879
rect 4433 21839 4491 21845
rect 4706 21836 4712 21888
rect 4764 21876 4770 21888
rect 4801 21879 4859 21885
rect 4801 21876 4813 21879
rect 4764 21848 4813 21876
rect 4764 21836 4770 21848
rect 4801 21845 4813 21848
rect 4847 21845 4859 21879
rect 4801 21839 4859 21845
rect 4890 21836 4896 21888
rect 4948 21876 4954 21888
rect 5077 21879 5135 21885
rect 5077 21876 5089 21879
rect 4948 21848 5089 21876
rect 4948 21836 4954 21848
rect 5077 21845 5089 21848
rect 5123 21845 5135 21879
rect 5626 21876 5632 21888
rect 5587 21848 5632 21876
rect 5077 21839 5135 21845
rect 5626 21836 5632 21848
rect 5684 21836 5690 21888
rect 5920 21885 5948 21916
rect 7009 21913 7021 21916
rect 7055 21913 7067 21947
rect 7009 21907 7067 21913
rect 7374 21904 7380 21956
rect 7432 21904 7438 21956
rect 7469 21947 7527 21953
rect 7469 21913 7481 21947
rect 7515 21944 7527 21947
rect 8128 21944 8156 21984
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 9217 22015 9275 22021
rect 9217 22012 9229 22015
rect 9180 21984 9229 22012
rect 9180 21972 9186 21984
rect 9217 21981 9229 21984
rect 9263 21981 9275 22015
rect 9324 22012 9352 22052
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9646 22080 9674 22188
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 13357 22219 13415 22225
rect 13357 22185 13369 22219
rect 13403 22216 13415 22219
rect 13403 22188 13492 22216
rect 13403 22185 13415 22188
rect 13357 22179 13415 22185
rect 10781 22151 10839 22157
rect 10781 22117 10793 22151
rect 10827 22148 10839 22151
rect 13464 22148 13492 22188
rect 14366 22176 14372 22228
rect 14424 22216 14430 22228
rect 20901 22219 20959 22225
rect 20901 22216 20913 22219
rect 14424 22188 20913 22216
rect 14424 22176 14430 22188
rect 20901 22185 20913 22188
rect 20947 22216 20959 22219
rect 21634 22216 21640 22228
rect 20947 22188 21640 22216
rect 20947 22185 20959 22188
rect 20901 22179 20959 22185
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 22002 22216 22008 22228
rect 21963 22188 22008 22216
rect 22002 22176 22008 22188
rect 22060 22176 22066 22228
rect 14090 22148 14096 22160
rect 10827 22120 13216 22148
rect 13464 22120 14096 22148
rect 10827 22117 10839 22120
rect 10781 22111 10839 22117
rect 10226 22080 10232 22092
rect 9539 22052 9674 22080
rect 10187 22052 10232 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 10226 22040 10232 22052
rect 10284 22040 10290 22092
rect 12066 22080 12072 22092
rect 12027 22052 12072 22080
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 12158 22040 12164 22092
rect 12216 22080 12222 22092
rect 12216 22052 12261 22080
rect 12216 22040 12222 22052
rect 10870 22012 10876 22024
rect 9324 21984 10732 22012
rect 10831 21984 10876 22012
rect 9217 21975 9275 21981
rect 8481 21947 8539 21953
rect 8481 21944 8493 21947
rect 7515 21916 8064 21944
rect 8128 21916 8493 21944
rect 7515 21913 7527 21916
rect 7469 21907 7527 21913
rect 5905 21879 5963 21885
rect 5905 21845 5917 21879
rect 5951 21845 5963 21879
rect 5905 21839 5963 21845
rect 5994 21836 6000 21888
rect 6052 21876 6058 21888
rect 6052 21848 6097 21876
rect 6052 21836 6058 21848
rect 6178 21836 6184 21888
rect 6236 21876 6242 21888
rect 6365 21879 6423 21885
rect 6365 21876 6377 21879
rect 6236 21848 6377 21876
rect 6236 21836 6242 21848
rect 6365 21845 6377 21848
rect 6411 21845 6423 21879
rect 6365 21839 6423 21845
rect 6454 21836 6460 21888
rect 6512 21876 6518 21888
rect 6549 21879 6607 21885
rect 6549 21876 6561 21879
rect 6512 21848 6561 21876
rect 6512 21836 6518 21848
rect 6549 21845 6561 21848
rect 6595 21845 6607 21879
rect 6549 21839 6607 21845
rect 6638 21836 6644 21888
rect 6696 21876 6702 21888
rect 6917 21879 6975 21885
rect 6917 21876 6929 21879
rect 6696 21848 6929 21876
rect 6696 21836 6702 21848
rect 6917 21845 6929 21848
rect 6963 21845 6975 21879
rect 7558 21876 7564 21888
rect 7519 21848 7564 21876
rect 6917 21839 6975 21845
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 7926 21876 7932 21888
rect 7887 21848 7932 21876
rect 7926 21836 7932 21848
rect 7984 21836 7990 21888
rect 8036 21885 8064 21916
rect 8481 21913 8493 21916
rect 8527 21913 8539 21947
rect 8481 21907 8539 21913
rect 8662 21904 8668 21956
rect 8720 21944 8726 21956
rect 9677 21947 9735 21953
rect 9677 21944 9689 21947
rect 8720 21916 9689 21944
rect 8720 21904 8726 21916
rect 9677 21913 9689 21916
rect 9723 21913 9735 21947
rect 9677 21907 9735 21913
rect 10134 21904 10140 21956
rect 10192 21944 10198 21956
rect 10505 21947 10563 21953
rect 10505 21944 10517 21947
rect 10192 21916 10517 21944
rect 10192 21904 10198 21916
rect 10505 21913 10517 21916
rect 10551 21913 10563 21947
rect 10704 21944 10732 21984
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 11146 22012 11152 22024
rect 10980 21984 11152 22012
rect 10980 21944 11008 21984
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 22012 12955 22015
rect 13078 22012 13084 22024
rect 12943 21984 13084 22012
rect 12943 21981 12955 21984
rect 12897 21975 12955 21981
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 13188 22021 13216 22120
rect 14090 22108 14096 22120
rect 14148 22108 14154 22160
rect 14274 22108 14280 22160
rect 14332 22148 14338 22160
rect 14332 22120 16068 22148
rect 14332 22108 14338 22120
rect 13541 22083 13599 22089
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 14185 22083 14243 22089
rect 13587 22052 14136 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 22012 13231 22015
rect 13262 22012 13268 22024
rect 13219 21984 13268 22012
rect 13219 21981 13231 21984
rect 13173 21975 13231 21981
rect 13262 21972 13268 21984
rect 13320 21972 13326 22024
rect 13354 21972 13360 22024
rect 13412 22012 13418 22024
rect 13556 22012 13584 22043
rect 13412 21984 13584 22012
rect 13633 22015 13691 22021
rect 13412 21972 13418 21984
rect 13633 21981 13645 22015
rect 13679 21981 13691 22015
rect 14108 22012 14136 22052
rect 14185 22049 14197 22083
rect 14231 22080 14243 22083
rect 15562 22080 15568 22092
rect 14231 22052 15568 22080
rect 14231 22049 14243 22052
rect 14185 22043 14243 22049
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 16040 22080 16068 22120
rect 16114 22108 16120 22160
rect 16172 22148 16178 22160
rect 16172 22120 16804 22148
rect 16172 22108 16178 22120
rect 16776 22089 16804 22120
rect 18414 22108 18420 22160
rect 18472 22148 18478 22160
rect 19245 22151 19303 22157
rect 19245 22148 19257 22151
rect 18472 22120 19257 22148
rect 18472 22108 18478 22120
rect 19245 22117 19257 22120
rect 19291 22117 19303 22151
rect 20806 22148 20812 22160
rect 20767 22120 20812 22148
rect 19245 22111 19303 22117
rect 20806 22108 20812 22120
rect 20864 22108 20870 22160
rect 21726 22148 21732 22160
rect 21468 22120 21732 22148
rect 16301 22083 16359 22089
rect 16301 22080 16313 22083
rect 16040 22052 16313 22080
rect 16301 22049 16313 22052
rect 16347 22049 16359 22083
rect 16301 22043 16359 22049
rect 16761 22083 16819 22089
rect 16761 22049 16773 22083
rect 16807 22080 16819 22083
rect 17586 22080 17592 22092
rect 16807 22052 16841 22080
rect 17547 22052 17592 22080
rect 16807 22049 16819 22052
rect 16761 22043 16819 22049
rect 17586 22040 17592 22052
rect 17644 22040 17650 22092
rect 18509 22083 18567 22089
rect 18509 22049 18521 22083
rect 18555 22080 18567 22083
rect 18782 22080 18788 22092
rect 18555 22052 18788 22080
rect 18555 22049 18567 22052
rect 18509 22043 18567 22049
rect 18782 22040 18788 22052
rect 18840 22040 18846 22092
rect 19150 22040 19156 22092
rect 19208 22080 19214 22092
rect 19797 22083 19855 22089
rect 19797 22080 19809 22083
rect 19208 22052 19809 22080
rect 19208 22040 19214 22052
rect 19797 22049 19809 22052
rect 19843 22049 19855 22083
rect 20162 22080 20168 22092
rect 20123 22052 20168 22080
rect 19797 22043 19855 22049
rect 20162 22040 20168 22052
rect 20220 22040 20226 22092
rect 21468 22089 21496 22120
rect 21726 22108 21732 22120
rect 21784 22108 21790 22160
rect 21453 22083 21511 22089
rect 21453 22049 21465 22083
rect 21499 22080 21511 22083
rect 21499 22052 21533 22080
rect 21499 22049 21511 22052
rect 21453 22043 21511 22049
rect 22278 22040 22284 22092
rect 22336 22080 22342 22092
rect 22336 22052 22692 22080
rect 22336 22040 22342 22052
rect 14458 22012 14464 22024
rect 14108 21984 14464 22012
rect 13633 21975 13691 21981
rect 12437 21947 12495 21953
rect 12437 21944 12449 21947
rect 10704 21916 11008 21944
rect 11072 21916 12449 21944
rect 10505 21907 10563 21913
rect 8021 21879 8079 21885
rect 8021 21845 8033 21879
rect 8067 21845 8079 21879
rect 8021 21839 8079 21845
rect 8110 21836 8116 21888
rect 8168 21876 8174 21888
rect 8389 21879 8447 21885
rect 8389 21876 8401 21879
rect 8168 21848 8401 21876
rect 8168 21836 8174 21848
rect 8389 21845 8401 21848
rect 8435 21845 8447 21879
rect 8389 21839 8447 21845
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 9033 21879 9091 21885
rect 9033 21876 9045 21879
rect 8628 21848 9045 21876
rect 8628 21836 8634 21848
rect 9033 21845 9045 21848
rect 9079 21845 9091 21879
rect 9033 21839 9091 21845
rect 9306 21836 9312 21888
rect 9364 21876 9370 21888
rect 9585 21879 9643 21885
rect 9585 21876 9597 21879
rect 9364 21848 9597 21876
rect 9364 21836 9370 21848
rect 9585 21845 9597 21848
rect 9631 21845 9643 21879
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 9585 21839 9643 21845
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10410 21876 10416 21888
rect 10371 21848 10416 21876
rect 10410 21836 10416 21848
rect 10468 21836 10474 21888
rect 11072 21885 11100 21916
rect 12437 21913 12449 21916
rect 12483 21913 12495 21947
rect 12618 21944 12624 21956
rect 12579 21916 12624 21944
rect 12437 21907 12495 21913
rect 12618 21904 12624 21916
rect 12676 21904 12682 21956
rect 12805 21947 12863 21953
rect 12805 21913 12817 21947
rect 12851 21944 12863 21947
rect 13648 21944 13676 21975
rect 14458 21972 14464 21984
rect 14516 21972 14522 22024
rect 14642 21972 14648 22024
rect 14700 22012 14706 22024
rect 14921 22015 14979 22021
rect 14921 22012 14933 22015
rect 14700 21984 14933 22012
rect 14700 21972 14706 21984
rect 14921 21981 14933 21984
rect 14967 21981 14979 22015
rect 14921 21975 14979 21981
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 21981 15347 22015
rect 15289 21975 15347 21981
rect 12851 21916 13676 21944
rect 14553 21947 14611 21953
rect 12851 21913 12863 21916
rect 12805 21907 12863 21913
rect 14553 21913 14565 21947
rect 14599 21944 14611 21947
rect 15304 21944 15332 21975
rect 15470 21972 15476 22024
rect 15528 22012 15534 22024
rect 16666 22012 16672 22024
rect 15528 21984 15573 22012
rect 15856 21984 16672 22012
rect 15528 21972 15534 21984
rect 15856 21944 15884 21984
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 21818 22012 21824 22024
rect 18104 21984 19564 22012
rect 21779 21984 21824 22012
rect 18104 21972 18110 21984
rect 14599 21916 15884 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 15930 21904 15936 21956
rect 15988 21944 15994 21956
rect 16209 21947 16267 21953
rect 16209 21944 16221 21947
rect 15988 21916 16221 21944
rect 15988 21904 15994 21916
rect 16209 21913 16221 21916
rect 16255 21913 16267 21947
rect 16209 21907 16267 21913
rect 16945 21947 17003 21953
rect 16945 21913 16957 21947
rect 16991 21944 17003 21947
rect 17126 21944 17132 21956
rect 16991 21916 17132 21944
rect 16991 21913 17003 21916
rect 16945 21907 17003 21913
rect 17126 21904 17132 21916
rect 17184 21904 17190 21956
rect 17310 21904 17316 21956
rect 17368 21944 17374 21956
rect 17865 21947 17923 21953
rect 17865 21944 17877 21947
rect 17368 21916 17877 21944
rect 17368 21904 17374 21916
rect 17865 21913 17877 21916
rect 17911 21913 17923 21947
rect 17865 21907 17923 21913
rect 18138 21904 18144 21956
rect 18196 21944 18202 21956
rect 19334 21944 19340 21956
rect 18196 21916 19340 21944
rect 18196 21904 18202 21916
rect 19334 21904 19340 21916
rect 19392 21904 19398 21956
rect 19536 21944 19564 21984
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22189 22015 22247 22021
rect 22189 22012 22201 22015
rect 22152 21984 22201 22012
rect 22152 21972 22158 21984
rect 22189 21981 22201 21984
rect 22235 21981 22247 22015
rect 22554 22012 22560 22024
rect 22515 21984 22560 22012
rect 22189 21975 22247 21981
rect 22554 21972 22560 21984
rect 22612 21972 22618 22024
rect 20622 21944 20628 21956
rect 19536 21916 20628 21944
rect 20622 21904 20628 21916
rect 20680 21904 20686 21956
rect 20898 21904 20904 21956
rect 20956 21944 20962 21956
rect 20956 21916 22416 21944
rect 20956 21904 20962 21916
rect 11057 21879 11115 21885
rect 11057 21845 11069 21879
rect 11103 21845 11115 21879
rect 11330 21876 11336 21888
rect 11291 21848 11336 21876
rect 11057 21839 11115 21845
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 11609 21879 11667 21885
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11698 21876 11704 21888
rect 11655 21848 11704 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 11974 21876 11980 21888
rect 11935 21848 11980 21876
rect 11974 21836 11980 21848
rect 12032 21836 12038 21888
rect 13078 21876 13084 21888
rect 13039 21848 13084 21876
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 13817 21879 13875 21885
rect 13817 21845 13829 21879
rect 13863 21876 13875 21879
rect 14734 21876 14740 21888
rect 13863 21848 14740 21876
rect 13863 21845 13875 21848
rect 13817 21839 13875 21845
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 15102 21836 15108 21888
rect 15160 21876 15166 21888
rect 15197 21879 15255 21885
rect 15197 21876 15209 21879
rect 15160 21848 15209 21876
rect 15160 21836 15166 21848
rect 15197 21845 15209 21848
rect 15243 21845 15255 21879
rect 15654 21876 15660 21888
rect 15615 21848 15660 21876
rect 15197 21839 15255 21845
rect 15654 21836 15660 21848
rect 15712 21836 15718 21888
rect 15749 21879 15807 21885
rect 15749 21845 15761 21879
rect 15795 21876 15807 21879
rect 15838 21876 15844 21888
rect 15795 21848 15844 21876
rect 15795 21845 15807 21848
rect 15749 21839 15807 21845
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 16117 21879 16175 21885
rect 16117 21845 16129 21879
rect 16163 21876 16175 21879
rect 16298 21876 16304 21888
rect 16163 21848 16304 21876
rect 16163 21845 16175 21848
rect 16117 21839 16175 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 17037 21879 17095 21885
rect 17037 21845 17049 21879
rect 17083 21876 17095 21879
rect 17218 21876 17224 21888
rect 17083 21848 17224 21876
rect 17083 21845 17095 21848
rect 17037 21839 17095 21845
rect 17218 21836 17224 21848
rect 17276 21836 17282 21888
rect 17402 21876 17408 21888
rect 17363 21848 17408 21876
rect 17402 21836 17408 21848
rect 17460 21836 17466 21888
rect 17494 21836 17500 21888
rect 17552 21876 17558 21888
rect 17773 21879 17831 21885
rect 17773 21876 17785 21879
rect 17552 21848 17785 21876
rect 17552 21836 17558 21848
rect 17773 21845 17785 21848
rect 17819 21845 17831 21879
rect 18230 21876 18236 21888
rect 18191 21848 18236 21876
rect 17773 21839 17831 21845
rect 18230 21836 18236 21848
rect 18288 21836 18294 21888
rect 18598 21876 18604 21888
rect 18559 21848 18604 21876
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 18690 21836 18696 21888
rect 18748 21876 18754 21888
rect 19058 21876 19064 21888
rect 18748 21848 18793 21876
rect 19019 21848 19064 21876
rect 18748 21836 18754 21848
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19610 21876 19616 21888
rect 19571 21848 19616 21876
rect 19610 21836 19616 21848
rect 19668 21836 19674 21888
rect 19702 21836 19708 21888
rect 19760 21876 19766 21888
rect 20346 21876 20352 21888
rect 19760 21848 19805 21876
rect 20307 21848 20352 21876
rect 19760 21836 19766 21848
rect 20346 21836 20352 21848
rect 20404 21836 20410 21888
rect 20438 21836 20444 21888
rect 20496 21876 20502 21888
rect 21266 21876 21272 21888
rect 20496 21848 20541 21876
rect 21227 21848 21272 21876
rect 20496 21836 20502 21848
rect 21266 21836 21272 21848
rect 21324 21836 21330 21888
rect 21358 21836 21364 21888
rect 21416 21876 21422 21888
rect 22388 21885 22416 21916
rect 22373 21879 22431 21885
rect 21416 21848 21461 21876
rect 21416 21836 21422 21848
rect 22373 21845 22385 21879
rect 22419 21845 22431 21879
rect 22664 21876 22692 22052
rect 23109 22015 23167 22021
rect 23109 21981 23121 22015
rect 23155 22012 23167 22015
rect 23198 22012 23204 22024
rect 23155 21984 23204 22012
rect 23155 21981 23167 21984
rect 23109 21975 23167 21981
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 22741 21879 22799 21885
rect 22741 21876 22753 21879
rect 22664 21848 22753 21876
rect 22373 21839 22431 21845
rect 22741 21845 22753 21848
rect 22787 21845 22799 21879
rect 22741 21839 22799 21845
rect 22925 21879 22983 21885
rect 22925 21845 22937 21879
rect 22971 21876 22983 21879
rect 23382 21876 23388 21888
rect 22971 21848 23388 21876
rect 22971 21845 22983 21848
rect 22925 21839 22983 21845
rect 23382 21836 23388 21848
rect 23440 21836 23446 21888
rect 1104 21786 23460 21808
rect 1104 21734 6548 21786
rect 6600 21734 6612 21786
rect 6664 21734 6676 21786
rect 6728 21734 6740 21786
rect 6792 21734 6804 21786
rect 6856 21734 12146 21786
rect 12198 21734 12210 21786
rect 12262 21734 12274 21786
rect 12326 21734 12338 21786
rect 12390 21734 12402 21786
rect 12454 21734 17744 21786
rect 17796 21734 17808 21786
rect 17860 21734 17872 21786
rect 17924 21734 17936 21786
rect 17988 21734 18000 21786
rect 18052 21734 23460 21786
rect 1104 21712 23460 21734
rect 290 21632 296 21684
rect 348 21672 354 21684
rect 1489 21675 1547 21681
rect 1489 21672 1501 21675
rect 348 21644 1501 21672
rect 348 21632 354 21644
rect 1489 21641 1501 21644
rect 1535 21641 1547 21675
rect 2133 21675 2191 21681
rect 2133 21672 2145 21675
rect 1489 21635 1547 21641
rect 1688 21644 2145 21672
rect 1688 21545 1716 21644
rect 2133 21641 2145 21644
rect 2179 21641 2191 21675
rect 2133 21635 2191 21641
rect 2409 21675 2467 21681
rect 2409 21641 2421 21675
rect 2455 21641 2467 21675
rect 2409 21635 2467 21641
rect 2424 21604 2452 21635
rect 2682 21632 2688 21684
rect 2740 21672 2746 21684
rect 2869 21675 2927 21681
rect 2869 21672 2881 21675
rect 2740 21644 2881 21672
rect 2740 21632 2746 21644
rect 2869 21641 2881 21644
rect 2915 21641 2927 21675
rect 2869 21635 2927 21641
rect 3234 21632 3240 21684
rect 3292 21672 3298 21684
rect 3513 21675 3571 21681
rect 3513 21672 3525 21675
rect 3292 21644 3525 21672
rect 3292 21632 3298 21644
rect 3513 21641 3525 21644
rect 3559 21641 3571 21675
rect 3513 21635 3571 21641
rect 4062 21632 4068 21684
rect 4120 21672 4126 21684
rect 4341 21675 4399 21681
rect 4341 21672 4353 21675
rect 4120 21644 4353 21672
rect 4120 21632 4126 21644
rect 4341 21641 4353 21644
rect 4387 21641 4399 21675
rect 5442 21672 5448 21684
rect 4341 21635 4399 21641
rect 4448 21644 5448 21672
rect 2056 21576 2452 21604
rect 2777 21607 2835 21613
rect 2056 21545 2084 21576
rect 2777 21573 2789 21607
rect 2823 21604 2835 21607
rect 3142 21604 3148 21616
rect 2823 21576 3148 21604
rect 2823 21573 2835 21576
rect 2777 21567 2835 21573
rect 3142 21564 3148 21576
rect 3200 21564 3206 21616
rect 4448 21604 4476 21644
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 5905 21675 5963 21681
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 7558 21672 7564 21684
rect 5951 21644 7564 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 7558 21632 7564 21644
rect 7616 21632 7622 21684
rect 8573 21675 8631 21681
rect 8573 21641 8585 21675
rect 8619 21672 8631 21675
rect 9306 21672 9312 21684
rect 8619 21644 9312 21672
rect 8619 21641 8631 21644
rect 8573 21635 8631 21641
rect 9306 21632 9312 21644
rect 9364 21632 9370 21684
rect 9398 21632 9404 21684
rect 9456 21672 9462 21684
rect 10226 21672 10232 21684
rect 9456 21644 9501 21672
rect 9600 21644 10232 21672
rect 9456 21632 9462 21644
rect 3252 21576 4476 21604
rect 3252 21548 3280 21576
rect 4706 21564 4712 21616
rect 4764 21604 4770 21616
rect 6549 21607 6607 21613
rect 4764 21576 5764 21604
rect 4764 21564 4770 21576
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21505 2099 21539
rect 2314 21536 2320 21548
rect 2275 21508 2320 21536
rect 2041 21499 2099 21505
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21536 2651 21539
rect 2682 21536 2688 21548
rect 2639 21508 2688 21536
rect 2639 21505 2651 21508
rect 2593 21499 2651 21505
rect 2682 21496 2688 21508
rect 2740 21496 2746 21548
rect 3050 21536 3056 21548
rect 3011 21508 3056 21536
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 3234 21496 3240 21548
rect 3292 21496 3298 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 3344 21508 3433 21536
rect 2866 21428 2872 21480
rect 2924 21468 2930 21480
rect 3344 21468 3372 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 3510 21496 3516 21548
rect 3568 21536 3574 21548
rect 3697 21539 3755 21545
rect 3697 21536 3709 21539
rect 3568 21508 3709 21536
rect 3568 21496 3574 21508
rect 3697 21505 3709 21508
rect 3743 21505 3755 21539
rect 3697 21499 3755 21505
rect 3786 21496 3792 21548
rect 3844 21536 3850 21548
rect 3844 21508 3889 21536
rect 3844 21496 3850 21508
rect 3970 21496 3976 21548
rect 4028 21536 4034 21548
rect 4065 21539 4123 21545
rect 4065 21536 4077 21539
rect 4028 21508 4077 21536
rect 4028 21496 4034 21508
rect 4065 21505 4077 21508
rect 4111 21505 4123 21539
rect 4522 21536 4528 21548
rect 4483 21508 4528 21536
rect 4065 21499 4123 21505
rect 4522 21496 4528 21508
rect 4580 21496 4586 21548
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21536 4675 21539
rect 4982 21536 4988 21548
rect 4663 21508 4988 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 2924 21440 3372 21468
rect 2924 21428 2930 21440
rect 934 21360 940 21412
rect 992 21400 998 21412
rect 1857 21403 1915 21409
rect 1857 21400 1869 21403
rect 992 21372 1869 21400
rect 992 21360 998 21372
rect 1857 21369 1869 21372
rect 1903 21369 1915 21403
rect 1857 21363 1915 21369
rect 2590 21360 2596 21412
rect 2648 21400 2654 21412
rect 3237 21403 3295 21409
rect 3237 21400 3249 21403
rect 2648 21372 3249 21400
rect 2648 21360 2654 21372
rect 3237 21369 3249 21372
rect 3283 21369 3295 21403
rect 3344 21400 3372 21440
rect 4154 21428 4160 21480
rect 4212 21468 4218 21480
rect 4632 21468 4660 21499
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 5077 21539 5135 21545
rect 5077 21505 5089 21539
rect 5123 21505 5135 21539
rect 5077 21499 5135 21505
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21536 5411 21539
rect 5442 21536 5448 21548
rect 5399 21508 5448 21536
rect 5399 21505 5411 21508
rect 5353 21499 5411 21505
rect 4212 21440 4660 21468
rect 4212 21428 4218 21440
rect 4890 21428 4896 21480
rect 4948 21468 4954 21480
rect 5092 21468 5120 21499
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 5626 21536 5632 21548
rect 5587 21508 5632 21536
rect 5626 21496 5632 21508
rect 5684 21496 5690 21548
rect 5736 21536 5764 21576
rect 6549 21573 6561 21607
rect 6595 21604 6607 21607
rect 9033 21607 9091 21613
rect 9033 21604 9045 21607
rect 6595 21576 9045 21604
rect 6595 21573 6607 21576
rect 6549 21567 6607 21573
rect 9033 21573 9045 21576
rect 9079 21573 9091 21607
rect 9600 21604 9628 21644
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 10502 21632 10508 21684
rect 10560 21672 10566 21684
rect 11793 21675 11851 21681
rect 11793 21672 11805 21675
rect 10560 21644 11805 21672
rect 10560 21632 10566 21644
rect 11793 21641 11805 21644
rect 11839 21641 11851 21675
rect 11793 21635 11851 21641
rect 12066 21632 12072 21684
rect 12124 21672 12130 21684
rect 12253 21675 12311 21681
rect 12253 21672 12265 21675
rect 12124 21644 12265 21672
rect 12124 21632 12130 21644
rect 12253 21641 12265 21644
rect 12299 21641 12311 21675
rect 13906 21672 13912 21684
rect 12253 21635 12311 21641
rect 12406 21644 13912 21672
rect 9033 21567 9091 21573
rect 9324 21576 9628 21604
rect 6825 21539 6883 21545
rect 6825 21536 6837 21539
rect 5736 21508 6837 21536
rect 6825 21505 6837 21508
rect 6871 21505 6883 21539
rect 7374 21536 7380 21548
rect 7335 21508 7380 21536
rect 6825 21499 6883 21505
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 8018 21536 8024 21548
rect 7944 21508 8024 21536
rect 6086 21468 6092 21480
rect 4948 21440 6092 21468
rect 4948 21428 4954 21440
rect 6086 21428 6092 21440
rect 6144 21428 6150 21480
rect 6181 21471 6239 21477
rect 6181 21437 6193 21471
rect 6227 21468 6239 21471
rect 7282 21468 7288 21480
rect 6227 21440 6500 21468
rect 6227 21437 6239 21440
rect 6181 21431 6239 21437
rect 6472 21412 6500 21440
rect 6748 21440 7288 21468
rect 4430 21400 4436 21412
rect 3344 21372 4436 21400
rect 3237 21363 3295 21369
rect 4430 21360 4436 21372
rect 4488 21360 4494 21412
rect 4798 21400 4804 21412
rect 4759 21372 4804 21400
rect 4798 21360 4804 21372
rect 4856 21360 4862 21412
rect 5166 21400 5172 21412
rect 5127 21372 5172 21400
rect 5166 21360 5172 21372
rect 5224 21360 5230 21412
rect 5350 21360 5356 21412
rect 5408 21400 5414 21412
rect 5994 21400 6000 21412
rect 5408 21372 6000 21400
rect 5408 21360 5414 21372
rect 5994 21360 6000 21372
rect 6052 21360 6058 21412
rect 6454 21360 6460 21412
rect 6512 21360 6518 21412
rect 6638 21400 6644 21412
rect 6599 21372 6644 21400
rect 6638 21360 6644 21372
rect 6696 21360 6702 21412
rect 2498 21292 2504 21344
rect 2556 21332 2562 21344
rect 3878 21332 3884 21344
rect 2556 21304 3884 21332
rect 2556 21292 2562 21304
rect 3878 21292 3884 21304
rect 3936 21292 3942 21344
rect 3973 21335 4031 21341
rect 3973 21301 3985 21335
rect 4019 21332 4031 21335
rect 4062 21332 4068 21344
rect 4019 21304 4068 21332
rect 4019 21301 4031 21304
rect 3973 21295 4031 21301
rect 4062 21292 4068 21304
rect 4120 21292 4126 21344
rect 4246 21332 4252 21344
rect 4207 21304 4252 21332
rect 4246 21292 4252 21304
rect 4304 21292 4310 21344
rect 4338 21292 4344 21344
rect 4396 21332 4402 21344
rect 4893 21335 4951 21341
rect 4893 21332 4905 21335
rect 4396 21304 4905 21332
rect 4396 21292 4402 21304
rect 4893 21301 4905 21304
rect 4939 21301 4951 21335
rect 4893 21295 4951 21301
rect 4982 21292 4988 21344
rect 5040 21332 5046 21344
rect 5258 21332 5264 21344
rect 5040 21304 5264 21332
rect 5040 21292 5046 21304
rect 5258 21292 5264 21304
rect 5316 21292 5322 21344
rect 5442 21332 5448 21344
rect 5403 21304 5448 21332
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 5534 21292 5540 21344
rect 5592 21332 5598 21344
rect 6748 21332 6776 21440
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 7469 21471 7527 21477
rect 7469 21437 7481 21471
rect 7515 21437 7527 21471
rect 7469 21431 7527 21437
rect 7484 21400 7512 21431
rect 7558 21428 7564 21480
rect 7616 21468 7622 21480
rect 7944 21477 7972 21508
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 8202 21536 8208 21548
rect 8163 21508 8208 21536
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 9324 21536 9352 21576
rect 11146 21564 11152 21616
rect 11204 21604 11210 21616
rect 12406 21604 12434 21644
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 14553 21675 14611 21681
rect 14553 21641 14565 21675
rect 14599 21641 14611 21675
rect 14553 21635 14611 21641
rect 11204 21576 12434 21604
rect 11204 21564 11210 21576
rect 12526 21564 12532 21616
rect 12584 21604 12590 21616
rect 12621 21607 12679 21613
rect 12621 21604 12633 21607
rect 12584 21576 12633 21604
rect 12584 21564 12590 21576
rect 12621 21573 12633 21576
rect 12667 21604 12679 21607
rect 12710 21604 12716 21616
rect 12667 21576 12716 21604
rect 12667 21573 12679 21576
rect 12621 21567 12679 21573
rect 12710 21564 12716 21576
rect 12768 21564 12774 21616
rect 14568 21604 14596 21635
rect 15654 21632 15660 21684
rect 15712 21672 15718 21684
rect 16025 21675 16083 21681
rect 16025 21672 16037 21675
rect 15712 21644 16037 21672
rect 15712 21632 15718 21644
rect 16025 21641 16037 21644
rect 16071 21641 16083 21675
rect 16025 21635 16083 21641
rect 16298 21632 16304 21684
rect 16356 21672 16362 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16356 21644 17049 21672
rect 16356 21632 16362 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 17037 21635 17095 21641
rect 17405 21675 17463 21681
rect 17405 21641 17417 21675
rect 17451 21672 17463 21675
rect 17494 21672 17500 21684
rect 17451 21644 17500 21672
rect 17451 21641 17463 21644
rect 17405 21635 17463 21641
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 18322 21632 18328 21684
rect 18380 21672 18386 21684
rect 18699 21675 18757 21681
rect 18699 21672 18711 21675
rect 18380 21644 18711 21672
rect 18380 21632 18386 21644
rect 18699 21641 18711 21644
rect 18745 21641 18757 21675
rect 18699 21635 18757 21641
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 19116 21644 19748 21672
rect 19116 21632 19122 21644
rect 14568 21576 16804 21604
rect 10229 21539 10287 21545
rect 10229 21536 10241 21539
rect 8772 21508 9352 21536
rect 9416 21508 10241 21536
rect 7929 21471 7987 21477
rect 7616 21440 7661 21468
rect 7616 21428 7622 21440
rect 7929 21437 7941 21471
rect 7975 21437 7987 21471
rect 8110 21468 8116 21480
rect 8071 21440 8116 21468
rect 7929 21431 7987 21437
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 8772 21477 8800 21508
rect 8757 21471 8815 21477
rect 8757 21437 8769 21471
rect 8803 21437 8815 21471
rect 8938 21468 8944 21480
rect 8899 21440 8944 21468
rect 8757 21431 8815 21437
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9416 21400 9444 21508
rect 10229 21505 10241 21508
rect 10275 21536 10287 21539
rect 10686 21536 10692 21548
rect 10275 21508 10692 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 11606 21496 11612 21548
rect 11664 21536 11670 21548
rect 11885 21539 11943 21545
rect 11885 21536 11897 21539
rect 11664 21508 11897 21536
rect 11664 21496 11670 21508
rect 11885 21505 11897 21508
rect 11931 21505 11943 21539
rect 12437 21539 12495 21545
rect 12437 21536 12449 21539
rect 11885 21499 11943 21505
rect 11992 21508 12449 21536
rect 9490 21428 9496 21480
rect 9548 21468 9554 21480
rect 9858 21477 9864 21480
rect 9816 21471 9864 21477
rect 9548 21440 9593 21468
rect 9548 21428 9554 21440
rect 9816 21437 9828 21471
rect 9862 21437 9864 21471
rect 9816 21431 9864 21437
rect 9858 21428 9864 21431
rect 9916 21428 9922 21480
rect 9999 21471 10057 21477
rect 9999 21437 10011 21471
rect 10045 21468 10057 21471
rect 10318 21468 10324 21480
rect 10045 21440 10324 21468
rect 10045 21437 10057 21440
rect 9999 21431 10057 21437
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 10410 21428 10416 21480
rect 10468 21468 10474 21480
rect 11701 21471 11759 21477
rect 10468 21440 11652 21468
rect 10468 21428 10474 21440
rect 7484 21372 9444 21400
rect 11624 21400 11652 21440
rect 11701 21437 11713 21471
rect 11747 21468 11759 21471
rect 11790 21468 11796 21480
rect 11747 21440 11796 21468
rect 11747 21437 11759 21440
rect 11701 21431 11759 21437
rect 11790 21428 11796 21440
rect 11848 21428 11854 21480
rect 11992 21400 12020 21508
rect 12437 21505 12449 21508
rect 12483 21505 12495 21539
rect 12728 21536 12756 21564
rect 12728 21508 13079 21536
rect 12437 21499 12495 21505
rect 12713 21471 12771 21477
rect 12713 21437 12725 21471
rect 12759 21468 12771 21471
rect 12894 21468 12900 21480
rect 12759 21440 12900 21468
rect 12759 21437 12771 21440
rect 12713 21431 12771 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 13051 21477 13079 21508
rect 14458 21496 14464 21548
rect 14516 21536 14522 21548
rect 14921 21539 14979 21545
rect 14921 21536 14933 21539
rect 14516 21508 14933 21536
rect 14516 21496 14522 21508
rect 14921 21505 14933 21508
rect 14967 21505 14979 21539
rect 14921 21499 14979 21505
rect 15013 21539 15071 21545
rect 15013 21505 15025 21539
rect 15059 21505 15071 21539
rect 16114 21536 16120 21548
rect 15013 21499 15071 21505
rect 15856 21508 16120 21536
rect 13036 21471 13094 21477
rect 13036 21437 13048 21471
rect 13082 21437 13094 21471
rect 13036 21431 13094 21437
rect 13176 21471 13234 21477
rect 13176 21437 13188 21471
rect 13222 21468 13234 21471
rect 13262 21468 13268 21480
rect 13222 21440 13268 21468
rect 13222 21437 13234 21440
rect 13176 21431 13234 21437
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 13446 21468 13452 21480
rect 13407 21440 13452 21468
rect 13446 21428 13452 21440
rect 13504 21468 13510 21480
rect 14366 21468 14372 21480
rect 13504 21440 14372 21468
rect 13504 21428 13510 21440
rect 14366 21428 14372 21440
rect 14424 21428 14430 21480
rect 14734 21468 14740 21480
rect 14695 21440 14740 21468
rect 14734 21428 14740 21440
rect 14792 21428 14798 21480
rect 11624 21372 12020 21400
rect 7006 21332 7012 21344
rect 5592 21304 6776 21332
rect 6967 21304 7012 21332
rect 5592 21292 5598 21304
rect 7006 21292 7012 21304
rect 7064 21292 7070 21344
rect 8110 21292 8116 21344
rect 8168 21332 8174 21344
rect 9674 21332 9680 21344
rect 8168 21304 9680 21332
rect 8168 21292 8174 21304
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11333 21335 11391 21341
rect 11333 21332 11345 21335
rect 11112 21304 11345 21332
rect 11112 21292 11118 21304
rect 11333 21301 11345 21304
rect 11379 21332 11391 21335
rect 12066 21332 12072 21344
rect 11379 21304 12072 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 15028 21332 15056 21499
rect 15856 21480 15884 21508
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 16776 21536 16804 21576
rect 16850 21564 16856 21616
rect 16908 21604 16914 21616
rect 17681 21607 17739 21613
rect 17681 21604 17693 21607
rect 16908 21576 17693 21604
rect 16908 21564 16914 21576
rect 17681 21573 17693 21576
rect 17727 21573 17739 21607
rect 19720 21604 19748 21644
rect 19794 21632 19800 21684
rect 19852 21672 19858 21684
rect 20438 21672 20444 21684
rect 19852 21644 20444 21672
rect 19852 21632 19858 21644
rect 20438 21632 20444 21644
rect 20496 21632 20502 21684
rect 20533 21675 20591 21681
rect 20533 21641 20545 21675
rect 20579 21672 20591 21675
rect 20806 21672 20812 21684
rect 20579 21644 20812 21672
rect 20579 21641 20591 21644
rect 20533 21635 20591 21641
rect 20806 21632 20812 21644
rect 20864 21632 20870 21684
rect 20901 21675 20959 21681
rect 20901 21641 20913 21675
rect 20947 21672 20959 21675
rect 21358 21672 21364 21684
rect 20947 21644 21364 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 21542 21632 21548 21684
rect 21600 21672 21606 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 21600 21644 22017 21672
rect 21600 21632 21606 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22005 21635 22063 21641
rect 22189 21675 22247 21681
rect 22189 21641 22201 21675
rect 22235 21641 22247 21675
rect 22189 21635 22247 21641
rect 22649 21675 22707 21681
rect 22649 21641 22661 21675
rect 22695 21672 22707 21675
rect 22830 21672 22836 21684
rect 22695 21644 22836 21672
rect 22695 21641 22707 21644
rect 22649 21635 22707 21641
rect 21910 21604 21916 21616
rect 19720 21576 21916 21604
rect 17681 21567 17739 21573
rect 21910 21564 21916 21576
rect 21968 21564 21974 21616
rect 22204 21604 22232 21635
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 22020 21576 22232 21604
rect 16945 21539 17003 21545
rect 16945 21536 16957 21539
rect 16776 21508 16957 21536
rect 16945 21505 16957 21508
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 15838 21468 15844 21480
rect 15799 21440 15844 21468
rect 15838 21428 15844 21440
rect 15896 21428 15902 21480
rect 15933 21471 15991 21477
rect 15933 21437 15945 21471
rect 15979 21437 15991 21471
rect 15933 21431 15991 21437
rect 15381 21403 15439 21409
rect 15381 21369 15393 21403
rect 15427 21400 15439 21403
rect 15948 21400 15976 21431
rect 16574 21428 16580 21480
rect 16632 21468 16638 21480
rect 16761 21471 16819 21477
rect 16761 21468 16773 21471
rect 16632 21440 16773 21468
rect 16632 21428 16638 21440
rect 16761 21437 16773 21440
rect 16807 21437 16819 21471
rect 16960 21468 16988 21499
rect 17034 21496 17040 21548
rect 17092 21536 17098 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17092 21508 17509 21536
rect 17092 21496 17098 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 18138 21536 18144 21548
rect 18099 21508 18144 21536
rect 17497 21499 17555 21505
rect 18138 21496 18144 21508
rect 18196 21496 18202 21548
rect 18506 21536 18512 21548
rect 18248 21508 18512 21536
rect 18046 21468 18052 21480
rect 16960 21440 18052 21468
rect 16761 21431 16819 21437
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 18248 21477 18276 21508
rect 18506 21496 18512 21508
rect 18564 21496 18570 21548
rect 19242 21496 19248 21548
rect 19300 21496 19306 21548
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 19392 21508 21005 21536
rect 19392 21496 19398 21508
rect 20993 21505 21005 21508
rect 21039 21505 21051 21539
rect 21358 21536 21364 21548
rect 21319 21508 21364 21536
rect 20993 21499 21051 21505
rect 21358 21496 21364 21508
rect 21416 21496 21422 21548
rect 21450 21496 21456 21548
rect 21508 21536 21514 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21508 21508 21833 21536
rect 21508 21496 21514 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 18233 21471 18291 21477
rect 18233 21437 18245 21471
rect 18279 21437 18291 21471
rect 18233 21431 18291 21437
rect 18414 21428 18420 21480
rect 18472 21468 18478 21480
rect 18739 21473 18797 21479
rect 18739 21468 18751 21473
rect 18472 21440 18751 21468
rect 18472 21428 18478 21440
rect 18739 21439 18751 21440
rect 18785 21439 18797 21473
rect 18739 21433 18797 21439
rect 18969 21471 19027 21477
rect 18969 21437 18981 21471
rect 19015 21470 19027 21471
rect 19015 21468 19104 21470
rect 19260 21468 19288 21496
rect 19886 21468 19892 21480
rect 19015 21442 19892 21468
rect 19015 21437 19027 21442
rect 19076 21440 19892 21442
rect 18969 21431 19027 21437
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 19978 21428 19984 21480
rect 20036 21468 20042 21480
rect 20257 21471 20315 21477
rect 20257 21468 20269 21471
rect 20036 21440 20269 21468
rect 20036 21428 20042 21440
rect 20257 21437 20269 21440
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 20441 21471 20499 21477
rect 20441 21437 20453 21471
rect 20487 21437 20499 21471
rect 20441 21431 20499 21437
rect 17957 21403 18015 21409
rect 17957 21400 17969 21403
rect 15427 21372 15884 21400
rect 15948 21372 17969 21400
rect 15427 21369 15439 21372
rect 15381 21363 15439 21369
rect 15562 21332 15568 21344
rect 12768 21304 15056 21332
rect 15523 21304 15568 21332
rect 12768 21292 12774 21304
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 15856 21332 15884 21372
rect 17957 21369 17969 21372
rect 18003 21369 18015 21403
rect 17957 21363 18015 21369
rect 16298 21332 16304 21344
rect 15856 21304 16304 21332
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 16393 21335 16451 21341
rect 16393 21301 16405 21335
rect 16439 21332 16451 21335
rect 16482 21332 16488 21344
rect 16439 21304 16488 21332
rect 16439 21301 16451 21304
rect 16393 21295 16451 21301
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 17865 21335 17923 21341
rect 17865 21301 17877 21335
rect 17911 21332 17923 21335
rect 18230 21332 18236 21344
rect 17911 21304 18236 21332
rect 17911 21301 17923 21304
rect 17865 21295 17923 21301
rect 18230 21292 18236 21304
rect 18288 21292 18294 21344
rect 18414 21292 18420 21344
rect 18472 21332 18478 21344
rect 20073 21335 20131 21341
rect 20073 21332 20085 21335
rect 18472 21304 20085 21332
rect 18472 21292 18478 21304
rect 20073 21301 20085 21304
rect 20119 21332 20131 21335
rect 20456 21332 20484 21431
rect 21082 21428 21088 21480
rect 21140 21468 21146 21480
rect 22020 21468 22048 21576
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22244 21508 22385 21536
rect 22244 21496 22250 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22462 21496 22468 21548
rect 22520 21536 22526 21548
rect 22520 21508 22565 21536
rect 22520 21496 22526 21508
rect 22738 21496 22744 21548
rect 22796 21536 22802 21548
rect 22833 21539 22891 21545
rect 22833 21536 22845 21539
rect 22796 21508 22845 21536
rect 22796 21496 22802 21508
rect 22833 21505 22845 21508
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 21140 21440 22048 21468
rect 21140 21428 21146 21440
rect 20714 21360 20720 21412
rect 20772 21400 20778 21412
rect 21545 21403 21603 21409
rect 21545 21400 21557 21403
rect 20772 21372 21557 21400
rect 20772 21360 20778 21372
rect 21545 21369 21557 21372
rect 21591 21369 21603 21403
rect 21545 21363 21603 21369
rect 20119 21304 20484 21332
rect 20119 21301 20131 21304
rect 20073 21295 20131 21301
rect 20806 21292 20812 21344
rect 20864 21332 20870 21344
rect 21177 21335 21235 21341
rect 21177 21332 21189 21335
rect 20864 21304 21189 21332
rect 20864 21292 20870 21304
rect 21177 21301 21189 21304
rect 21223 21301 21235 21335
rect 23014 21332 23020 21344
rect 22975 21304 23020 21332
rect 21177 21295 21235 21301
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 1104 21242 23460 21264
rect 1104 21190 3749 21242
rect 3801 21190 3813 21242
rect 3865 21190 3877 21242
rect 3929 21190 3941 21242
rect 3993 21190 4005 21242
rect 4057 21190 9347 21242
rect 9399 21190 9411 21242
rect 9463 21190 9475 21242
rect 9527 21190 9539 21242
rect 9591 21190 9603 21242
rect 9655 21190 14945 21242
rect 14997 21190 15009 21242
rect 15061 21190 15073 21242
rect 15125 21190 15137 21242
rect 15189 21190 15201 21242
rect 15253 21190 20543 21242
rect 20595 21190 20607 21242
rect 20659 21190 20671 21242
rect 20723 21190 20735 21242
rect 20787 21190 20799 21242
rect 20851 21190 23460 21242
rect 1104 21168 23460 21190
rect 2498 21128 2504 21140
rect 2459 21100 2504 21128
rect 2498 21088 2504 21100
rect 2556 21088 2562 21140
rect 2774 21088 2780 21140
rect 2832 21128 2838 21140
rect 3053 21131 3111 21137
rect 2832 21100 2877 21128
rect 2832 21088 2838 21100
rect 3053 21097 3065 21131
rect 3099 21128 3111 21131
rect 3234 21128 3240 21140
rect 3099 21100 3240 21128
rect 3099 21097 3111 21100
rect 3053 21091 3111 21097
rect 3234 21088 3240 21100
rect 3292 21088 3298 21140
rect 3329 21131 3387 21137
rect 3329 21097 3341 21131
rect 3375 21128 3387 21131
rect 5718 21128 5724 21140
rect 3375 21100 5724 21128
rect 3375 21097 3387 21100
rect 3329 21091 3387 21097
rect 5718 21088 5724 21100
rect 5776 21088 5782 21140
rect 5997 21131 6055 21137
rect 5997 21097 6009 21131
rect 6043 21128 6055 21131
rect 7374 21128 7380 21140
rect 6043 21100 7380 21128
rect 6043 21097 6055 21100
rect 5997 21091 6055 21097
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 7926 21088 7932 21140
rect 7984 21128 7990 21140
rect 7984 21100 8800 21128
rect 7984 21088 7990 21100
rect 3786 21020 3792 21072
rect 3844 21060 3850 21072
rect 6822 21060 6828 21072
rect 3844 21032 6828 21060
rect 3844 21020 3850 21032
rect 6822 21020 6828 21032
rect 6880 21020 6886 21072
rect 6917 21063 6975 21069
rect 6917 21029 6929 21063
rect 6963 21060 6975 21063
rect 6963 21032 7420 21060
rect 6963 21029 6975 21032
rect 6917 21023 6975 21029
rect 2961 20995 3019 21001
rect 2961 20961 2973 20995
rect 3007 20992 3019 20995
rect 3142 20992 3148 21004
rect 3007 20964 3148 20992
rect 3007 20961 3019 20964
rect 2961 20955 3019 20961
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 5445 20995 5503 21001
rect 5445 20961 5457 20995
rect 5491 20992 5503 20995
rect 5534 20992 5540 21004
rect 5491 20964 5540 20992
rect 5491 20961 5503 20964
rect 5445 20955 5503 20961
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 5718 20992 5724 21004
rect 5644 20964 5724 20992
rect 2038 20924 2044 20936
rect 1999 20896 2044 20924
rect 2038 20884 2044 20896
rect 2096 20884 2102 20936
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20924 2283 20927
rect 3050 20924 3056 20936
rect 2271 20896 3056 20924
rect 2271 20893 2283 20896
rect 2225 20887 2283 20893
rect 3050 20884 3056 20896
rect 3108 20924 3114 20936
rect 3418 20924 3424 20936
rect 3108 20896 3424 20924
rect 3108 20884 3114 20896
rect 3418 20884 3424 20896
rect 3476 20884 3482 20936
rect 3602 20924 3608 20936
rect 3563 20896 3608 20924
rect 3602 20884 3608 20896
rect 3660 20884 3666 20936
rect 3694 20884 3700 20936
rect 3752 20924 3758 20936
rect 3881 20927 3939 20933
rect 3881 20924 3893 20927
rect 3752 20896 3893 20924
rect 3752 20884 3758 20896
rect 3881 20893 3893 20896
rect 3927 20893 3939 20927
rect 4338 20924 4344 20936
rect 4299 20896 4344 20924
rect 3881 20887 3939 20893
rect 4338 20884 4344 20896
rect 4396 20884 4402 20936
rect 4893 20927 4951 20933
rect 4893 20893 4905 20927
rect 4939 20924 4951 20927
rect 4982 20924 4988 20936
rect 4939 20896 4988 20924
rect 4939 20893 4951 20896
rect 4893 20887 4951 20893
rect 4982 20884 4988 20896
rect 5040 20884 5046 20936
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20924 5227 20927
rect 5350 20924 5356 20936
rect 5215 20896 5356 20924
rect 5215 20893 5227 20896
rect 5169 20887 5227 20893
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 5644 20933 5672 20964
rect 5718 20952 5724 20964
rect 5776 20952 5782 21004
rect 6178 20992 6184 21004
rect 6139 20964 6184 20992
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6365 20995 6423 21001
rect 6365 20961 6377 20995
rect 6411 20992 6423 20995
rect 7006 20992 7012 21004
rect 6411 20964 7012 20992
rect 6411 20961 6423 20964
rect 6365 20955 6423 20961
rect 7006 20952 7012 20964
rect 7064 20952 7070 21004
rect 7392 20992 7420 21032
rect 8110 20992 8116 21004
rect 7392 20964 8116 20992
rect 8110 20952 8116 20964
rect 8168 20952 8174 21004
rect 8202 20952 8208 21004
rect 8260 20992 8266 21004
rect 8294 20995 8352 21001
rect 8294 20992 8306 20995
rect 8260 20964 8306 20992
rect 8260 20952 8266 20964
rect 8294 20961 8306 20964
rect 8340 20961 8352 20995
rect 8772 20992 8800 21100
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 9214 21128 9220 21140
rect 8904 21100 9220 21128
rect 8904 21088 8910 21100
rect 9214 21088 9220 21100
rect 9272 21088 9278 21140
rect 9490 21088 9496 21140
rect 9548 21128 9554 21140
rect 11057 21131 11115 21137
rect 11057 21128 11069 21131
rect 9548 21100 11069 21128
rect 9548 21088 9554 21100
rect 11057 21097 11069 21100
rect 11103 21097 11115 21131
rect 11057 21091 11115 21097
rect 11330 21088 11336 21140
rect 11388 21128 11394 21140
rect 11388 21100 16160 21128
rect 11388 21088 11394 21100
rect 10686 21020 10692 21072
rect 10744 21060 10750 21072
rect 10781 21063 10839 21069
rect 10781 21060 10793 21063
rect 10744 21032 10793 21060
rect 10744 21020 10750 21032
rect 10781 21029 10793 21032
rect 10827 21029 10839 21063
rect 13722 21060 13728 21072
rect 13683 21032 13728 21060
rect 10781 21023 10839 21029
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 13909 21063 13967 21069
rect 13909 21060 13921 21063
rect 13872 21032 13921 21060
rect 13872 21020 13878 21032
rect 13909 21029 13921 21032
rect 13955 21060 13967 21063
rect 14550 21060 14556 21072
rect 13955 21032 14556 21060
rect 13955 21029 13967 21032
rect 13909 21023 13967 21029
rect 14550 21020 14556 21032
rect 14608 21020 14614 21072
rect 14829 21063 14887 21069
rect 14829 21029 14841 21063
rect 14875 21060 14887 21063
rect 15286 21060 15292 21072
rect 14875 21032 15292 21060
rect 14875 21029 14887 21032
rect 14829 21023 14887 21029
rect 15286 21020 15292 21032
rect 15344 21020 15350 21072
rect 15488 21032 15976 21060
rect 9404 20995 9462 21001
rect 9404 20992 9416 20995
rect 8772 20964 9416 20992
rect 8294 20955 8352 20961
rect 9404 20961 9416 20964
rect 9450 20961 9462 20995
rect 9674 20992 9680 21004
rect 9635 20964 9680 20992
rect 9404 20955 9462 20961
rect 9674 20952 9680 20964
rect 9732 20952 9738 21004
rect 11698 20952 11704 21004
rect 11756 20992 11762 21004
rect 12391 20995 12449 21001
rect 12391 20992 12403 20995
rect 11756 20964 12403 20992
rect 11756 20952 11762 20964
rect 12391 20961 12403 20964
rect 12437 20961 12449 20995
rect 12391 20955 12449 20961
rect 12986 20952 12992 21004
rect 13044 20992 13050 21004
rect 13081 20995 13139 21001
rect 13081 20992 13093 20995
rect 13044 20964 13093 20992
rect 13044 20952 13050 20964
rect 13081 20961 13093 20964
rect 13127 20961 13139 20995
rect 13081 20955 13139 20961
rect 14185 20995 14243 21001
rect 14185 20961 14197 20995
rect 14231 20961 14243 20995
rect 14185 20955 14243 20961
rect 5629 20927 5687 20933
rect 5629 20893 5641 20927
rect 5675 20893 5687 20927
rect 6454 20924 6460 20936
rect 6415 20896 6460 20924
rect 5629 20887 5687 20893
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 6546 20884 6552 20936
rect 6604 20924 6610 20936
rect 6822 20924 6828 20936
rect 6604 20896 6828 20924
rect 6604 20884 6610 20896
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 8021 20927 8079 20933
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 8757 20927 8815 20933
rect 8067 20896 8708 20924
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 2409 20859 2467 20865
rect 2409 20825 2421 20859
rect 2455 20856 2467 20859
rect 2958 20856 2964 20868
rect 2455 20828 2964 20856
rect 2455 20825 2467 20828
rect 2409 20819 2467 20825
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 4617 20859 4675 20865
rect 3068 20828 4108 20856
rect 2774 20748 2780 20800
rect 2832 20788 2838 20800
rect 3068 20788 3096 20828
rect 3418 20788 3424 20800
rect 2832 20760 3096 20788
rect 3379 20760 3424 20788
rect 2832 20748 2838 20760
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 4080 20797 4108 20828
rect 4617 20825 4629 20859
rect 4663 20856 4675 20859
rect 7282 20856 7288 20868
rect 4663 20828 7288 20856
rect 4663 20825 4675 20828
rect 4617 20819 4675 20825
rect 7282 20816 7288 20828
rect 7340 20816 7346 20868
rect 8680 20856 8708 20896
rect 8757 20893 8769 20927
rect 8803 20924 8815 20927
rect 8846 20924 8852 20936
rect 8803 20896 8852 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 8846 20884 8852 20896
rect 8904 20924 8910 20936
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8904 20896 8953 20924
rect 8904 20884 8910 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 9490 20924 9496 20936
rect 8941 20887 8999 20893
rect 9048 20896 9496 20924
rect 9048 20856 9076 20896
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 9766 20884 9772 20936
rect 9824 20924 9830 20936
rect 10502 20924 10508 20936
rect 9824 20896 10508 20924
rect 9824 20884 9830 20896
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 11882 20884 11888 20936
rect 11940 20924 11946 20936
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 11940 20896 12173 20924
rect 11940 20884 11946 20896
rect 12161 20893 12173 20896
rect 12207 20893 12219 20927
rect 12894 20924 12900 20936
rect 12855 20896 12900 20924
rect 12161 20887 12219 20893
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 13262 20884 13268 20936
rect 13320 20884 13326 20936
rect 13280 20856 13308 20884
rect 8680 20828 9076 20856
rect 12820 20828 13308 20856
rect 12820 20800 12848 20828
rect 14200 20800 14228 20955
rect 14366 20952 14372 21004
rect 14424 20992 14430 21004
rect 15488 20992 15516 21032
rect 14424 20964 14469 20992
rect 15212 20964 15516 20992
rect 15565 20995 15623 21001
rect 14424 20952 14430 20964
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 15212 20924 15240 20964
rect 15565 20961 15577 20995
rect 15611 20961 15623 20995
rect 15565 20955 15623 20961
rect 15378 20924 15384 20936
rect 14516 20896 15240 20924
rect 15339 20896 15384 20924
rect 14516 20884 14522 20896
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 14550 20816 14556 20868
rect 14608 20856 14614 20868
rect 14826 20856 14832 20868
rect 14608 20828 14832 20856
rect 14608 20816 14614 20828
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 15289 20859 15347 20865
rect 15289 20825 15301 20859
rect 15335 20825 15347 20859
rect 15580 20856 15608 20955
rect 15948 20933 15976 21032
rect 16132 20933 16160 21100
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 16356 21100 19656 21128
rect 16356 21088 16362 21100
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20961 16543 20995
rect 16485 20955 16543 20961
rect 15933 20927 15991 20933
rect 15933 20893 15945 20927
rect 15979 20893 15991 20927
rect 15933 20887 15991 20893
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 16298 20856 16304 20868
rect 15580 20828 15976 20856
rect 16259 20828 16304 20856
rect 15289 20819 15347 20825
rect 4065 20791 4123 20797
rect 4065 20757 4077 20791
rect 4111 20757 4123 20791
rect 4246 20788 4252 20800
rect 4207 20760 4252 20788
rect 4065 20751 4123 20757
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 4706 20788 4712 20800
rect 4667 20760 4712 20788
rect 4706 20748 4712 20760
rect 4764 20748 4770 20800
rect 4890 20748 4896 20800
rect 4948 20788 4954 20800
rect 4985 20791 5043 20797
rect 4985 20788 4997 20791
rect 4948 20760 4997 20788
rect 4948 20748 4954 20760
rect 4985 20757 4997 20760
rect 5031 20757 5043 20791
rect 4985 20751 5043 20757
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20788 5595 20791
rect 5902 20788 5908 20800
rect 5583 20760 5908 20788
rect 5583 20757 5595 20760
rect 5537 20751 5595 20757
rect 5902 20748 5908 20760
rect 5960 20748 5966 20800
rect 6270 20748 6276 20800
rect 6328 20788 6334 20800
rect 6546 20788 6552 20800
rect 6328 20760 6552 20788
rect 6328 20748 6334 20760
rect 6546 20748 6552 20760
rect 6604 20748 6610 20800
rect 6825 20791 6883 20797
rect 6825 20757 6837 20791
rect 6871 20788 6883 20791
rect 6914 20788 6920 20800
rect 6871 20760 6920 20788
rect 6871 20757 6883 20760
rect 6825 20751 6883 20757
rect 6914 20748 6920 20760
rect 6972 20788 6978 20800
rect 7190 20788 7196 20800
rect 6972 20760 7196 20788
rect 6972 20748 6978 20760
rect 7190 20748 7196 20760
rect 7248 20748 7254 20800
rect 7650 20748 7656 20800
rect 7708 20788 7714 20800
rect 8110 20788 8116 20800
rect 7708 20760 8116 20788
rect 7708 20748 7714 20760
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 8290 20791 8348 20797
rect 8290 20757 8302 20791
rect 8336 20788 8348 20791
rect 9407 20791 9465 20797
rect 9407 20788 9419 20791
rect 8336 20760 9419 20788
rect 8336 20757 8348 20760
rect 8290 20751 8348 20757
rect 9407 20757 9419 20760
rect 9453 20788 9465 20791
rect 10410 20788 10416 20800
rect 9453 20760 10416 20788
rect 9453 20757 9465 20760
rect 9407 20751 9465 20757
rect 10410 20748 10416 20760
rect 10468 20788 10474 20800
rect 10686 20788 10692 20800
rect 10468 20760 10692 20788
rect 10468 20748 10474 20760
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 10870 20788 10876 20800
rect 10831 20760 10876 20788
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 12430 20791 12488 20797
rect 12430 20757 12442 20791
rect 12476 20788 12488 20791
rect 12526 20788 12532 20800
rect 12476 20760 12532 20788
rect 12476 20757 12488 20760
rect 12430 20751 12488 20757
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 12802 20748 12808 20800
rect 12860 20748 12866 20800
rect 13262 20788 13268 20800
rect 13223 20760 13268 20788
rect 13262 20748 13268 20760
rect 13320 20748 13326 20800
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 13412 20760 13457 20788
rect 13412 20748 13418 20760
rect 14182 20748 14188 20800
rect 14240 20748 14246 20800
rect 14461 20791 14519 20797
rect 14461 20757 14473 20791
rect 14507 20788 14519 20791
rect 14734 20788 14740 20800
rect 14507 20760 14740 20788
rect 14507 20757 14519 20760
rect 14461 20751 14519 20757
rect 14734 20748 14740 20760
rect 14792 20748 14798 20800
rect 14918 20788 14924 20800
rect 14879 20760 14924 20788
rect 14918 20748 14924 20760
rect 14976 20748 14982 20800
rect 15304 20788 15332 20819
rect 15948 20800 15976 20828
rect 16298 20816 16304 20828
rect 16356 20856 16362 20868
rect 16500 20856 16528 20955
rect 16666 20952 16672 21004
rect 16724 20992 16730 21004
rect 18325 20995 18383 21001
rect 16724 20964 17540 20992
rect 16724 20952 16730 20964
rect 16761 20927 16819 20933
rect 16761 20893 16773 20927
rect 16807 20924 16819 20927
rect 17402 20924 17408 20936
rect 16807 20896 17408 20924
rect 16807 20893 16819 20896
rect 16761 20887 16819 20893
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 17512 20924 17540 20964
rect 18325 20961 18337 20995
rect 18371 20992 18383 20995
rect 18414 20992 18420 21004
rect 18371 20964 18420 20992
rect 18371 20961 18383 20964
rect 18325 20955 18383 20961
rect 18414 20952 18420 20964
rect 18472 20952 18478 21004
rect 18598 20995 18656 21001
rect 18598 20961 18610 20995
rect 18644 20992 18656 20995
rect 19150 20992 19156 21004
rect 18644 20964 19156 20992
rect 18644 20961 18656 20964
rect 18598 20955 18656 20961
rect 19150 20952 19156 20964
rect 19208 20952 19214 21004
rect 18506 20924 18512 20936
rect 17512 20896 18512 20924
rect 18506 20884 18512 20896
rect 18564 20924 18570 20936
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 18564 20896 19073 20924
rect 18564 20884 18570 20896
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19628 20924 19656 21100
rect 19702 21088 19708 21140
rect 19760 21128 19766 21140
rect 20717 21131 20775 21137
rect 20717 21128 20729 21131
rect 19760 21100 20729 21128
rect 19760 21088 19766 21100
rect 20717 21097 20729 21100
rect 20763 21097 20775 21131
rect 20717 21091 20775 21097
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 21450 21128 21456 21140
rect 21048 21100 21456 21128
rect 21048 21088 21054 21100
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 22646 21128 22652 21140
rect 22607 21100 22652 21128
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 21545 21063 21603 21069
rect 21545 21060 21557 21063
rect 21192 21032 21557 21060
rect 20898 20952 20904 21004
rect 20956 20992 20962 21004
rect 21192 21001 21220 21032
rect 21545 21029 21557 21032
rect 21591 21029 21603 21063
rect 21545 21023 21603 21029
rect 21818 21020 21824 21072
rect 21876 21060 21882 21072
rect 21876 21032 22140 21060
rect 21876 21020 21882 21032
rect 22112 21001 22140 21032
rect 21177 20995 21235 21001
rect 21177 20992 21189 20995
rect 20956 20964 21189 20992
rect 20956 20952 20962 20964
rect 21177 20961 21189 20964
rect 21223 20961 21235 20995
rect 21177 20955 21235 20961
rect 21269 20995 21327 21001
rect 21269 20961 21281 20995
rect 21315 20961 21327 20995
rect 21269 20955 21327 20961
rect 22097 20995 22155 21001
rect 22097 20961 22109 20995
rect 22143 20961 22155 20995
rect 22097 20955 22155 20961
rect 19628 20896 20484 20924
rect 19061 20887 19119 20893
rect 16666 20856 16672 20868
rect 16356 20828 16528 20856
rect 16627 20828 16672 20856
rect 16356 20816 16362 20828
rect 16666 20816 16672 20828
rect 16724 20816 16730 20868
rect 16942 20816 16948 20868
rect 17000 20856 17006 20868
rect 17000 20828 17264 20856
rect 17000 20816 17006 20828
rect 15749 20791 15807 20797
rect 15749 20788 15761 20791
rect 15304 20760 15761 20788
rect 15749 20757 15761 20760
rect 15795 20757 15807 20791
rect 15749 20751 15807 20757
rect 15930 20748 15936 20800
rect 15988 20748 15994 20800
rect 17126 20788 17132 20800
rect 17087 20760 17132 20788
rect 17126 20748 17132 20760
rect 17184 20748 17190 20800
rect 17236 20797 17264 20828
rect 20254 20816 20260 20868
rect 20312 20856 20318 20868
rect 20358 20859 20416 20865
rect 20358 20856 20370 20859
rect 20312 20828 20370 20856
rect 20312 20816 20318 20828
rect 20358 20825 20370 20828
rect 20404 20825 20416 20859
rect 20456 20856 20484 20896
rect 20530 20884 20536 20936
rect 20588 20924 20594 20936
rect 20625 20927 20683 20933
rect 20625 20924 20637 20927
rect 20588 20896 20637 20924
rect 20588 20884 20594 20896
rect 20625 20893 20637 20896
rect 20671 20893 20683 20927
rect 20625 20887 20683 20893
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 21284 20924 21312 20955
rect 21048 20896 21312 20924
rect 21048 20884 21054 20896
rect 22278 20884 22284 20936
rect 22336 20924 22342 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22336 20896 22477 20924
rect 22336 20884 22342 20896
rect 22465 20893 22477 20896
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20924 22891 20927
rect 23658 20924 23664 20936
rect 22879 20896 23664 20924
rect 22879 20893 22891 20896
rect 22833 20887 22891 20893
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 22186 20856 22192 20868
rect 20456 20828 22192 20856
rect 20358 20819 20416 20825
rect 22186 20816 22192 20828
rect 22244 20816 22250 20868
rect 17221 20791 17279 20797
rect 17221 20757 17233 20791
rect 17267 20757 17279 20791
rect 17221 20751 17279 20757
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 18594 20791 18652 20797
rect 18594 20788 18606 20791
rect 18380 20760 18606 20788
rect 18380 20748 18386 20760
rect 18594 20757 18606 20760
rect 18640 20757 18652 20791
rect 19242 20788 19248 20800
rect 19203 20760 19248 20788
rect 18594 20751 18652 20757
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 19886 20748 19892 20800
rect 19944 20788 19950 20800
rect 21085 20791 21143 20797
rect 21085 20788 21097 20791
rect 19944 20760 21097 20788
rect 19944 20748 19950 20760
rect 21085 20757 21097 20760
rect 21131 20757 21143 20791
rect 21085 20751 21143 20757
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21913 20791 21971 20797
rect 21913 20788 21925 20791
rect 21232 20760 21925 20788
rect 21232 20748 21238 20760
rect 21913 20757 21925 20760
rect 21959 20757 21971 20791
rect 21913 20751 21971 20757
rect 22002 20748 22008 20800
rect 22060 20788 22066 20800
rect 23014 20788 23020 20800
rect 22060 20760 22105 20788
rect 22975 20760 23020 20788
rect 22060 20748 22066 20760
rect 23014 20748 23020 20760
rect 23072 20748 23078 20800
rect 1104 20698 23460 20720
rect 1104 20646 6548 20698
rect 6600 20646 6612 20698
rect 6664 20646 6676 20698
rect 6728 20646 6740 20698
rect 6792 20646 6804 20698
rect 6856 20646 12146 20698
rect 12198 20646 12210 20698
rect 12262 20646 12274 20698
rect 12326 20646 12338 20698
rect 12390 20646 12402 20698
rect 12454 20646 17744 20698
rect 17796 20646 17808 20698
rect 17860 20646 17872 20698
rect 17924 20646 17936 20698
rect 17988 20646 18000 20698
rect 18052 20646 23460 20698
rect 1104 20624 23460 20646
rect 2314 20544 2320 20596
rect 2372 20584 2378 20596
rect 2409 20587 2467 20593
rect 2409 20584 2421 20587
rect 2372 20556 2421 20584
rect 2372 20544 2378 20556
rect 2409 20553 2421 20556
rect 2455 20553 2467 20587
rect 2866 20584 2872 20596
rect 2827 20556 2872 20584
rect 2409 20547 2467 20553
rect 2866 20544 2872 20556
rect 2924 20544 2930 20596
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 3510 20584 3516 20596
rect 3099 20556 3516 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3510 20544 3516 20556
rect 3568 20544 3574 20596
rect 3973 20587 4031 20593
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 4338 20584 4344 20596
rect 4019 20556 4344 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 4338 20544 4344 20556
rect 4396 20544 4402 20596
rect 5077 20587 5135 20593
rect 5077 20553 5089 20587
rect 5123 20553 5135 20587
rect 5077 20547 5135 20553
rect 3237 20519 3295 20525
rect 3237 20485 3249 20519
rect 3283 20516 3295 20519
rect 4614 20516 4620 20528
rect 3283 20488 4620 20516
rect 3283 20485 3295 20488
rect 3237 20479 3295 20485
rect 4614 20476 4620 20488
rect 4672 20476 4678 20528
rect 5092 20516 5120 20547
rect 5626 20544 5632 20596
rect 5684 20584 5690 20596
rect 5997 20587 6055 20593
rect 5997 20584 6009 20587
rect 5684 20556 6009 20584
rect 5684 20544 5690 20556
rect 5997 20553 6009 20556
rect 6043 20553 6055 20587
rect 5997 20547 6055 20553
rect 6730 20544 6736 20596
rect 6788 20584 6794 20596
rect 8113 20587 8171 20593
rect 6788 20556 8064 20584
rect 6788 20544 6794 20556
rect 5718 20516 5724 20528
rect 5092 20488 5724 20516
rect 5718 20476 5724 20488
rect 5776 20476 5782 20528
rect 5810 20476 5816 20528
rect 5868 20516 5874 20528
rect 8036 20516 8064 20556
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8662 20584 8668 20596
rect 8159 20556 8668 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 8941 20587 8999 20593
rect 8941 20553 8953 20587
rect 8987 20584 8999 20587
rect 9490 20584 9496 20596
rect 8987 20556 9352 20584
rect 9451 20556 9496 20584
rect 8987 20553 8999 20556
rect 8941 20547 8999 20553
rect 9324 20516 9352 20556
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 9953 20587 10011 20593
rect 9953 20553 9965 20587
rect 9999 20584 10011 20587
rect 10594 20584 10600 20596
rect 9999 20556 10600 20584
rect 9999 20553 10011 20556
rect 9953 20547 10011 20553
rect 10594 20544 10600 20556
rect 10652 20544 10658 20596
rect 11333 20587 11391 20593
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 13354 20584 13360 20596
rect 11379 20556 13360 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 13449 20587 13507 20593
rect 13449 20553 13461 20587
rect 13495 20553 13507 20587
rect 13449 20547 13507 20553
rect 13909 20587 13967 20593
rect 13909 20553 13921 20587
rect 13955 20584 13967 20587
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 13955 20556 14289 20584
rect 13955 20553 13967 20556
rect 13909 20547 13967 20553
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 15933 20587 15991 20593
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 18138 20584 18144 20596
rect 15979 20556 18144 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 9401 20519 9459 20525
rect 9401 20516 9413 20519
rect 5868 20488 7788 20516
rect 8036 20488 9168 20516
rect 9324 20488 9413 20516
rect 5868 20476 5874 20488
rect 3326 20408 3332 20460
rect 3384 20448 3390 20460
rect 3881 20451 3939 20457
rect 3881 20448 3893 20451
rect 3384 20420 3893 20448
rect 3384 20408 3390 20420
rect 3881 20417 3893 20420
rect 3927 20417 3939 20451
rect 3881 20411 3939 20417
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 4709 20451 4767 20457
rect 4709 20448 4721 20451
rect 4212 20420 4721 20448
rect 4212 20408 4218 20420
rect 4709 20417 4721 20420
rect 4755 20417 4767 20451
rect 4709 20411 4767 20417
rect 5629 20451 5687 20457
rect 5629 20417 5641 20451
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20380 3479 20383
rect 3786 20380 3792 20392
rect 3467 20352 3792 20380
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20349 4123 20383
rect 4065 20343 4123 20349
rect 4080 20312 4108 20343
rect 4430 20340 4436 20392
rect 4488 20380 4494 20392
rect 4614 20380 4620 20392
rect 4488 20352 4533 20380
rect 4575 20352 4620 20380
rect 4488 20340 4494 20352
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 4798 20312 4804 20324
rect 3436 20284 3924 20312
rect 4080 20284 4804 20312
rect 3436 20256 3464 20284
rect 3418 20204 3424 20256
rect 3476 20204 3482 20256
rect 3513 20247 3571 20253
rect 3513 20213 3525 20247
rect 3559 20244 3571 20247
rect 3602 20244 3608 20256
rect 3559 20216 3608 20244
rect 3559 20213 3571 20216
rect 3513 20207 3571 20213
rect 3602 20204 3608 20216
rect 3660 20204 3666 20256
rect 3896 20244 3924 20284
rect 4798 20272 4804 20284
rect 4856 20312 4862 20324
rect 5445 20315 5503 20321
rect 5445 20312 5457 20315
rect 4856 20284 5457 20312
rect 4856 20272 4862 20284
rect 5445 20281 5457 20284
rect 5491 20281 5503 20315
rect 5644 20312 5672 20411
rect 5994 20408 6000 20460
rect 6052 20448 6058 20460
rect 7760 20457 7788 20488
rect 7478 20451 7536 20457
rect 7478 20448 7490 20451
rect 6052 20420 7490 20448
rect 6052 20408 6058 20420
rect 7478 20417 7490 20420
rect 7524 20417 7536 20451
rect 7478 20411 7536 20417
rect 7745 20451 7803 20457
rect 7745 20417 7757 20451
rect 7791 20417 7803 20451
rect 8570 20448 8576 20460
rect 8531 20420 8576 20448
rect 7745 20411 7803 20417
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 9140 20448 9168 20488
rect 9401 20485 9413 20488
rect 9447 20516 9459 20519
rect 9766 20516 9772 20528
rect 9447 20488 9772 20516
rect 9447 20485 9459 20488
rect 9401 20479 9459 20485
rect 9766 20476 9772 20488
rect 9824 20476 9830 20528
rect 11146 20516 11152 20528
rect 10244 20488 11152 20516
rect 10244 20457 10272 20488
rect 11146 20476 11152 20488
rect 11204 20476 11210 20528
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 9140 20420 10241 20448
rect 10229 20417 10241 20420
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 10689 20451 10747 20457
rect 10689 20448 10701 20451
rect 10376 20420 10701 20448
rect 10376 20408 10382 20420
rect 10689 20417 10701 20420
rect 10735 20417 10747 20451
rect 10689 20411 10747 20417
rect 10778 20408 10784 20460
rect 10836 20448 10842 20460
rect 11840 20451 11898 20457
rect 11840 20448 11852 20451
rect 10836 20420 11852 20448
rect 10836 20408 10842 20420
rect 11840 20417 11852 20420
rect 11886 20417 11898 20451
rect 13464 20448 13492 20547
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 18874 20584 18880 20596
rect 18564 20556 18880 20584
rect 18564 20544 18570 20556
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 19150 20544 19156 20596
rect 19208 20584 19214 20596
rect 20165 20587 20223 20593
rect 20165 20584 20177 20587
rect 19208 20556 20177 20584
rect 19208 20544 19214 20556
rect 20165 20553 20177 20556
rect 20211 20584 20223 20587
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 20211 20556 21465 20584
rect 20211 20553 20223 20556
rect 20165 20547 20223 20553
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 21821 20587 21879 20593
rect 21821 20584 21833 20587
rect 21600 20556 21833 20584
rect 21600 20544 21606 20556
rect 21821 20553 21833 20556
rect 21867 20553 21879 20587
rect 21821 20547 21879 20553
rect 22281 20587 22339 20593
rect 22281 20553 22293 20587
rect 22327 20584 22339 20587
rect 22370 20584 22376 20596
rect 22327 20556 22376 20584
rect 22327 20553 22339 20556
rect 22281 20547 22339 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 14645 20519 14703 20525
rect 14645 20516 14657 20519
rect 11840 20411 11898 20417
rect 12176 20420 13492 20448
rect 13556 20488 14657 20516
rect 5905 20383 5963 20389
rect 5905 20349 5917 20383
rect 5951 20380 5963 20383
rect 6730 20380 6736 20392
rect 5951 20352 6736 20380
rect 5951 20349 5963 20352
rect 5905 20343 5963 20349
rect 6730 20340 6736 20352
rect 6788 20340 6794 20392
rect 8294 20380 8300 20392
rect 8255 20352 8300 20380
rect 8294 20340 8300 20352
rect 8352 20340 8358 20392
rect 8481 20383 8539 20389
rect 8481 20349 8493 20383
rect 8527 20380 8539 20383
rect 8662 20380 8668 20392
rect 8527 20352 8668 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 8662 20340 8668 20352
rect 8720 20340 8726 20392
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 5644 20284 6500 20312
rect 5445 20275 5503 20281
rect 4430 20244 4436 20256
rect 3896 20216 4436 20244
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 5353 20247 5411 20253
rect 5353 20213 5365 20247
rect 5399 20244 5411 20247
rect 5810 20244 5816 20256
rect 5399 20216 5816 20244
rect 5399 20213 5411 20216
rect 5353 20207 5411 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 6086 20204 6092 20256
rect 6144 20244 6150 20256
rect 6365 20247 6423 20253
rect 6365 20244 6377 20247
rect 6144 20216 6377 20244
rect 6144 20204 6150 20216
rect 6365 20213 6377 20216
rect 6411 20213 6423 20247
rect 6472 20244 6500 20284
rect 8938 20272 8944 20324
rect 8996 20312 9002 20324
rect 9033 20315 9091 20321
rect 9033 20312 9045 20315
rect 8996 20284 9045 20312
rect 8996 20272 9002 20284
rect 9033 20281 9045 20284
rect 9079 20281 9091 20315
rect 9033 20275 9091 20281
rect 9214 20272 9220 20324
rect 9272 20312 9278 20324
rect 9600 20312 9628 20343
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 10413 20383 10471 20389
rect 10413 20380 10425 20383
rect 9732 20352 10425 20380
rect 9732 20340 9738 20352
rect 10413 20349 10425 20352
rect 10459 20349 10471 20383
rect 10413 20343 10471 20349
rect 10597 20383 10655 20389
rect 10597 20349 10609 20383
rect 10643 20380 10655 20383
rect 11054 20380 11060 20392
rect 10643 20352 11060 20380
rect 10643 20349 10655 20352
rect 10597 20343 10655 20349
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 11517 20383 11575 20389
rect 11517 20380 11529 20383
rect 11204 20352 11529 20380
rect 11204 20340 11210 20352
rect 11517 20349 11529 20352
rect 11563 20349 11575 20383
rect 11517 20343 11575 20349
rect 12023 20383 12081 20389
rect 12023 20349 12035 20383
rect 12069 20380 12081 20383
rect 12176 20380 12204 20420
rect 12069 20352 12204 20380
rect 12069 20349 12081 20352
rect 12023 20343 12081 20349
rect 12250 20340 12256 20392
rect 12308 20380 12314 20392
rect 13556 20380 13584 20488
rect 14645 20485 14657 20488
rect 14691 20485 14703 20519
rect 14645 20479 14703 20485
rect 14936 20488 16252 20516
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20448 13875 20451
rect 14090 20448 14096 20460
rect 13863 20420 14096 20448
rect 13863 20417 13875 20420
rect 13817 20411 13875 20417
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 12308 20352 13584 20380
rect 14001 20383 14059 20389
rect 12308 20340 12314 20352
rect 14001 20349 14013 20383
rect 14047 20349 14059 20383
rect 14734 20380 14740 20392
rect 14695 20352 14740 20380
rect 14001 20343 14059 20349
rect 9272 20284 9628 20312
rect 13357 20315 13415 20321
rect 9272 20272 9278 20284
rect 13357 20281 13369 20315
rect 13403 20312 13415 20315
rect 13446 20312 13452 20324
rect 13403 20284 13452 20312
rect 13403 20281 13415 20284
rect 13357 20275 13415 20281
rect 13446 20272 13452 20284
rect 13504 20272 13510 20324
rect 14016 20312 14044 20343
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 14936 20389 14964 20488
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 16022 20448 16028 20460
rect 15611 20420 16028 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 14921 20383 14979 20389
rect 14921 20349 14933 20383
rect 14967 20349 14979 20383
rect 15286 20380 15292 20392
rect 15247 20352 15292 20380
rect 14921 20343 14979 20349
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 15470 20380 15476 20392
rect 15431 20352 15476 20380
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 16224 20380 16252 20488
rect 16408 20488 17264 20516
rect 16408 20460 16436 20488
rect 16390 20448 16396 20460
rect 16351 20420 16396 20448
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 17034 20448 17040 20460
rect 16995 20420 17040 20448
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 16666 20380 16672 20392
rect 16224 20352 16672 20380
rect 16666 20340 16672 20352
rect 16724 20340 16730 20392
rect 16942 20340 16948 20392
rect 17000 20380 17006 20392
rect 17236 20389 17264 20488
rect 17494 20476 17500 20528
rect 17552 20516 17558 20528
rect 17862 20516 17868 20528
rect 17552 20488 17868 20516
rect 17552 20476 17558 20488
rect 17862 20476 17868 20488
rect 17920 20476 17926 20528
rect 18592 20519 18650 20525
rect 18592 20485 18604 20519
rect 18638 20516 18650 20519
rect 19242 20516 19248 20528
rect 18638 20488 19248 20516
rect 18638 20485 18650 20488
rect 18592 20479 18650 20485
rect 19242 20476 19248 20488
rect 19300 20516 19306 20528
rect 20901 20519 20959 20525
rect 20901 20516 20913 20519
rect 19300 20488 20913 20516
rect 19300 20476 19306 20488
rect 20901 20485 20913 20488
rect 20947 20485 20959 20519
rect 20901 20479 20959 20485
rect 19058 20408 19064 20460
rect 19116 20448 19122 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 19116 20420 20085 20448
rect 19116 20408 19122 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20073 20411 20131 20417
rect 20456 20420 21005 20448
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 17000 20352 17141 20380
rect 17000 20340 17006 20352
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 17221 20383 17279 20389
rect 17221 20349 17233 20383
rect 17267 20349 17279 20383
rect 17402 20380 17408 20392
rect 17221 20343 17279 20349
rect 17328 20352 17408 20380
rect 14826 20312 14832 20324
rect 14016 20284 14832 20312
rect 14826 20272 14832 20284
rect 14884 20272 14890 20324
rect 15654 20272 15660 20324
rect 15712 20312 15718 20324
rect 16209 20315 16267 20321
rect 16209 20312 16221 20315
rect 15712 20284 16221 20312
rect 15712 20272 15718 20284
rect 16209 20281 16221 20284
rect 16255 20281 16267 20315
rect 16209 20275 16267 20281
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 6472 20216 10057 20244
rect 6365 20207 6423 20213
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 11057 20247 11115 20253
rect 11057 20213 11069 20247
rect 11103 20244 11115 20247
rect 13262 20244 13268 20256
rect 11103 20216 13268 20244
rect 11103 20213 11115 20216
rect 11057 20207 11115 20213
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 14918 20244 14924 20256
rect 13596 20216 14924 20244
rect 13596 20204 13602 20216
rect 14918 20204 14924 20216
rect 14976 20204 14982 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 16025 20247 16083 20253
rect 16025 20244 16037 20247
rect 15620 20216 16037 20244
rect 15620 20204 15626 20216
rect 16025 20213 16037 20216
rect 16071 20213 16083 20247
rect 16025 20207 16083 20213
rect 16669 20247 16727 20253
rect 16669 20213 16681 20247
rect 16715 20244 16727 20247
rect 17328 20244 17356 20352
rect 17402 20340 17408 20352
rect 17460 20340 17466 20392
rect 17954 20380 17960 20392
rect 17915 20352 17960 20380
rect 17954 20340 17960 20352
rect 18012 20340 18018 20392
rect 18138 20380 18144 20392
rect 18099 20352 18144 20380
rect 18138 20340 18144 20352
rect 18196 20340 18202 20392
rect 18325 20383 18383 20389
rect 18325 20349 18337 20383
rect 18371 20349 18383 20383
rect 19886 20380 19892 20392
rect 19847 20352 19892 20380
rect 18325 20343 18383 20349
rect 16715 20216 17356 20244
rect 16715 20213 16727 20216
rect 16669 20207 16727 20213
rect 17402 20204 17408 20256
rect 17460 20244 17466 20256
rect 17497 20247 17555 20253
rect 17497 20244 17509 20247
rect 17460 20216 17509 20244
rect 17460 20204 17466 20216
rect 17497 20213 17509 20216
rect 17543 20213 17555 20247
rect 18340 20244 18368 20343
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 19705 20315 19763 20321
rect 19705 20281 19717 20315
rect 19751 20312 19763 20315
rect 20456 20312 20484 20420
rect 20916 20392 20944 20420
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 21358 20408 21364 20460
rect 21416 20448 21422 20460
rect 21637 20451 21695 20457
rect 21637 20448 21649 20451
rect 21416 20420 21649 20448
rect 21416 20408 21422 20420
rect 21637 20417 21649 20420
rect 21683 20417 21695 20451
rect 21637 20411 21695 20417
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20448 22155 20451
rect 22186 20448 22192 20460
rect 22143 20420 22192 20448
rect 22143 20417 22155 20420
rect 22097 20411 22155 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 22465 20451 22523 20457
rect 22465 20417 22477 20451
rect 22511 20417 22523 20451
rect 22465 20411 22523 20417
rect 22833 20451 22891 20457
rect 22833 20417 22845 20451
rect 22879 20448 22891 20451
rect 22922 20448 22928 20460
rect 22879 20420 22928 20448
rect 22879 20417 22891 20420
rect 22833 20411 22891 20417
rect 20809 20383 20867 20389
rect 20809 20349 20821 20383
rect 20855 20349 20867 20383
rect 20809 20343 20867 20349
rect 19751 20284 20484 20312
rect 20533 20315 20591 20321
rect 19751 20281 19763 20284
rect 19705 20275 19763 20281
rect 20533 20281 20545 20315
rect 20579 20312 20591 20315
rect 20622 20312 20628 20324
rect 20579 20284 20628 20312
rect 20579 20281 20591 20284
rect 20533 20275 20591 20281
rect 20622 20272 20628 20284
rect 20680 20272 20686 20324
rect 20824 20312 20852 20343
rect 20898 20340 20904 20392
rect 20956 20340 20962 20392
rect 22480 20380 22508 20411
rect 22922 20408 22928 20420
rect 22980 20408 22986 20460
rect 23566 20380 23572 20392
rect 22480 20352 23572 20380
rect 23566 20340 23572 20352
rect 23624 20340 23630 20392
rect 22649 20315 22707 20321
rect 20824 20284 20944 20312
rect 19334 20244 19340 20256
rect 18340 20216 19340 20244
rect 17497 20207 17555 20213
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 20916 20244 20944 20284
rect 22649 20281 22661 20315
rect 22695 20312 22707 20315
rect 23106 20312 23112 20324
rect 22695 20284 23112 20312
rect 22695 20281 22707 20284
rect 22649 20275 22707 20281
rect 23106 20272 23112 20284
rect 23164 20272 23170 20324
rect 21082 20244 21088 20256
rect 20916 20216 21088 20244
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21358 20244 21364 20256
rect 21319 20216 21364 20244
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 23017 20247 23075 20253
rect 23017 20213 23029 20247
rect 23063 20244 23075 20247
rect 23290 20244 23296 20256
rect 23063 20216 23296 20244
rect 23063 20213 23075 20216
rect 23017 20207 23075 20213
rect 23290 20204 23296 20216
rect 23348 20204 23354 20256
rect 1104 20154 23460 20176
rect 1104 20102 3749 20154
rect 3801 20102 3813 20154
rect 3865 20102 3877 20154
rect 3929 20102 3941 20154
rect 3993 20102 4005 20154
rect 4057 20102 9347 20154
rect 9399 20102 9411 20154
rect 9463 20102 9475 20154
rect 9527 20102 9539 20154
rect 9591 20102 9603 20154
rect 9655 20102 14945 20154
rect 14997 20102 15009 20154
rect 15061 20102 15073 20154
rect 15125 20102 15137 20154
rect 15189 20102 15201 20154
rect 15253 20102 20543 20154
rect 20595 20102 20607 20154
rect 20659 20102 20671 20154
rect 20723 20102 20735 20154
rect 20787 20102 20799 20154
rect 20851 20102 23460 20154
rect 1104 20080 23460 20102
rect 4154 20040 4160 20052
rect 4115 20012 4160 20040
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 4338 20040 4344 20052
rect 4299 20012 4344 20040
rect 4338 20000 4344 20012
rect 4396 20000 4402 20052
rect 5074 20040 5080 20052
rect 4908 20012 5080 20040
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19904 4859 19907
rect 4908 19904 4936 20012
rect 5074 20000 5080 20012
rect 5132 20040 5138 20052
rect 5994 20040 6000 20052
rect 5132 20012 6000 20040
rect 5132 20000 5138 20012
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6178 20000 6184 20052
rect 6236 20040 6242 20052
rect 8386 20040 8392 20052
rect 6236 20012 8392 20040
rect 6236 20000 6242 20012
rect 8386 20000 8392 20012
rect 8444 20040 8450 20052
rect 8573 20043 8631 20049
rect 8573 20040 8585 20043
rect 8444 20012 8585 20040
rect 8444 20000 8450 20012
rect 8573 20009 8585 20012
rect 8619 20009 8631 20043
rect 8573 20003 8631 20009
rect 10226 20000 10232 20052
rect 10284 20040 10290 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10284 20012 10333 20040
rect 10284 20000 10290 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10321 20003 10379 20009
rect 12437 20043 12495 20049
rect 12437 20009 12449 20043
rect 12483 20040 12495 20043
rect 12802 20040 12808 20052
rect 12483 20012 12808 20040
rect 12483 20009 12495 20012
rect 12437 20003 12495 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13354 20040 13360 20052
rect 13136 20012 13360 20040
rect 13136 20000 13142 20012
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 13909 20043 13967 20049
rect 13909 20009 13921 20043
rect 13955 20040 13967 20043
rect 14734 20040 14740 20052
rect 13955 20012 14740 20040
rect 13955 20009 13967 20012
rect 13909 20003 13967 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 15252 20012 15976 20040
rect 15252 20000 15258 20012
rect 5350 19972 5356 19984
rect 5000 19944 5356 19972
rect 5000 19913 5028 19944
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 12066 19932 12072 19984
rect 12124 19972 12130 19984
rect 14182 19972 14188 19984
rect 12124 19944 14188 19972
rect 12124 19932 12130 19944
rect 14182 19932 14188 19944
rect 14240 19932 14246 19984
rect 4847 19876 4936 19904
rect 4985 19907 5043 19913
rect 4847 19873 4859 19876
rect 4801 19867 4859 19873
rect 4985 19873 4997 19907
rect 5031 19873 5043 19907
rect 6086 19904 6092 19916
rect 4985 19867 5043 19873
rect 5184 19876 6092 19904
rect 3602 19836 3608 19848
rect 3563 19808 3608 19836
rect 3602 19796 3608 19808
rect 3660 19796 3666 19848
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19836 4031 19839
rect 4338 19836 4344 19848
rect 4019 19808 4344 19836
rect 4019 19805 4031 19808
rect 3973 19799 4031 19805
rect 4338 19796 4344 19808
rect 4396 19796 4402 19848
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 5184 19836 5212 19876
rect 6086 19864 6092 19876
rect 6144 19864 6150 19916
rect 12158 19864 12164 19916
rect 12216 19904 12222 19916
rect 12529 19907 12587 19913
rect 12529 19904 12541 19907
rect 12216 19876 12541 19904
rect 12216 19864 12222 19876
rect 12529 19873 12541 19876
rect 12575 19873 12587 19907
rect 12529 19867 12587 19873
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 13265 19907 13323 19913
rect 13265 19904 13277 19907
rect 12860 19876 13277 19904
rect 12860 19864 12866 19876
rect 13265 19873 13277 19876
rect 13311 19873 13323 19907
rect 13265 19867 13323 19873
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 13538 19904 13544 19916
rect 13495 19876 13544 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 14090 19904 14096 19916
rect 14051 19876 14096 19904
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 15948 19904 15976 20012
rect 17678 20000 17684 20052
rect 17736 20040 17742 20052
rect 19058 20040 19064 20052
rect 17736 20012 19064 20040
rect 17736 20000 17742 20012
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 20806 20000 20812 20052
rect 20864 20040 20870 20052
rect 21266 20040 21272 20052
rect 20864 20012 21272 20040
rect 20864 20000 20870 20012
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 21821 20043 21879 20049
rect 21821 20009 21833 20043
rect 21867 20040 21879 20043
rect 23474 20040 23480 20052
rect 21867 20012 23480 20040
rect 21867 20009 21879 20012
rect 21821 20003 21879 20009
rect 23474 20000 23480 20012
rect 23532 20000 23538 20052
rect 16209 19975 16267 19981
rect 16209 19941 16221 19975
rect 16255 19972 16267 19975
rect 17494 19972 17500 19984
rect 16255 19944 17500 19972
rect 16255 19941 16267 19944
rect 16209 19935 16267 19941
rect 17494 19932 17500 19944
rect 17552 19932 17558 19984
rect 21082 19972 21088 19984
rect 20916 19944 21088 19972
rect 16298 19904 16304 19916
rect 15948 19876 16304 19904
rect 16298 19864 16304 19876
rect 16356 19904 16362 19916
rect 16393 19907 16451 19913
rect 16393 19904 16405 19907
rect 16356 19876 16405 19904
rect 16356 19864 16362 19876
rect 16393 19873 16405 19876
rect 16439 19873 16451 19907
rect 16393 19867 16451 19873
rect 16758 19864 16764 19916
rect 16816 19864 16822 19916
rect 17310 19904 17316 19916
rect 17271 19876 17316 19904
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 20916 19913 20944 19944
rect 21082 19932 21088 19944
rect 21140 19972 21146 19984
rect 22738 19972 22744 19984
rect 21140 19944 22744 19972
rect 21140 19932 21146 19944
rect 22738 19932 22744 19944
rect 22796 19932 22802 19984
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 22094 19864 22100 19916
rect 22152 19904 22158 19916
rect 22152 19876 22197 19904
rect 22152 19864 22158 19876
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 4755 19808 5212 19836
rect 5276 19808 5549 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 5276 19768 5304 19808
rect 5537 19805 5549 19808
rect 5583 19836 5595 19839
rect 5810 19836 5816 19848
rect 5583 19808 5816 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 5810 19796 5816 19808
rect 5868 19836 5874 19848
rect 7101 19839 7159 19845
rect 7101 19836 7113 19839
rect 5868 19808 7113 19836
rect 5868 19796 5874 19808
rect 7101 19805 7113 19808
rect 7147 19836 7159 19839
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 7147 19808 7205 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 7193 19805 7205 19808
rect 7239 19836 7251 19839
rect 8665 19839 8723 19845
rect 8665 19836 8677 19839
rect 7239 19808 8677 19836
rect 7239 19805 7251 19808
rect 7193 19799 7251 19805
rect 8665 19805 8677 19808
rect 8711 19836 8723 19839
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 8711 19808 8953 19836
rect 8711 19805 8723 19808
rect 8665 19799 8723 19805
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 10594 19836 10600 19848
rect 10555 19808 10600 19836
rect 8941 19799 8999 19805
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 10870 19796 10876 19848
rect 10928 19836 10934 19848
rect 12069 19839 12127 19845
rect 12069 19836 12081 19839
rect 10928 19808 12081 19836
rect 10928 19796 10934 19808
rect 12069 19805 12081 19808
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 12710 19836 12716 19848
rect 12299 19808 12716 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 13170 19836 13176 19848
rect 12943 19808 13176 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 13354 19796 13360 19848
rect 13412 19836 13418 19848
rect 14829 19839 14887 19845
rect 13412 19808 14780 19836
rect 13412 19796 13418 19808
rect 3804 19740 5304 19768
rect 3050 19660 3056 19712
rect 3108 19700 3114 19712
rect 3421 19703 3479 19709
rect 3421 19700 3433 19703
rect 3108 19672 3433 19700
rect 3108 19660 3114 19672
rect 3421 19669 3433 19672
rect 3467 19669 3479 19703
rect 3421 19663 3479 19669
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 3804 19709 3832 19740
rect 5350 19728 5356 19780
rect 5408 19768 5414 19780
rect 5408 19740 5453 19768
rect 5408 19728 5414 19740
rect 6086 19728 6092 19780
rect 6144 19768 6150 19780
rect 6834 19771 6892 19777
rect 6834 19768 6846 19771
rect 6144 19740 6846 19768
rect 6144 19728 6150 19740
rect 6834 19737 6846 19740
rect 6880 19737 6892 19771
rect 6834 19731 6892 19737
rect 7282 19728 7288 19780
rect 7340 19768 7346 19780
rect 7438 19771 7496 19777
rect 7438 19768 7450 19771
rect 7340 19740 7450 19768
rect 7340 19728 7346 19740
rect 7438 19737 7450 19740
rect 7484 19768 7496 19771
rect 7558 19768 7564 19780
rect 7484 19740 7564 19768
rect 7484 19737 7496 19740
rect 7438 19731 7496 19737
rect 7558 19728 7564 19740
rect 7616 19728 7622 19780
rect 8754 19728 8760 19780
rect 8812 19768 8818 19780
rect 9214 19777 9220 19780
rect 9186 19771 9220 19777
rect 9186 19768 9198 19771
rect 8812 19740 9198 19768
rect 8812 19728 8818 19740
rect 9186 19737 9198 19740
rect 9272 19768 9278 19780
rect 11146 19768 11152 19780
rect 9272 19740 9334 19768
rect 9416 19740 11152 19768
rect 9186 19731 9220 19737
rect 9214 19728 9220 19731
rect 9272 19728 9278 19740
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3568 19672 3801 19700
rect 3568 19660 3574 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 5258 19700 5264 19712
rect 5219 19672 5264 19700
rect 3789 19663 3847 19669
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 5718 19700 5724 19712
rect 5679 19672 5724 19700
rect 5718 19660 5724 19672
rect 5776 19660 5782 19712
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 9416 19700 9444 19740
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 11824 19771 11882 19777
rect 11824 19737 11836 19771
rect 11870 19768 11882 19771
rect 11974 19768 11980 19780
rect 11870 19740 11980 19768
rect 11870 19737 11882 19740
rect 11824 19731 11882 19737
rect 11974 19728 11980 19740
rect 12032 19728 12038 19780
rect 13541 19771 13599 19777
rect 13541 19737 13553 19771
rect 13587 19768 13599 19771
rect 14369 19771 14427 19777
rect 14369 19768 14381 19771
rect 13587 19740 14381 19768
rect 13587 19737 13599 19740
rect 13541 19731 13599 19737
rect 14369 19737 14381 19740
rect 14415 19737 14427 19771
rect 14369 19731 14427 19737
rect 8904 19672 9444 19700
rect 8904 19660 8910 19672
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 10686 19700 10692 19712
rect 10468 19672 10513 19700
rect 10647 19672 10692 19700
rect 10468 19660 10474 19672
rect 10686 19660 10692 19672
rect 10744 19660 10750 19712
rect 13078 19700 13084 19712
rect 13039 19672 13084 19700
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 13170 19660 13176 19712
rect 13228 19700 13234 19712
rect 14645 19703 14703 19709
rect 14645 19700 14657 19703
rect 13228 19672 14657 19700
rect 13228 19660 13234 19672
rect 14645 19669 14657 19672
rect 14691 19669 14703 19703
rect 14752 19700 14780 19808
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 15562 19836 15568 19848
rect 14875 19808 15568 19836
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 15930 19836 15936 19848
rect 15712 19808 15936 19836
rect 15712 19796 15718 19808
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 15096 19771 15154 19777
rect 15096 19737 15108 19771
rect 15142 19768 15154 19771
rect 15286 19768 15292 19780
rect 15142 19740 15292 19768
rect 15142 19737 15154 19740
rect 15096 19731 15154 19737
rect 15286 19728 15292 19740
rect 15344 19768 15350 19780
rect 16482 19768 16488 19780
rect 15344 19740 16488 19768
rect 15344 19728 15350 19740
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 16776 19768 16804 19864
rect 17402 19836 17408 19848
rect 17363 19808 17408 19836
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 17727 19808 19257 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 19245 19805 19257 19808
rect 19291 19836 19303 19839
rect 19334 19836 19340 19848
rect 19291 19808 19340 19836
rect 19291 19805 19303 19808
rect 19245 19799 19303 19805
rect 19334 19796 19340 19808
rect 19392 19836 19398 19848
rect 20438 19836 20444 19848
rect 19392 19808 20444 19836
rect 19392 19796 19398 19808
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 20993 19839 21051 19845
rect 20993 19836 21005 19839
rect 20772 19808 21005 19836
rect 20772 19796 20778 19808
rect 20993 19805 21005 19808
rect 21039 19805 21051 19839
rect 20993 19799 21051 19805
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 21637 19839 21695 19845
rect 21637 19836 21649 19839
rect 21508 19808 21649 19836
rect 21508 19796 21514 19808
rect 21637 19805 21649 19808
rect 21683 19805 21695 19839
rect 22830 19836 22836 19848
rect 22791 19808 22836 19836
rect 21637 19799 21695 19805
rect 22830 19796 22836 19808
rect 22888 19796 22894 19848
rect 17954 19777 17960 19780
rect 17948 19768 17960 19777
rect 16776 19740 17356 19768
rect 17915 19740 17960 19768
rect 15930 19700 15936 19712
rect 14752 19672 15936 19700
rect 14645 19663 14703 19669
rect 15930 19660 15936 19672
rect 15988 19660 15994 19712
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16298 19700 16304 19712
rect 16080 19672 16304 19700
rect 16080 19660 16086 19672
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 16574 19700 16580 19712
rect 16535 19672 16580 19700
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19700 16727 19703
rect 16850 19700 16856 19712
rect 16715 19672 16856 19700
rect 16715 19669 16727 19672
rect 16669 19663 16727 19669
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 17037 19703 17095 19709
rect 17037 19669 17049 19703
rect 17083 19700 17095 19703
rect 17218 19700 17224 19712
rect 17083 19672 17224 19700
rect 17083 19669 17095 19672
rect 17037 19663 17095 19669
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 17328 19700 17356 19740
rect 17948 19731 17960 19740
rect 17954 19728 17960 19731
rect 18012 19728 18018 19780
rect 19512 19771 19570 19777
rect 19512 19737 19524 19771
rect 19558 19768 19570 19771
rect 19610 19768 19616 19780
rect 19558 19740 19616 19768
rect 19558 19737 19570 19740
rect 19512 19731 19570 19737
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 20254 19768 20260 19780
rect 20167 19740 20260 19768
rect 17402 19700 17408 19712
rect 17328 19672 17408 19700
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 17589 19703 17647 19709
rect 17589 19669 17601 19703
rect 17635 19700 17647 19703
rect 18598 19700 18604 19712
rect 17635 19672 18604 19700
rect 17635 19669 17647 19672
rect 17589 19663 17647 19669
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 19061 19703 19119 19709
rect 19061 19669 19073 19703
rect 19107 19700 19119 19703
rect 20180 19700 20208 19740
rect 20254 19728 20260 19740
rect 20312 19768 20318 19780
rect 21085 19771 21143 19777
rect 21085 19768 21097 19771
rect 20312 19740 21097 19768
rect 20312 19728 20318 19740
rect 21085 19737 21097 19740
rect 21131 19737 21143 19771
rect 21085 19731 21143 19737
rect 19107 19672 20208 19700
rect 19107 19669 19119 19672
rect 19061 19663 19119 19669
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 20625 19703 20683 19709
rect 20625 19700 20637 19703
rect 20404 19672 20637 19700
rect 20404 19660 20410 19672
rect 20625 19669 20637 19672
rect 20671 19669 20683 19703
rect 21450 19700 21456 19712
rect 21411 19672 21456 19700
rect 20625 19663 20683 19669
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 22278 19700 22284 19712
rect 22239 19672 22284 19700
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 22428 19672 22473 19700
rect 22428 19660 22434 19672
rect 22554 19660 22560 19712
rect 22612 19700 22618 19712
rect 22741 19703 22799 19709
rect 22741 19700 22753 19703
rect 22612 19672 22753 19700
rect 22612 19660 22618 19672
rect 22741 19669 22753 19672
rect 22787 19669 22799 19703
rect 23014 19700 23020 19712
rect 22975 19672 23020 19700
rect 22741 19663 22799 19669
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 1104 19610 23460 19632
rect 1104 19558 6548 19610
rect 6600 19558 6612 19610
rect 6664 19558 6676 19610
rect 6728 19558 6740 19610
rect 6792 19558 6804 19610
rect 6856 19558 12146 19610
rect 12198 19558 12210 19610
rect 12262 19558 12274 19610
rect 12326 19558 12338 19610
rect 12390 19558 12402 19610
rect 12454 19558 17744 19610
rect 17796 19558 17808 19610
rect 17860 19558 17872 19610
rect 17924 19558 17936 19610
rect 17988 19558 18000 19610
rect 18052 19558 23460 19610
rect 1104 19536 23460 19558
rect 3050 19496 3056 19508
rect 3011 19468 3056 19496
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 3513 19499 3571 19505
rect 3513 19496 3525 19499
rect 3292 19468 3525 19496
rect 3292 19456 3298 19468
rect 3513 19465 3525 19468
rect 3559 19465 3571 19499
rect 4338 19496 4344 19508
rect 4299 19468 4344 19496
rect 3513 19459 3571 19465
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 4614 19496 4620 19508
rect 4575 19468 4620 19496
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 5350 19456 5356 19508
rect 5408 19496 5414 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 5408 19468 7849 19496
rect 5408 19456 5414 19468
rect 7837 19465 7849 19468
rect 7883 19465 7895 19499
rect 7837 19459 7895 19465
rect 9493 19499 9551 19505
rect 9493 19465 9505 19499
rect 9539 19496 9551 19499
rect 9674 19496 9680 19508
rect 9539 19468 9680 19496
rect 9539 19465 9551 19468
rect 9493 19459 9551 19465
rect 9674 19456 9680 19468
rect 9732 19496 9738 19508
rect 9858 19496 9864 19508
rect 9732 19468 9864 19496
rect 9732 19456 9738 19468
rect 9858 19456 9864 19468
rect 9916 19456 9922 19508
rect 10962 19496 10968 19508
rect 10923 19468 10968 19496
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11146 19496 11152 19508
rect 11107 19468 11152 19496
rect 11146 19456 11152 19468
rect 11204 19456 11210 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 12066 19496 12072 19508
rect 11563 19468 12072 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 12066 19456 12072 19468
rect 12124 19456 12130 19508
rect 13262 19496 13268 19508
rect 13223 19468 13268 19496
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 13541 19499 13599 19505
rect 13541 19465 13553 19499
rect 13587 19496 13599 19499
rect 13630 19496 13636 19508
rect 13587 19468 13636 19496
rect 13587 19465 13599 19468
rect 13541 19459 13599 19465
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 14369 19499 14427 19505
rect 14369 19465 14381 19499
rect 14415 19496 14427 19499
rect 15378 19496 15384 19508
rect 14415 19468 15384 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 15378 19456 15384 19468
rect 15436 19456 15442 19508
rect 15841 19499 15899 19505
rect 15841 19465 15853 19499
rect 15887 19465 15899 19499
rect 15841 19459 15899 19465
rect 16117 19499 16175 19505
rect 16117 19465 16129 19499
rect 16163 19496 16175 19499
rect 16390 19496 16396 19508
rect 16163 19468 16396 19496
rect 16163 19465 16175 19468
rect 16117 19459 16175 19465
rect 5810 19388 5816 19440
rect 5868 19428 5874 19440
rect 10410 19428 10416 19440
rect 5868 19400 8156 19428
rect 5868 19388 5874 19400
rect 3142 19360 3148 19372
rect 3103 19332 3148 19360
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 3602 19320 3608 19372
rect 3660 19360 3666 19372
rect 3881 19363 3939 19369
rect 3881 19360 3893 19363
rect 3660 19332 3893 19360
rect 3660 19320 3666 19332
rect 3881 19329 3893 19332
rect 3927 19329 3939 19363
rect 3881 19323 3939 19329
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19360 4031 19363
rect 4062 19360 4068 19372
rect 4019 19332 4068 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 4430 19360 4436 19372
rect 4391 19332 4436 19360
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 4522 19320 4528 19372
rect 4580 19360 4586 19372
rect 5166 19360 5172 19372
rect 4580 19332 5172 19360
rect 4580 19320 4586 19332
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 5925 19363 5983 19369
rect 5925 19329 5937 19363
rect 5971 19360 5983 19363
rect 6086 19360 6092 19372
rect 5971 19332 6092 19360
rect 5971 19329 5983 19332
rect 5925 19323 5983 19329
rect 6086 19320 6092 19332
rect 6144 19320 6150 19372
rect 6196 19369 6224 19400
rect 8128 19369 8156 19400
rect 8220 19400 10416 19428
rect 6181 19363 6239 19369
rect 6181 19329 6193 19363
rect 6227 19360 6239 19363
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 6227 19332 6377 19360
rect 6227 19329 6239 19332
rect 6181 19323 6239 19329
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6621 19363 6679 19369
rect 6621 19360 6633 19363
rect 6365 19323 6423 19329
rect 6472 19332 6633 19360
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 3418 19292 3424 19304
rect 3007 19264 3424 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3418 19252 3424 19264
rect 3476 19252 3482 19304
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 4338 19292 4344 19304
rect 3835 19264 4344 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 4338 19252 4344 19264
rect 4396 19292 4402 19304
rect 4798 19292 4804 19304
rect 4396 19264 4804 19292
rect 4396 19252 4402 19264
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 6472 19292 6500 19332
rect 6621 19329 6633 19332
rect 6667 19329 6679 19363
rect 6621 19323 6679 19329
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 6380 19264 6500 19292
rect 8036 19292 8064 19323
rect 8220 19292 8248 19400
rect 10410 19388 10416 19400
rect 10468 19388 10474 19440
rect 10870 19388 10876 19440
rect 10928 19428 10934 19440
rect 15562 19428 15568 19440
rect 10928 19400 15568 19428
rect 10928 19388 10934 19400
rect 8386 19369 8392 19372
rect 8380 19360 8392 19369
rect 8347 19332 8392 19360
rect 8380 19323 8392 19332
rect 8386 19320 8392 19323
rect 8444 19320 8450 19372
rect 9582 19360 9588 19372
rect 9543 19332 9588 19360
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 9841 19363 9899 19369
rect 9841 19360 9853 19363
rect 9692 19332 9853 19360
rect 9692 19292 9720 19332
rect 9841 19329 9853 19332
rect 9887 19329 9899 19363
rect 11330 19360 11336 19372
rect 11291 19332 11336 19360
rect 9841 19323 9899 19329
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 12641 19363 12699 19369
rect 12641 19329 12653 19363
rect 12687 19360 12699 19363
rect 12802 19360 12808 19372
rect 12687 19332 12808 19360
rect 12687 19329 12699 19332
rect 12641 19323 12699 19329
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 12912 19369 12940 19400
rect 12897 19363 12955 19369
rect 12897 19329 12909 19363
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19360 13139 19363
rect 13170 19360 13176 19372
rect 13127 19332 13176 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13170 19320 13176 19332
rect 13228 19360 13234 19372
rect 13357 19363 13415 19369
rect 13228 19332 13308 19360
rect 13228 19320 13234 19332
rect 8036 19264 8248 19292
rect 9600 19264 9720 19292
rect 13280 19292 13308 19332
rect 13357 19329 13369 19363
rect 13403 19360 13415 19363
rect 13630 19360 13636 19372
rect 13403 19332 13636 19360
rect 13403 19329 13415 19332
rect 13357 19323 13415 19329
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 13906 19360 13912 19372
rect 13867 19332 13912 19360
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 14366 19360 14372 19372
rect 14047 19332 14372 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 14476 19369 14504 19400
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 15856 19428 15884 19459
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 16666 19496 16672 19508
rect 16627 19468 16672 19496
rect 16666 19456 16672 19468
rect 16724 19456 16730 19508
rect 18141 19499 18199 19505
rect 18141 19465 18153 19499
rect 18187 19496 18199 19499
rect 18322 19496 18328 19508
rect 18187 19468 18328 19496
rect 18187 19465 18199 19468
rect 18141 19459 18199 19465
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 19610 19496 19616 19508
rect 19571 19468 19616 19496
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 21082 19496 21088 19508
rect 21043 19468 21088 19496
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 21358 19456 21364 19508
rect 21416 19456 21422 19508
rect 21450 19456 21456 19508
rect 21508 19496 21514 19508
rect 22281 19499 22339 19505
rect 22281 19496 22293 19499
rect 21508 19468 22293 19496
rect 21508 19456 21514 19468
rect 22281 19465 22293 19468
rect 22327 19465 22339 19499
rect 22281 19459 22339 19465
rect 16022 19428 16028 19440
rect 15856 19400 16028 19428
rect 16022 19388 16028 19400
rect 16080 19428 16086 19440
rect 16758 19428 16764 19440
rect 16080 19400 16764 19428
rect 16080 19388 16086 19400
rect 16758 19388 16764 19400
rect 16816 19388 16822 19440
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 17782 19431 17840 19437
rect 17782 19428 17794 19431
rect 17644 19400 17794 19428
rect 17644 19388 17650 19400
rect 17782 19397 17794 19400
rect 17828 19397 17840 19431
rect 17782 19391 17840 19397
rect 18064 19400 19564 19428
rect 14734 19369 14740 19372
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 14728 19323 14740 19369
rect 14792 19360 14798 19372
rect 15930 19360 15936 19372
rect 14792 19332 14828 19360
rect 15891 19332 15936 19360
rect 13722 19292 13728 19304
rect 13280 19264 13728 19292
rect 3234 19184 3240 19236
rect 3292 19224 3298 19236
rect 3292 19196 3648 19224
rect 3292 19184 3298 19196
rect 2685 19159 2743 19165
rect 2685 19125 2697 19159
rect 2731 19156 2743 19159
rect 3510 19156 3516 19168
rect 2731 19128 3516 19156
rect 2731 19125 2743 19128
rect 2685 19119 2743 19125
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 3620 19156 3648 19196
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 3620 19128 4813 19156
rect 4801 19125 4813 19128
rect 4847 19156 4859 19159
rect 6380 19156 6408 19264
rect 7742 19156 7748 19168
rect 4847 19128 6408 19156
rect 7703 19128 7748 19156
rect 4847 19125 4859 19128
rect 4801 19119 4859 19125
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 8478 19116 8484 19168
rect 8536 19156 8542 19168
rect 9600 19156 9628 19264
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 13817 19295 13875 19301
rect 13817 19261 13829 19295
rect 13863 19261 13875 19295
rect 13817 19255 13875 19261
rect 8536 19128 9628 19156
rect 13832 19156 13860 19255
rect 14182 19252 14188 19304
rect 14240 19292 14246 19304
rect 14476 19292 14504 19323
rect 14734 19320 14740 19323
rect 14792 19320 14798 19332
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16390 19360 16396 19372
rect 16172 19332 16252 19360
rect 16351 19332 16396 19360
rect 16172 19320 16178 19332
rect 14240 19264 14504 19292
rect 14240 19252 14246 19264
rect 16224 19233 16252 19332
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 18064 19369 18092 19400
rect 18049 19363 18107 19369
rect 16540 19332 16804 19360
rect 16540 19320 16546 19332
rect 16776 19304 16804 19332
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 19265 19363 19323 19369
rect 19265 19329 19277 19363
rect 19311 19360 19323 19363
rect 19426 19360 19432 19372
rect 19311 19332 19432 19360
rect 19311 19329 19323 19332
rect 19265 19323 19323 19329
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 19536 19369 19564 19400
rect 20438 19388 20444 19440
rect 20496 19428 20502 19440
rect 21376 19428 21404 19456
rect 22189 19431 22247 19437
rect 22189 19428 22201 19431
rect 20496 19400 21036 19428
rect 21376 19400 22201 19428
rect 20496 19388 20502 19400
rect 19521 19363 19579 19369
rect 19521 19329 19533 19363
rect 19567 19360 19579 19363
rect 20456 19360 20484 19388
rect 19567 19332 20484 19360
rect 20737 19363 20795 19369
rect 19567 19329 19579 19332
rect 19521 19323 19579 19329
rect 20737 19329 20749 19363
rect 20783 19360 20795 19363
rect 20898 19360 20904 19372
rect 20783 19332 20904 19360
rect 20783 19329 20795 19332
rect 20737 19323 20795 19329
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 21008 19369 21036 19400
rect 22189 19397 22201 19400
rect 22235 19397 22247 19431
rect 24118 19428 24124 19440
rect 22189 19391 22247 19397
rect 22664 19400 24124 19428
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19329 21051 19363
rect 21266 19360 21272 19372
rect 21227 19332 21272 19360
rect 20993 19323 21051 19329
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 21361 19363 21419 19369
rect 21361 19329 21373 19363
rect 21407 19360 21419 19363
rect 22664 19360 22692 19400
rect 24118 19388 24124 19400
rect 24176 19388 24182 19440
rect 22830 19360 22836 19372
rect 21407 19332 21496 19360
rect 21407 19329 21419 19332
rect 21361 19323 21419 19329
rect 16758 19252 16764 19304
rect 16816 19252 16822 19304
rect 16209 19227 16267 19233
rect 16209 19193 16221 19227
rect 16255 19193 16267 19227
rect 16209 19187 16267 19193
rect 19527 19196 20116 19224
rect 15194 19156 15200 19168
rect 13832 19128 15200 19156
rect 8536 19116 8542 19128
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 15654 19156 15660 19168
rect 15436 19128 15660 19156
rect 15436 19116 15442 19128
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 18506 19116 18512 19168
rect 18564 19156 18570 19168
rect 19527 19156 19555 19196
rect 18564 19128 19555 19156
rect 20088 19156 20116 19196
rect 21266 19156 21272 19168
rect 20088 19128 21272 19156
rect 18564 19116 18570 19128
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21468 19156 21496 19332
rect 21560 19332 22692 19360
rect 22791 19332 22836 19360
rect 21560 19233 21588 19332
rect 22830 19320 22836 19332
rect 22888 19320 22894 19372
rect 21726 19252 21732 19304
rect 21784 19252 21790 19304
rect 22462 19292 22468 19304
rect 22423 19264 22468 19292
rect 22462 19252 22468 19264
rect 22520 19252 22526 19304
rect 22741 19295 22799 19301
rect 22741 19261 22753 19295
rect 22787 19292 22799 19295
rect 23106 19292 23112 19304
rect 22787 19264 23112 19292
rect 22787 19261 22799 19264
rect 22741 19255 22799 19261
rect 23106 19252 23112 19264
rect 23164 19252 23170 19304
rect 21545 19227 21603 19233
rect 21545 19193 21557 19227
rect 21591 19193 21603 19227
rect 21545 19187 21603 19193
rect 21744 19168 21772 19252
rect 21827 19233 21833 19236
rect 21821 19187 21833 19233
rect 21885 19224 21891 19236
rect 21885 19196 21921 19224
rect 21827 19184 21833 19187
rect 21885 19184 21891 19196
rect 21634 19156 21640 19168
rect 21468 19128 21640 19156
rect 21634 19116 21640 19128
rect 21692 19116 21698 19168
rect 21726 19116 21732 19168
rect 21784 19116 21790 19168
rect 23017 19159 23075 19165
rect 23017 19125 23029 19159
rect 23063 19156 23075 19159
rect 23106 19156 23112 19168
rect 23063 19128 23112 19156
rect 23063 19125 23075 19128
rect 23017 19119 23075 19125
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 1104 19066 23460 19088
rect 1104 19014 3749 19066
rect 3801 19014 3813 19066
rect 3865 19014 3877 19066
rect 3929 19014 3941 19066
rect 3993 19014 4005 19066
rect 4057 19014 9347 19066
rect 9399 19014 9411 19066
rect 9463 19014 9475 19066
rect 9527 19014 9539 19066
rect 9591 19014 9603 19066
rect 9655 19014 14945 19066
rect 14997 19014 15009 19066
rect 15061 19014 15073 19066
rect 15125 19014 15137 19066
rect 15189 19014 15201 19066
rect 15253 19014 20543 19066
rect 20595 19014 20607 19066
rect 20659 19014 20671 19066
rect 20723 19014 20735 19066
rect 20787 19014 20799 19066
rect 20851 19014 23460 19066
rect 1104 18992 23460 19014
rect 3510 18912 3516 18964
rect 3568 18952 3574 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3568 18924 3801 18952
rect 3568 18912 3574 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 3789 18915 3847 18921
rect 4154 18912 4160 18964
rect 4212 18952 4218 18964
rect 4798 18952 4804 18964
rect 4212 18924 4804 18952
rect 4212 18912 4218 18924
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 6362 18952 6368 18964
rect 4908 18924 6368 18952
rect 3602 18884 3608 18896
rect 3563 18856 3608 18884
rect 3602 18844 3608 18856
rect 3660 18844 3666 18896
rect 4908 18884 4936 18924
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 8754 18952 8760 18964
rect 8715 18924 8760 18952
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 11790 18912 11796 18964
rect 11848 18952 11854 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 11848 18924 12449 18952
rect 11848 18912 11854 18924
rect 12437 18921 12449 18924
rect 12483 18921 12495 18955
rect 12437 18915 12495 18921
rect 12529 18955 12587 18961
rect 12529 18921 12541 18955
rect 12575 18952 12587 18955
rect 12802 18952 12808 18964
rect 12575 18924 12808 18952
rect 12575 18921 12587 18924
rect 12529 18915 12587 18921
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14148 18924 15056 18952
rect 14148 18912 14154 18924
rect 4816 18856 4936 18884
rect 15028 18884 15056 18924
rect 15286 18912 15292 18964
rect 15344 18952 15350 18964
rect 15473 18955 15531 18961
rect 15473 18952 15485 18955
rect 15344 18924 15485 18952
rect 15344 18912 15350 18924
rect 15473 18921 15485 18924
rect 15519 18921 15531 18955
rect 17034 18952 17040 18964
rect 15473 18915 15531 18921
rect 15580 18924 16620 18952
rect 16995 18924 17040 18952
rect 15580 18884 15608 18924
rect 15028 18856 15608 18884
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18816 3111 18819
rect 3418 18816 3424 18828
rect 3099 18788 3424 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 3973 18751 4031 18757
rect 3973 18748 3985 18751
rect 2823 18720 3985 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 3973 18717 3985 18720
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 4341 18751 4399 18757
rect 4341 18717 4353 18751
rect 4387 18748 4399 18751
rect 4816 18748 4844 18856
rect 5810 18816 5816 18828
rect 5771 18788 5816 18816
rect 5810 18776 5816 18788
rect 5868 18776 5874 18828
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8628 18788 8953 18816
rect 8628 18776 8634 18788
rect 8941 18785 8953 18788
rect 8987 18785 8999 18819
rect 8941 18779 8999 18785
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 11020 18788 11192 18816
rect 11020 18776 11026 18788
rect 4387 18720 4844 18748
rect 4387 18717 4399 18720
rect 4341 18711 4399 18717
rect 5166 18708 5172 18760
rect 5224 18748 5230 18760
rect 5546 18751 5604 18757
rect 5546 18748 5558 18751
rect 5224 18720 5558 18748
rect 5224 18708 5230 18720
rect 5546 18717 5558 18720
rect 5592 18748 5604 18751
rect 5718 18748 5724 18760
rect 5592 18720 5724 18748
rect 5592 18717 5604 18720
rect 5546 18711 5604 18717
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 5828 18748 5856 18776
rect 7285 18751 7343 18757
rect 7285 18748 7297 18751
rect 5828 18720 7297 18748
rect 7285 18717 7297 18720
rect 7331 18748 7343 18751
rect 7374 18748 7380 18760
rect 7331 18720 7380 18748
rect 7331 18717 7343 18720
rect 7285 18711 7343 18717
rect 7374 18708 7380 18720
rect 7432 18748 7438 18760
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 7432 18720 9229 18748
rect 7432 18708 7438 18720
rect 9217 18717 9229 18720
rect 9263 18748 9275 18751
rect 9401 18751 9459 18757
rect 9401 18748 9413 18751
rect 9263 18720 9413 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 9401 18717 9413 18720
rect 9447 18748 9459 18751
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9447 18720 9597 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9585 18717 9597 18720
rect 9631 18748 9643 18751
rect 9674 18748 9680 18760
rect 9631 18720 9680 18748
rect 9631 18717 9643 18720
rect 9585 18711 9643 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 9858 18757 9864 18760
rect 9852 18748 9864 18757
rect 9819 18720 9864 18748
rect 9852 18711 9864 18720
rect 9858 18708 9864 18711
rect 9916 18708 9922 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18717 11115 18751
rect 11164 18748 11192 18788
rect 11313 18751 11371 18757
rect 11313 18748 11325 18751
rect 11164 18720 11325 18748
rect 11057 18711 11115 18717
rect 11313 18717 11325 18720
rect 11359 18717 11371 18751
rect 11313 18711 11371 18717
rect 13909 18751 13967 18757
rect 13909 18717 13921 18751
rect 13955 18748 13967 18751
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 13955 18720 14105 18748
rect 13955 18717 13967 18720
rect 13909 18711 13967 18717
rect 14093 18717 14105 18720
rect 14139 18748 14151 18751
rect 14182 18748 14188 18760
rect 14139 18720 14188 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 3234 18680 3240 18692
rect 3195 18652 3240 18680
rect 3234 18640 3240 18652
rect 3292 18640 3298 18692
rect 4157 18683 4215 18689
rect 4157 18649 4169 18683
rect 4203 18649 4215 18683
rect 7006 18680 7012 18692
rect 7064 18689 7070 18692
rect 4157 18643 4215 18649
rect 4356 18652 5488 18680
rect 6976 18652 7012 18680
rect 2593 18615 2651 18621
rect 2593 18581 2605 18615
rect 2639 18612 2651 18615
rect 2958 18612 2964 18624
rect 2639 18584 2964 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 3145 18615 3203 18621
rect 3145 18581 3157 18615
rect 3191 18612 3203 18615
rect 3510 18612 3516 18624
rect 3191 18584 3516 18612
rect 3191 18581 3203 18584
rect 3145 18575 3203 18581
rect 3510 18572 3516 18584
rect 3568 18572 3574 18624
rect 4172 18612 4200 18643
rect 4356 18612 4384 18652
rect 4172 18584 4384 18612
rect 4433 18615 4491 18621
rect 4433 18581 4445 18615
rect 4479 18612 4491 18615
rect 5350 18612 5356 18624
rect 4479 18584 5356 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 5460 18612 5488 18652
rect 7006 18640 7012 18652
rect 7064 18643 7076 18689
rect 7644 18683 7702 18689
rect 7644 18649 7656 18683
rect 7690 18680 7702 18683
rect 8294 18680 8300 18692
rect 7690 18652 8300 18680
rect 7690 18649 7702 18652
rect 7644 18643 7702 18649
rect 7064 18640 7070 18643
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 9692 18680 9720 18708
rect 10870 18680 10876 18692
rect 9692 18652 10876 18680
rect 10870 18640 10876 18652
rect 10928 18680 10934 18692
rect 11072 18680 11100 18711
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 15378 18748 15384 18760
rect 14292 18720 15384 18748
rect 10928 18652 11100 18680
rect 10928 18640 10934 18652
rect 11422 18640 11428 18692
rect 11480 18680 11486 18692
rect 13664 18683 13722 18689
rect 13664 18680 13676 18683
rect 11480 18652 13676 18680
rect 11480 18640 11486 18652
rect 13664 18649 13676 18652
rect 13710 18680 13722 18683
rect 14292 18680 14320 18720
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 15562 18748 15568 18760
rect 15475 18720 15568 18748
rect 15562 18708 15568 18720
rect 15620 18748 15626 18760
rect 16390 18748 16396 18760
rect 15620 18720 16396 18748
rect 15620 18708 15626 18720
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 13710 18652 14320 18680
rect 14360 18683 14418 18689
rect 13710 18649 13722 18652
rect 13664 18643 13722 18649
rect 14360 18649 14372 18683
rect 14406 18680 14418 18683
rect 14918 18680 14924 18692
rect 14406 18652 14924 18680
rect 14406 18649 14418 18652
rect 14360 18643 14418 18649
rect 14918 18640 14924 18652
rect 14976 18640 14982 18692
rect 15832 18683 15890 18689
rect 15396 18652 15792 18680
rect 5905 18615 5963 18621
rect 5905 18612 5917 18615
rect 5460 18584 5917 18612
rect 5905 18581 5917 18584
rect 5951 18612 5963 18615
rect 5994 18612 6000 18624
rect 5951 18584 6000 18612
rect 5951 18581 5963 18584
rect 5905 18575 5963 18581
rect 5994 18572 6000 18584
rect 6052 18572 6058 18624
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7742 18612 7748 18624
rect 7156 18584 7748 18612
rect 7156 18572 7162 18584
rect 7742 18572 7748 18584
rect 7800 18572 7806 18624
rect 10965 18615 11023 18621
rect 10965 18581 10977 18615
rect 11011 18612 11023 18615
rect 12986 18612 12992 18624
rect 11011 18584 12992 18612
rect 11011 18581 11023 18584
rect 10965 18575 11023 18581
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 15396 18612 15424 18652
rect 13136 18584 15424 18612
rect 15764 18612 15792 18652
rect 15832 18649 15844 18683
rect 15878 18680 15890 18683
rect 16022 18680 16028 18692
rect 15878 18652 16028 18680
rect 15878 18649 15890 18652
rect 15832 18643 15890 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 16114 18612 16120 18624
rect 15764 18584 16120 18612
rect 13136 18572 13142 18584
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16592 18612 16620 18924
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 18046 18952 18052 18964
rect 17512 18924 18052 18952
rect 16945 18887 17003 18893
rect 16945 18853 16957 18887
rect 16991 18884 17003 18887
rect 17512 18884 17540 18924
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 18196 18924 18521 18952
rect 18196 18912 18202 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 18785 18955 18843 18961
rect 18785 18952 18797 18955
rect 18748 18924 18797 18952
rect 18748 18912 18754 18924
rect 18785 18921 18797 18924
rect 18831 18921 18843 18955
rect 18785 18915 18843 18921
rect 19610 18912 19616 18964
rect 19668 18952 19674 18964
rect 19668 18924 22692 18952
rect 19668 18912 19674 18924
rect 16991 18856 17540 18884
rect 20717 18887 20775 18893
rect 16991 18853 17003 18856
rect 16945 18847 17003 18853
rect 20717 18853 20729 18887
rect 20763 18884 20775 18887
rect 20990 18884 20996 18896
rect 20763 18856 20996 18884
rect 20763 18853 20775 18856
rect 20717 18847 20775 18853
rect 20990 18844 20996 18856
rect 21048 18844 21054 18896
rect 22664 18825 22692 18924
rect 18417 18819 18475 18825
rect 18417 18785 18429 18819
rect 18463 18816 18475 18819
rect 22649 18819 22707 18825
rect 18463 18788 19104 18816
rect 18463 18785 18475 18788
rect 18417 18779 18475 18785
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17000 18720 17540 18748
rect 17000 18708 17006 18720
rect 17512 18692 17540 18720
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18693 18751 18751 18757
rect 18693 18748 18705 18751
rect 18380 18720 18705 18748
rect 18380 18708 18386 18720
rect 18693 18717 18705 18720
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 18969 18751 19027 18757
rect 18969 18748 18981 18751
rect 18932 18720 18981 18748
rect 18932 18708 18938 18720
rect 18969 18717 18981 18720
rect 19015 18717 19027 18751
rect 19076 18748 19104 18788
rect 22649 18785 22661 18819
rect 22695 18785 22707 18819
rect 22649 18779 22707 18785
rect 22738 18776 22744 18828
rect 22796 18816 22802 18828
rect 22796 18788 22841 18816
rect 22796 18776 22802 18788
rect 19334 18748 19340 18760
rect 19076 18720 19340 18748
rect 18969 18711 19027 18717
rect 19334 18708 19340 18720
rect 19392 18748 19398 18760
rect 20530 18748 20536 18760
rect 19392 18720 20536 18748
rect 19392 18708 19398 18720
rect 20530 18708 20536 18720
rect 20588 18748 20594 18760
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 20588 18720 20637 18748
rect 20588 18708 20594 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 21830 18751 21888 18757
rect 21830 18748 21842 18751
rect 20772 18720 21842 18748
rect 20772 18708 20778 18720
rect 21830 18717 21842 18720
rect 21876 18717 21888 18751
rect 21830 18711 21888 18717
rect 22097 18751 22155 18757
rect 22097 18717 22109 18751
rect 22143 18748 22155 18751
rect 23014 18748 23020 18760
rect 22143 18720 23020 18748
rect 22143 18717 22155 18720
rect 22097 18711 22155 18717
rect 23014 18708 23020 18720
rect 23072 18708 23078 18760
rect 17494 18640 17500 18692
rect 17552 18680 17558 18692
rect 18150 18683 18208 18689
rect 18150 18680 18162 18683
rect 17552 18652 18162 18680
rect 17552 18640 17558 18652
rect 18150 18649 18162 18652
rect 18196 18649 18208 18683
rect 18150 18643 18208 18649
rect 18598 18640 18604 18692
rect 18656 18680 18662 18692
rect 18656 18652 20300 18680
rect 18656 18640 18662 18652
rect 17586 18612 17592 18624
rect 16592 18584 17592 18612
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 19245 18615 19303 18621
rect 19245 18581 19257 18615
rect 19291 18612 19303 18615
rect 19610 18612 19616 18624
rect 19291 18584 19616 18612
rect 19291 18581 19303 18584
rect 19245 18575 19303 18581
rect 19610 18572 19616 18584
rect 19668 18572 19674 18624
rect 20272 18612 20300 18652
rect 20346 18640 20352 18692
rect 20404 18689 20410 18692
rect 20404 18683 20438 18689
rect 20426 18680 20438 18683
rect 22557 18683 22615 18689
rect 22557 18680 22569 18683
rect 20426 18652 22569 18680
rect 20426 18649 20438 18652
rect 20404 18643 20438 18649
rect 22557 18649 22569 18652
rect 22603 18649 22615 18683
rect 22557 18643 22615 18649
rect 20404 18640 20410 18643
rect 21910 18612 21916 18624
rect 20272 18584 21916 18612
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 22189 18615 22247 18621
rect 22189 18581 22201 18615
rect 22235 18612 22247 18615
rect 22278 18612 22284 18624
rect 22235 18584 22284 18612
rect 22235 18581 22247 18584
rect 22189 18575 22247 18581
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 1104 18522 23460 18544
rect 1104 18470 6548 18522
rect 6600 18470 6612 18522
rect 6664 18470 6676 18522
rect 6728 18470 6740 18522
rect 6792 18470 6804 18522
rect 6856 18470 12146 18522
rect 12198 18470 12210 18522
rect 12262 18470 12274 18522
rect 12326 18470 12338 18522
rect 12390 18470 12402 18522
rect 12454 18470 17744 18522
rect 17796 18470 17808 18522
rect 17860 18470 17872 18522
rect 17924 18470 17936 18522
rect 17988 18470 18000 18522
rect 18052 18470 23460 18522
rect 1104 18448 23460 18470
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18408 2099 18411
rect 2866 18408 2872 18420
rect 2087 18380 2872 18408
rect 2087 18377 2099 18380
rect 2041 18371 2099 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3326 18368 3332 18420
rect 3384 18408 3390 18420
rect 3973 18411 4031 18417
rect 3973 18408 3985 18411
rect 3384 18380 3985 18408
rect 3384 18368 3390 18380
rect 3973 18377 3985 18380
rect 4019 18377 4031 18411
rect 4433 18411 4491 18417
rect 4433 18408 4445 18411
rect 3973 18371 4031 18377
rect 4080 18380 4445 18408
rect 2148 18312 2912 18340
rect 2148 18281 2176 18312
rect 2884 18281 2912 18312
rect 3510 18300 3516 18352
rect 3568 18340 3574 18352
rect 4080 18340 4108 18380
rect 4433 18377 4445 18380
rect 4479 18377 4491 18411
rect 4433 18371 4491 18377
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 4856 18380 4905 18408
rect 4856 18368 4862 18380
rect 4893 18377 4905 18380
rect 4939 18377 4951 18411
rect 4893 18371 4951 18377
rect 5261 18411 5319 18417
rect 5261 18377 5273 18411
rect 5307 18408 5319 18411
rect 5307 18380 7328 18408
rect 5307 18377 5319 18380
rect 5261 18371 5319 18377
rect 3568 18312 4108 18340
rect 5353 18343 5411 18349
rect 3568 18300 3574 18312
rect 5353 18309 5365 18343
rect 5399 18340 5411 18343
rect 7098 18340 7104 18352
rect 5399 18312 7104 18340
rect 5399 18309 5411 18312
rect 5353 18303 5411 18309
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 7300 18340 7328 18380
rect 7374 18368 7380 18420
rect 7432 18408 7438 18420
rect 7837 18411 7895 18417
rect 7837 18408 7849 18411
rect 7432 18380 7849 18408
rect 7432 18368 7438 18380
rect 7837 18377 7849 18380
rect 7883 18408 7895 18411
rect 8113 18411 8171 18417
rect 8113 18408 8125 18411
rect 7883 18380 8125 18408
rect 7883 18377 7895 18380
rect 7837 18371 7895 18377
rect 8113 18377 8125 18380
rect 8159 18408 8171 18411
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 8159 18380 8309 18408
rect 8159 18377 8171 18380
rect 8113 18371 8171 18377
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8478 18408 8484 18420
rect 8439 18380 8484 18408
rect 8297 18371 8355 18377
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 10226 18368 10232 18420
rect 10284 18368 10290 18420
rect 10870 18368 10876 18420
rect 10928 18408 10934 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 10928 18380 11529 18408
rect 10928 18368 10934 18380
rect 11517 18377 11529 18380
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 9030 18340 9036 18352
rect 7300 18312 9036 18340
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 9616 18343 9674 18349
rect 9616 18309 9628 18343
rect 9662 18340 9674 18343
rect 10244 18340 10272 18368
rect 9662 18312 10272 18340
rect 9662 18309 9674 18312
rect 9616 18303 9674 18309
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18241 2835 18275
rect 2777 18235 2835 18241
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 3234 18272 3240 18284
rect 2915 18244 3240 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 1872 18204 1900 18235
rect 2792 18204 2820 18235
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 3418 18232 3424 18284
rect 3476 18232 3482 18284
rect 3605 18275 3663 18281
rect 5815 18276 5873 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 5736 18275 5873 18276
rect 3651 18244 4108 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 1872 18176 2452 18204
rect 2792 18176 2912 18204
rect 2424 18145 2452 18176
rect 2409 18139 2467 18145
rect 2409 18105 2421 18139
rect 2455 18105 2467 18139
rect 2884 18136 2912 18176
rect 2958 18164 2964 18216
rect 3016 18204 3022 18216
rect 3329 18207 3387 18213
rect 3016 18176 3061 18204
rect 3016 18164 3022 18176
rect 3329 18173 3341 18207
rect 3375 18204 3387 18207
rect 3436 18204 3464 18232
rect 3375 18176 3464 18204
rect 3513 18207 3571 18213
rect 3375 18173 3387 18176
rect 3329 18167 3387 18173
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3878 18204 3884 18216
rect 3559 18176 3884 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 3418 18136 3424 18148
rect 2884 18108 3424 18136
rect 2409 18099 2467 18105
rect 3418 18096 3424 18108
rect 3476 18096 3482 18148
rect 4080 18136 4108 18244
rect 5736 18248 5827 18275
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 4212 18176 4261 18204
rect 4212 18164 4218 18176
rect 4249 18173 4261 18176
rect 4295 18173 4307 18207
rect 4249 18167 4307 18173
rect 4341 18207 4399 18213
rect 4341 18173 4353 18207
rect 4387 18204 4399 18207
rect 4614 18204 4620 18216
rect 4387 18176 4620 18204
rect 4387 18173 4399 18176
rect 4341 18167 4399 18173
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5445 18207 5503 18213
rect 5445 18204 5457 18207
rect 5316 18176 5457 18204
rect 5316 18164 5322 18176
rect 5445 18173 5457 18176
rect 5491 18204 5503 18207
rect 5736 18204 5764 18248
rect 5815 18241 5827 18248
rect 5861 18241 5873 18275
rect 5815 18235 5873 18241
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 6621 18275 6679 18281
rect 6621 18272 6633 18275
rect 6512 18244 6633 18272
rect 6512 18232 6518 18244
rect 6621 18241 6633 18244
rect 6667 18241 6679 18275
rect 6621 18235 6679 18241
rect 9766 18232 9772 18284
rect 9824 18272 9830 18284
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9824 18244 9873 18272
rect 9824 18232 9830 18244
rect 9861 18241 9873 18244
rect 9907 18272 9919 18275
rect 9953 18275 10011 18281
rect 9953 18272 9965 18275
rect 9907 18244 9965 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 9953 18241 9965 18244
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10220 18275 10278 18281
rect 10220 18241 10232 18275
rect 10266 18272 10278 18275
rect 10502 18272 10508 18284
rect 10266 18244 10508 18272
rect 10266 18241 10278 18244
rect 10220 18235 10278 18241
rect 10502 18232 10508 18244
rect 10560 18272 10566 18284
rect 11532 18272 11560 18371
rect 13998 18368 14004 18420
rect 14056 18408 14062 18420
rect 14645 18411 14703 18417
rect 14645 18408 14657 18411
rect 14056 18380 14657 18408
rect 14056 18368 14062 18380
rect 14645 18377 14657 18380
rect 14691 18377 14703 18411
rect 14645 18371 14703 18377
rect 14734 18368 14740 18420
rect 14792 18408 14798 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 14792 18380 16681 18408
rect 14792 18368 14798 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 16669 18371 16727 18377
rect 17310 18368 17316 18420
rect 17368 18408 17374 18420
rect 17405 18411 17463 18417
rect 17405 18408 17417 18411
rect 17368 18380 17417 18408
rect 17368 18368 17374 18380
rect 17405 18377 17417 18380
rect 17451 18377 17463 18411
rect 17405 18371 17463 18377
rect 17586 18368 17592 18420
rect 17644 18408 17650 18420
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 17644 18380 21833 18408
rect 17644 18368 17650 18380
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 22278 18408 22284 18420
rect 22239 18380 22284 18408
rect 21821 18371 21879 18377
rect 22278 18368 22284 18380
rect 22336 18368 22342 18420
rect 22738 18408 22744 18420
rect 22699 18380 22744 18408
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 11968 18343 12026 18349
rect 11968 18309 11980 18343
rect 12014 18340 12026 18343
rect 12066 18340 12072 18352
rect 12014 18312 12072 18340
rect 12014 18309 12026 18312
rect 11968 18303 12026 18309
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 12618 18300 12624 18352
rect 12676 18300 12682 18352
rect 15562 18340 15568 18352
rect 14568 18312 15568 18340
rect 11701 18275 11759 18281
rect 11701 18272 11713 18275
rect 10560 18244 11192 18272
rect 11532 18244 11713 18272
rect 10560 18232 10566 18244
rect 6178 18204 6184 18216
rect 5491 18176 5764 18204
rect 6012 18176 6184 18204
rect 5491 18173 5503 18176
rect 5445 18167 5503 18173
rect 5350 18136 5356 18148
rect 4080 18108 5356 18136
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 6012 18145 6040 18176
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 6365 18207 6423 18213
rect 6365 18173 6377 18207
rect 6411 18173 6423 18207
rect 11164 18204 11192 18244
rect 11701 18241 11713 18244
rect 11747 18241 11759 18275
rect 12636 18272 12664 18300
rect 11701 18235 11759 18241
rect 11788 18244 12664 18272
rect 11788 18204 11816 18244
rect 14274 18232 14280 18284
rect 14332 18281 14338 18284
rect 14568 18281 14596 18312
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 16206 18300 16212 18352
rect 16264 18340 16270 18352
rect 16264 18312 16988 18340
rect 16264 18300 16270 18312
rect 14332 18272 14344 18281
rect 14553 18275 14611 18281
rect 14332 18244 14377 18272
rect 14332 18235 14344 18244
rect 14553 18241 14565 18275
rect 14599 18241 14611 18275
rect 15758 18275 15816 18281
rect 15758 18272 15770 18275
rect 14553 18235 14611 18241
rect 14660 18244 15770 18272
rect 14332 18232 14338 18235
rect 11164 18176 11816 18204
rect 6365 18167 6423 18173
rect 5997 18139 6055 18145
rect 5997 18105 6009 18139
rect 6043 18105 6055 18139
rect 6380 18136 6408 18167
rect 5997 18099 6055 18105
rect 6196 18108 6408 18136
rect 7745 18139 7803 18145
rect 2317 18071 2375 18077
rect 2317 18037 2329 18071
rect 2363 18068 2375 18071
rect 3050 18068 3056 18080
rect 2363 18040 3056 18068
rect 2363 18037 2375 18040
rect 2317 18031 2375 18037
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 4982 18068 4988 18080
rect 4847 18040 4988 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 6086 18068 6092 18080
rect 6047 18040 6092 18068
rect 6086 18028 6092 18040
rect 6144 18068 6150 18080
rect 6196 18068 6224 18108
rect 7745 18105 7757 18139
rect 7791 18136 7803 18139
rect 8294 18136 8300 18148
rect 7791 18108 8300 18136
rect 7791 18105 7803 18108
rect 7745 18099 7803 18105
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 11333 18139 11391 18145
rect 11333 18105 11345 18139
rect 11379 18136 11391 18139
rect 11422 18136 11428 18148
rect 11379 18108 11428 18136
rect 11379 18105 11391 18108
rect 11333 18099 11391 18105
rect 11422 18096 11428 18108
rect 11480 18096 11486 18148
rect 13078 18136 13084 18148
rect 13039 18108 13084 18136
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 13170 18096 13176 18148
rect 13228 18136 13234 18148
rect 14660 18136 14688 18244
rect 15758 18241 15770 18244
rect 15804 18241 15816 18275
rect 15758 18235 15816 18241
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16172 18244 16217 18272
rect 16172 18232 16178 18244
rect 16025 18207 16083 18213
rect 16025 18173 16037 18207
rect 16071 18204 16083 18207
rect 16390 18204 16396 18216
rect 16071 18176 16396 18204
rect 16071 18173 16083 18176
rect 16025 18167 16083 18173
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 16960 18204 16988 18312
rect 17126 18300 17132 18352
rect 17184 18340 17190 18352
rect 17184 18312 17632 18340
rect 17184 18300 17190 18312
rect 17034 18232 17040 18284
rect 17092 18272 17098 18284
rect 17604 18281 17632 18312
rect 18046 18300 18052 18352
rect 18104 18340 18110 18352
rect 18598 18340 18604 18352
rect 18104 18312 18604 18340
rect 18104 18300 18110 18312
rect 18598 18300 18604 18312
rect 18656 18300 18662 18352
rect 19334 18340 19340 18352
rect 18800 18312 19340 18340
rect 18800 18281 18828 18312
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 20162 18300 20168 18352
rect 20220 18340 20226 18352
rect 20622 18340 20628 18352
rect 20220 18312 20628 18340
rect 20220 18300 20226 18312
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 21726 18300 21732 18352
rect 21784 18340 21790 18352
rect 22833 18343 22891 18349
rect 22833 18340 22845 18343
rect 21784 18312 22845 18340
rect 21784 18300 21790 18312
rect 22833 18309 22845 18312
rect 22879 18309 22891 18343
rect 22833 18303 22891 18309
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 17092 18244 17233 18272
rect 17092 18232 17098 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18241 17647 18275
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 17589 18235 17647 18241
rect 17696 18244 18429 18272
rect 17696 18204 17724 18244
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 19052 18275 19110 18281
rect 19052 18241 19064 18275
rect 19098 18272 19110 18275
rect 19426 18272 19432 18284
rect 19098 18244 19432 18272
rect 19098 18241 19110 18244
rect 19052 18235 19110 18241
rect 19426 18232 19432 18244
rect 19484 18272 19490 18284
rect 19886 18272 19892 18284
rect 19484 18244 19892 18272
rect 19484 18232 19490 18244
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 20513 18275 20571 18281
rect 20513 18272 20525 18275
rect 19996 18244 20525 18272
rect 18230 18204 18236 18216
rect 16960 18176 17724 18204
rect 18191 18176 18236 18204
rect 18230 18164 18236 18176
rect 18288 18164 18294 18216
rect 18322 18136 18328 18148
rect 13228 18108 13273 18136
rect 14568 18108 14688 18136
rect 16040 18108 18328 18136
rect 13228 18096 13234 18108
rect 6144 18040 6224 18068
rect 6144 18028 6150 18040
rect 8846 18028 8852 18080
rect 8904 18068 8910 18080
rect 11238 18068 11244 18080
rect 8904 18040 11244 18068
rect 8904 18028 8910 18040
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 11698 18028 11704 18080
rect 11756 18068 11762 18080
rect 14568 18068 14596 18108
rect 11756 18040 14596 18068
rect 11756 18028 11762 18040
rect 14642 18028 14648 18080
rect 14700 18068 14706 18080
rect 16040 18068 16068 18108
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 14700 18040 16068 18068
rect 14700 18028 14706 18040
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16301 18071 16359 18077
rect 16301 18068 16313 18071
rect 16172 18040 16313 18068
rect 16172 18028 16178 18040
rect 16301 18037 16313 18040
rect 16347 18037 16359 18071
rect 16301 18031 16359 18037
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 16448 18040 16493 18068
rect 16448 18028 16454 18040
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 17681 18071 17739 18077
rect 17681 18068 17693 18071
rect 17644 18040 17693 18068
rect 17644 18028 17650 18040
rect 17681 18037 17693 18040
rect 17727 18037 17739 18071
rect 17681 18031 17739 18037
rect 18138 18028 18144 18080
rect 18196 18068 18202 18080
rect 18782 18068 18788 18080
rect 18196 18040 18788 18068
rect 18196 18028 18202 18040
rect 18782 18028 18788 18040
rect 18840 18068 18846 18080
rect 19996 18068 20024 18244
rect 20513 18241 20525 18244
rect 20559 18241 20571 18275
rect 20513 18235 20571 18241
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 21048 18244 22201 18272
rect 21048 18232 21054 18244
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 20128 18176 20269 18204
rect 20128 18164 20134 18176
rect 20257 18173 20269 18176
rect 20303 18173 20315 18207
rect 22462 18204 22468 18216
rect 22423 18176 22468 18204
rect 20257 18167 20315 18173
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 20162 18136 20168 18148
rect 20123 18108 20168 18136
rect 20162 18096 20168 18108
rect 20220 18096 20226 18148
rect 21266 18096 21272 18148
rect 21324 18136 21330 18148
rect 23017 18139 23075 18145
rect 23017 18136 23029 18139
rect 21324 18108 23029 18136
rect 21324 18096 21330 18108
rect 23017 18105 23029 18108
rect 23063 18105 23075 18139
rect 23017 18099 23075 18105
rect 18840 18040 20024 18068
rect 18840 18028 18846 18040
rect 20254 18028 20260 18080
rect 20312 18068 20318 18080
rect 21542 18068 21548 18080
rect 20312 18040 21548 18068
rect 20312 18028 20318 18040
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 21637 18071 21695 18077
rect 21637 18037 21649 18071
rect 21683 18068 21695 18071
rect 21910 18068 21916 18080
rect 21683 18040 21916 18068
rect 21683 18037 21695 18040
rect 21637 18031 21695 18037
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 1104 17978 23460 18000
rect 1104 17926 3749 17978
rect 3801 17926 3813 17978
rect 3865 17926 3877 17978
rect 3929 17926 3941 17978
rect 3993 17926 4005 17978
rect 4057 17926 9347 17978
rect 9399 17926 9411 17978
rect 9463 17926 9475 17978
rect 9527 17926 9539 17978
rect 9591 17926 9603 17978
rect 9655 17926 14945 17978
rect 14997 17926 15009 17978
rect 15061 17926 15073 17978
rect 15125 17926 15137 17978
rect 15189 17926 15201 17978
rect 15253 17926 20543 17978
rect 20595 17926 20607 17978
rect 20659 17926 20671 17978
rect 20723 17926 20735 17978
rect 20787 17926 20799 17978
rect 20851 17926 23460 17978
rect 1104 17904 23460 17926
rect 3142 17824 3148 17876
rect 3200 17864 3206 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3200 17836 3801 17864
rect 3200 17824 3206 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 5902 17864 5908 17876
rect 3789 17827 3847 17833
rect 4448 17836 5908 17864
rect 4448 17796 4476 17836
rect 5902 17824 5908 17836
rect 5960 17824 5966 17876
rect 6270 17824 6276 17876
rect 6328 17864 6334 17876
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 6328 17836 9689 17864
rect 6328 17824 6334 17836
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 9677 17827 9735 17833
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 13170 17864 13176 17876
rect 11296 17836 13176 17864
rect 11296 17824 11302 17836
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 13909 17867 13967 17873
rect 13909 17833 13921 17867
rect 13955 17864 13967 17867
rect 14458 17864 14464 17876
rect 13955 17836 14464 17864
rect 13955 17833 13967 17836
rect 13909 17827 13967 17833
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 15473 17867 15531 17873
rect 15473 17833 15485 17867
rect 15519 17864 15531 17867
rect 16574 17864 16580 17876
rect 15519 17836 16580 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 17313 17867 17371 17873
rect 17313 17833 17325 17867
rect 17359 17864 17371 17867
rect 18966 17864 18972 17876
rect 17359 17836 18972 17864
rect 17359 17833 17371 17836
rect 17313 17827 17371 17833
rect 18966 17824 18972 17836
rect 19024 17824 19030 17876
rect 19061 17867 19119 17873
rect 19061 17833 19073 17867
rect 19107 17864 19119 17867
rect 19518 17864 19524 17876
rect 19107 17836 19524 17864
rect 19107 17833 19119 17836
rect 19061 17827 19119 17833
rect 19518 17824 19524 17836
rect 19576 17864 19582 17876
rect 19978 17864 19984 17876
rect 19576 17836 19984 17864
rect 19576 17824 19582 17836
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 20438 17824 20444 17876
rect 20496 17864 20502 17876
rect 20496 17836 20668 17864
rect 20496 17824 20502 17836
rect 19242 17796 19248 17808
rect 2792 17768 4476 17796
rect 19203 17768 19248 17796
rect 2792 17737 2820 17768
rect 19242 17756 19248 17768
rect 19300 17756 19306 17808
rect 20640 17796 20668 17836
rect 21358 17824 21364 17876
rect 21416 17864 21422 17876
rect 21726 17864 21732 17876
rect 21416 17836 21732 17864
rect 21416 17824 21422 17836
rect 21726 17824 21732 17836
rect 21784 17824 21790 17876
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 22741 17867 22799 17873
rect 22741 17864 22753 17867
rect 22520 17836 22753 17864
rect 22520 17824 22526 17836
rect 22741 17833 22753 17836
rect 22787 17864 22799 17867
rect 23198 17864 23204 17876
rect 22787 17836 23204 17864
rect 22787 17833 22799 17836
rect 22741 17827 22799 17833
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 20640 17768 23152 17796
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17697 2835 17731
rect 2777 17691 2835 17697
rect 2866 17688 2872 17740
rect 2924 17728 2930 17740
rect 2961 17731 3019 17737
rect 2961 17728 2973 17731
rect 2924 17700 2973 17728
rect 2924 17688 2930 17700
rect 2961 17697 2973 17700
rect 3007 17697 3019 17731
rect 2961 17691 3019 17697
rect 3418 17688 3424 17740
rect 3476 17728 3482 17740
rect 16945 17731 17003 17737
rect 3476 17700 4200 17728
rect 3476 17688 3482 17700
rect 3050 17660 3056 17672
rect 3011 17632 3056 17660
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 3602 17620 3608 17672
rect 3660 17660 3666 17672
rect 4172 17669 4200 17700
rect 16945 17697 16957 17731
rect 16991 17728 17003 17731
rect 20901 17731 20959 17737
rect 16991 17700 17724 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3660 17632 3985 17660
rect 3660 17620 3666 17632
rect 3973 17629 3985 17632
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 6086 17660 6092 17672
rect 4479 17632 6092 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4816 17604 4844 17632
rect 6086 17620 6092 17632
rect 6144 17660 6150 17672
rect 7285 17663 7343 17669
rect 7285 17660 7297 17663
rect 6144 17632 7297 17660
rect 6144 17620 6150 17632
rect 7285 17629 7297 17632
rect 7331 17660 7343 17663
rect 8757 17663 8815 17669
rect 8757 17660 8769 17663
rect 7331 17632 8769 17660
rect 7331 17629 7343 17632
rect 7285 17623 7343 17629
rect 8757 17629 8769 17632
rect 8803 17660 8815 17663
rect 9033 17663 9091 17669
rect 9033 17660 9045 17663
rect 8803 17632 9045 17660
rect 8803 17629 8815 17632
rect 8757 17623 8815 17629
rect 9033 17629 9045 17632
rect 9079 17660 9091 17663
rect 9122 17660 9128 17672
rect 9079 17632 9128 17660
rect 9079 17629 9091 17632
rect 9033 17623 9091 17629
rect 9122 17620 9128 17632
rect 9180 17660 9186 17672
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 9180 17632 9229 17660
rect 9180 17620 9186 17632
rect 9217 17629 9229 17632
rect 9263 17660 9275 17663
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 9263 17632 9413 17660
rect 9263 17629 9275 17632
rect 9217 17623 9275 17629
rect 9401 17629 9413 17632
rect 9447 17660 9459 17663
rect 9585 17663 9643 17669
rect 9585 17660 9597 17663
rect 9447 17632 9597 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 9585 17629 9597 17632
rect 9631 17660 9643 17663
rect 11054 17660 11060 17672
rect 9631 17632 11060 17660
rect 9631 17629 9643 17632
rect 9585 17623 9643 17629
rect 11054 17620 11060 17632
rect 11112 17660 11118 17672
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 11112 17632 11253 17660
rect 11112 17620 11118 17632
rect 11241 17629 11253 17632
rect 11287 17660 11299 17663
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 11287 17632 11529 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11517 17629 11529 17632
rect 11563 17660 11575 17663
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11563 17632 11805 17660
rect 11563 17629 11575 17632
rect 11517 17623 11575 17629
rect 11793 17629 11805 17632
rect 11839 17660 11851 17663
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 11839 17632 11989 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 11977 17629 11989 17632
rect 12023 17660 12035 17663
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 12023 17632 12173 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 12161 17629 12173 17632
rect 12207 17660 12219 17663
rect 12253 17663 12311 17669
rect 12253 17660 12265 17663
rect 12207 17632 12265 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12253 17629 12265 17632
rect 12299 17660 12311 17663
rect 12986 17660 12992 17672
rect 12299 17632 12992 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 14090 17660 14096 17672
rect 13780 17632 13825 17660
rect 14051 17632 14096 17660
rect 13780 17620 13786 17632
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 16390 17620 16396 17672
rect 16448 17660 16454 17672
rect 16960 17660 16988 17691
rect 17126 17660 17132 17672
rect 16448 17632 16988 17660
rect 17087 17632 17132 17660
rect 16448 17620 16454 17632
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 17696 17669 17724 17700
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21358 17728 21364 17740
rect 20947 17700 21364 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22094 17728 22100 17740
rect 22051 17700 22100 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 17681 17663 17739 17669
rect 17681 17629 17693 17663
rect 17727 17660 17739 17663
rect 19334 17660 19340 17672
rect 17727 17632 19340 17660
rect 17727 17629 17739 17632
rect 17681 17623 17739 17629
rect 18156 17604 18184 17632
rect 19334 17620 19340 17632
rect 19392 17620 19398 17672
rect 20625 17663 20683 17669
rect 19444 17632 20484 17660
rect 4706 17601 4712 17604
rect 4700 17592 4712 17601
rect 3436 17564 4476 17592
rect 4667 17564 4712 17592
rect 3436 17533 3464 17564
rect 3421 17527 3479 17533
rect 3421 17493 3433 17527
rect 3467 17493 3479 17527
rect 3421 17487 3479 17493
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 4341 17527 4399 17533
rect 4341 17524 4353 17527
rect 4120 17496 4353 17524
rect 4120 17484 4126 17496
rect 4341 17493 4353 17496
rect 4387 17493 4399 17527
rect 4448 17524 4476 17564
rect 4700 17555 4712 17564
rect 4706 17552 4712 17555
rect 4764 17552 4770 17604
rect 4798 17552 4804 17604
rect 4856 17552 4862 17604
rect 5718 17592 5724 17604
rect 4908 17564 5724 17592
rect 4908 17524 4936 17564
rect 5718 17552 5724 17564
rect 5776 17552 5782 17604
rect 5994 17552 6000 17604
rect 6052 17592 6058 17604
rect 7018 17595 7076 17601
rect 7018 17592 7030 17595
rect 6052 17564 7030 17592
rect 6052 17552 6058 17564
rect 7018 17561 7030 17564
rect 7064 17561 7076 17595
rect 7018 17555 7076 17561
rect 7190 17552 7196 17604
rect 7248 17592 7254 17604
rect 8490 17595 8548 17601
rect 8490 17592 8502 17595
rect 7248 17564 8502 17592
rect 7248 17552 7254 17564
rect 8490 17561 8502 17564
rect 8536 17561 8548 17595
rect 8490 17555 8548 17561
rect 10226 17552 10232 17604
rect 10284 17592 10290 17604
rect 12526 17601 12532 17604
rect 10790 17595 10848 17601
rect 10790 17592 10802 17595
rect 10284 17564 10802 17592
rect 10284 17552 10290 17564
rect 10790 17561 10802 17564
rect 10836 17561 10848 17595
rect 10790 17555 10848 17561
rect 12520 17555 12532 17601
rect 12584 17592 12590 17604
rect 14360 17595 14418 17601
rect 14360 17592 14372 17595
rect 12584 17564 12620 17592
rect 13648 17564 14372 17592
rect 12526 17552 12532 17555
rect 12584 17552 12590 17564
rect 4448 17496 4936 17524
rect 4341 17487 4399 17493
rect 5074 17484 5080 17536
rect 5132 17524 5138 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5132 17496 5825 17524
rect 5132 17484 5138 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 7374 17524 7380 17536
rect 7335 17496 7380 17524
rect 5813 17487 5871 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 7466 17484 7472 17536
rect 7524 17524 7530 17536
rect 10318 17524 10324 17536
rect 7524 17496 10324 17524
rect 7524 17484 7530 17496
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 13648 17533 13676 17564
rect 14360 17561 14372 17564
rect 14406 17592 14418 17595
rect 14406 17564 15700 17592
rect 14406 17561 14418 17564
rect 14360 17555 14418 17561
rect 13633 17527 13691 17533
rect 13633 17493 13645 17527
rect 13679 17493 13691 17527
rect 13633 17487 13691 17493
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 14550 17524 14556 17536
rect 14240 17496 14556 17524
rect 14240 17484 14246 17496
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 14826 17484 14832 17536
rect 14884 17524 14890 17536
rect 15565 17527 15623 17533
rect 15565 17524 15577 17527
rect 14884 17496 15577 17524
rect 14884 17484 14890 17496
rect 15565 17493 15577 17496
rect 15611 17493 15623 17527
rect 15672 17524 15700 17564
rect 16666 17552 16672 17604
rect 16724 17601 16730 17604
rect 16724 17592 16736 17601
rect 17948 17595 18006 17601
rect 16724 17564 16769 17592
rect 16868 17564 17724 17592
rect 16724 17555 16736 17564
rect 16724 17552 16730 17555
rect 16868 17524 16896 17564
rect 15672 17496 16896 17524
rect 15565 17487 15623 17493
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 17460 17496 17601 17524
rect 17460 17484 17466 17496
rect 17589 17493 17601 17496
rect 17635 17493 17647 17527
rect 17696 17524 17724 17564
rect 17948 17561 17960 17595
rect 17994 17592 18006 17595
rect 18046 17592 18052 17604
rect 17994 17564 18052 17592
rect 17994 17561 18006 17564
rect 17948 17555 18006 17561
rect 18046 17552 18052 17564
rect 18104 17552 18110 17604
rect 18138 17552 18144 17604
rect 18196 17552 18202 17604
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 19444 17592 19472 17632
rect 18656 17564 19472 17592
rect 18656 17552 18662 17564
rect 19610 17552 19616 17604
rect 19668 17592 19674 17604
rect 20162 17592 20168 17604
rect 19668 17564 20168 17592
rect 19668 17552 19674 17564
rect 20162 17552 20168 17564
rect 20220 17552 20226 17604
rect 20346 17592 20352 17604
rect 20404 17601 20410 17604
rect 20316 17564 20352 17592
rect 20346 17552 20352 17564
rect 20404 17555 20416 17601
rect 20456 17592 20484 17632
rect 20625 17629 20637 17663
rect 20671 17660 20683 17663
rect 20714 17660 20720 17672
rect 20671 17632 20720 17660
rect 20671 17629 20683 17632
rect 20625 17623 20683 17629
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 21542 17660 21548 17672
rect 21503 17632 21548 17660
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 22833 17663 22891 17669
rect 22833 17660 22845 17663
rect 21652 17632 22845 17660
rect 21652 17592 21680 17632
rect 22833 17629 22845 17632
rect 22879 17629 22891 17663
rect 22833 17623 22891 17629
rect 20456 17564 21680 17592
rect 22097 17595 22155 17601
rect 22097 17561 22109 17595
rect 22143 17592 22155 17595
rect 22278 17592 22284 17604
rect 22143 17564 22284 17592
rect 22143 17561 22155 17564
rect 22097 17555 22155 17561
rect 20404 17552 20410 17555
rect 22278 17552 22284 17564
rect 22336 17552 22342 17604
rect 23124 17536 23152 17768
rect 20993 17527 21051 17533
rect 20993 17524 21005 17527
rect 17696 17496 21005 17524
rect 17589 17487 17647 17493
rect 20993 17493 21005 17496
rect 21039 17493 21051 17527
rect 20993 17487 21051 17493
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 21140 17496 21185 17524
rect 21140 17484 21146 17496
rect 21266 17484 21272 17536
rect 21324 17524 21330 17536
rect 21453 17527 21511 17533
rect 21453 17524 21465 17527
rect 21324 17496 21465 17524
rect 21324 17484 21330 17496
rect 21453 17493 21465 17496
rect 21499 17493 21511 17527
rect 21453 17487 21511 17493
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 22244 17496 22289 17524
rect 22244 17484 22250 17496
rect 22462 17484 22468 17536
rect 22520 17524 22526 17536
rect 22557 17527 22615 17533
rect 22557 17524 22569 17527
rect 22520 17496 22569 17524
rect 22520 17484 22526 17496
rect 22557 17493 22569 17496
rect 22603 17493 22615 17527
rect 23106 17524 23112 17536
rect 23067 17496 23112 17524
rect 22557 17487 22615 17493
rect 23106 17484 23112 17496
rect 23164 17484 23170 17536
rect 1104 17434 23460 17456
rect 1104 17382 6548 17434
rect 6600 17382 6612 17434
rect 6664 17382 6676 17434
rect 6728 17382 6740 17434
rect 6792 17382 6804 17434
rect 6856 17382 12146 17434
rect 12198 17382 12210 17434
rect 12262 17382 12274 17434
rect 12326 17382 12338 17434
rect 12390 17382 12402 17434
rect 12454 17382 17744 17434
rect 17796 17382 17808 17434
rect 17860 17382 17872 17434
rect 17924 17382 17936 17434
rect 17988 17382 18000 17434
rect 18052 17382 23460 17434
rect 1104 17360 23460 17382
rect 3881 17323 3939 17329
rect 3881 17289 3893 17323
rect 3927 17320 3939 17323
rect 4614 17320 4620 17332
rect 3927 17292 4620 17320
rect 3927 17289 3939 17292
rect 3881 17283 3939 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 6270 17320 6276 17332
rect 4816 17292 6276 17320
rect 4157 17255 4215 17261
rect 4157 17221 4169 17255
rect 4203 17252 4215 17255
rect 4816 17252 4844 17292
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6733 17323 6791 17329
rect 6733 17289 6745 17323
rect 6779 17320 6791 17323
rect 8018 17320 8024 17332
rect 6779 17292 8024 17320
rect 6779 17289 6791 17292
rect 6733 17283 6791 17289
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 9030 17320 9036 17332
rect 8991 17292 9036 17320
rect 9030 17280 9036 17292
rect 9088 17280 9094 17332
rect 10502 17320 10508 17332
rect 10463 17292 10508 17320
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 10689 17323 10747 17329
rect 10689 17289 10701 17323
rect 10735 17320 10747 17323
rect 10873 17323 10931 17329
rect 10873 17320 10885 17323
rect 10735 17292 10885 17320
rect 10735 17289 10747 17292
rect 10689 17283 10747 17289
rect 10873 17289 10885 17292
rect 10919 17320 10931 17323
rect 11054 17320 11060 17332
rect 10919 17292 11060 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11241 17323 11299 17329
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 11514 17320 11520 17332
rect 11287 17292 11520 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 15286 17320 15292 17332
rect 14231 17292 15292 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 16206 17320 16212 17332
rect 16167 17292 16212 17320
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 16669 17323 16727 17329
rect 16669 17289 16681 17323
rect 16715 17320 16727 17323
rect 17494 17320 17500 17332
rect 16715 17292 17500 17320
rect 16715 17289 16727 17292
rect 16669 17283 16727 17289
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 18141 17323 18199 17329
rect 18141 17289 18153 17323
rect 18187 17320 18199 17323
rect 18322 17320 18328 17332
rect 18187 17292 18328 17320
rect 18187 17289 18199 17292
rect 18141 17283 18199 17289
rect 18322 17280 18328 17292
rect 18380 17280 18386 17332
rect 18598 17320 18604 17332
rect 18559 17292 18604 17320
rect 18598 17280 18604 17292
rect 18656 17280 18662 17332
rect 18693 17323 18751 17329
rect 18693 17289 18705 17323
rect 18739 17320 18751 17323
rect 19426 17320 19432 17332
rect 18739 17292 19432 17320
rect 18739 17289 18751 17292
rect 18693 17283 18751 17289
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 19794 17280 19800 17332
rect 19852 17280 19858 17332
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 20220 17292 20545 17320
rect 20220 17280 20226 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 20990 17320 20996 17332
rect 20951 17292 20996 17320
rect 20533 17283 20591 17289
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 21637 17323 21695 17329
rect 21637 17320 21649 17323
rect 21192 17292 21649 17320
rect 4203 17224 4844 17252
rect 4203 17221 4215 17224
rect 4157 17215 4215 17221
rect 4890 17212 4896 17264
rect 4948 17252 4954 17264
rect 5068 17255 5126 17261
rect 5068 17252 5080 17255
rect 4948 17224 5080 17252
rect 4948 17212 4954 17224
rect 5068 17221 5080 17224
rect 5114 17252 5126 17255
rect 5534 17252 5540 17264
rect 5114 17224 5540 17252
rect 5114 17221 5126 17224
rect 5068 17215 5126 17221
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 8938 17252 8944 17264
rect 6236 17224 8944 17252
rect 6236 17212 6242 17224
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4522 17184 4528 17196
rect 4387 17156 4528 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 3712 17048 3740 17147
rect 4522 17144 4528 17156
rect 4580 17144 4586 17196
rect 4709 17188 4767 17193
rect 4632 17187 4767 17188
rect 4632 17160 4721 17187
rect 3973 17119 4031 17125
rect 3973 17085 3985 17119
rect 4019 17116 4031 17119
rect 4632 17116 4660 17160
rect 4709 17153 4721 17160
rect 4755 17153 4767 17187
rect 4709 17147 4767 17153
rect 4019 17088 4660 17116
rect 4019 17085 4031 17088
rect 3973 17079 4031 17085
rect 4798 17076 4804 17128
rect 4856 17116 4862 17128
rect 6822 17116 6828 17128
rect 4856 17088 4901 17116
rect 6783 17088 6828 17116
rect 4856 17076 4862 17088
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 6932 17125 6960 17224
rect 8938 17212 8944 17224
rect 8996 17212 9002 17264
rect 13173 17255 13231 17261
rect 13173 17221 13185 17255
rect 13219 17252 13231 17255
rect 13449 17255 13507 17261
rect 13449 17252 13461 17255
rect 13219 17224 13461 17252
rect 13219 17221 13231 17224
rect 13173 17215 13231 17221
rect 13449 17221 13461 17224
rect 13495 17252 13507 17255
rect 14090 17252 14096 17264
rect 13495 17224 14096 17252
rect 13495 17221 13507 17224
rect 13449 17215 13507 17221
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 7920 17187 7978 17193
rect 7920 17184 7932 17187
rect 7800 17156 7932 17184
rect 7800 17144 7806 17156
rect 7920 17153 7932 17156
rect 7966 17153 7978 17187
rect 9122 17184 9128 17196
rect 9083 17156 9128 17184
rect 7920 17147 7978 17153
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 9381 17187 9439 17193
rect 9381 17184 9393 17187
rect 9232 17156 9393 17184
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17085 6975 17119
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 6917 17079 6975 17085
rect 7392 17088 7665 17116
rect 4154 17048 4160 17060
rect 3712 17020 4160 17048
rect 4154 17008 4160 17020
rect 4212 17008 4218 17060
rect 6365 17051 6423 17057
rect 6365 17048 6377 17051
rect 5736 17020 6377 17048
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4706 16980 4712 16992
rect 4571 16952 4712 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5736 16980 5764 17020
rect 6365 17017 6377 17020
rect 6411 17017 6423 17051
rect 7282 17048 7288 17060
rect 6365 17011 6423 17017
rect 6472 17020 7288 17048
rect 5592 16952 5764 16980
rect 6181 16983 6239 16989
rect 5592 16940 5598 16952
rect 6181 16949 6193 16983
rect 6227 16980 6239 16983
rect 6472 16980 6500 17020
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 6227 16952 6500 16980
rect 6227 16949 6239 16952
rect 6181 16943 6239 16949
rect 6546 16940 6552 16992
rect 6604 16980 6610 16992
rect 7392 16989 7420 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 9030 17076 9036 17128
rect 9088 17116 9094 17128
rect 9232 17116 9260 17156
rect 9381 17153 9393 17156
rect 9427 17153 9439 17187
rect 12710 17184 12716 17196
rect 12768 17193 12774 17196
rect 12680 17156 12716 17184
rect 9381 17147 9439 17153
rect 12710 17144 12716 17156
rect 12768 17147 12780 17193
rect 12986 17184 12992 17196
rect 12899 17156 12992 17184
rect 12768 17144 12774 17147
rect 12986 17144 12992 17156
rect 13044 17184 13050 17196
rect 13188 17184 13216 17215
rect 14090 17212 14096 17224
rect 14148 17252 14154 17264
rect 16390 17252 16396 17264
rect 14148 17224 16396 17252
rect 14148 17212 14154 17224
rect 13044 17156 13216 17184
rect 13633 17187 13691 17193
rect 13044 17144 13050 17156
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13679 17156 13921 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 13909 17153 13921 17156
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 9088 17088 9260 17116
rect 13924 17116 13952 17147
rect 13998 17144 14004 17196
rect 14056 17184 14062 17196
rect 14277 17187 14335 17193
rect 14056 17156 14101 17184
rect 14056 17144 14062 17156
rect 14277 17153 14289 17187
rect 14323 17184 14335 17187
rect 14458 17184 14464 17196
rect 14323 17156 14464 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 14577 17193 14605 17224
rect 16390 17212 16396 17224
rect 16448 17212 16454 17264
rect 17310 17252 17316 17264
rect 16500 17224 17316 17252
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 14642 17144 14648 17196
rect 14700 17184 14706 17196
rect 14809 17187 14867 17193
rect 14809 17184 14821 17187
rect 14700 17156 14821 17184
rect 14700 17144 14706 17156
rect 14809 17153 14821 17156
rect 14855 17153 14867 17187
rect 16022 17184 16028 17196
rect 15983 17156 16028 17184
rect 14809 17147 14867 17153
rect 16022 17144 16028 17156
rect 16080 17144 16086 17196
rect 16500 17184 16528 17224
rect 17310 17212 17316 17224
rect 17368 17212 17374 17264
rect 17770 17212 17776 17264
rect 17828 17261 17834 17264
rect 17828 17252 17840 17261
rect 17828 17224 17873 17252
rect 17828 17215 17840 17224
rect 17828 17212 17834 17215
rect 18782 17212 18788 17264
rect 18840 17252 18846 17264
rect 19812 17252 19840 17280
rect 18840 17224 19840 17252
rect 18840 17212 18846 17224
rect 20070 17212 20076 17264
rect 20128 17252 20134 17264
rect 20714 17252 20720 17264
rect 20128 17224 20720 17252
rect 20128 17212 20134 17224
rect 20714 17212 20720 17224
rect 20772 17252 20778 17264
rect 21192 17252 21220 17292
rect 21637 17289 21649 17292
rect 21683 17320 21695 17323
rect 23014 17320 23020 17332
rect 21683 17292 23020 17320
rect 21683 17289 21695 17292
rect 21637 17283 21695 17289
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 21358 17252 21364 17264
rect 20772 17224 21220 17252
rect 21319 17224 21364 17252
rect 20772 17212 20778 17224
rect 21358 17212 21364 17224
rect 21416 17212 21422 17264
rect 22094 17212 22100 17264
rect 22152 17212 22158 17264
rect 22189 17255 22247 17261
rect 22189 17221 22201 17255
rect 22235 17252 22247 17255
rect 22462 17252 22468 17264
rect 22235 17224 22468 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 22462 17212 22468 17224
rect 22520 17212 22526 17264
rect 18049 17187 18107 17193
rect 16132 17156 16528 17184
rect 17052 17156 18000 17184
rect 16132 17116 16160 17156
rect 13924 17088 14136 17116
rect 9088 17076 9094 17088
rect 10226 17008 10232 17060
rect 10284 17048 10290 17060
rect 11609 17051 11667 17057
rect 11609 17048 11621 17051
rect 10284 17020 11621 17048
rect 10284 17008 10290 17020
rect 11609 17017 11621 17020
rect 11655 17017 11667 17051
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 11609 17011 11667 17017
rect 13096 17020 13737 17048
rect 7193 16983 7251 16989
rect 7193 16980 7205 16983
rect 6604 16952 7205 16980
rect 6604 16940 6610 16952
rect 7193 16949 7205 16952
rect 7239 16980 7251 16983
rect 7377 16983 7435 16989
rect 7377 16980 7389 16983
rect 7239 16952 7389 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7377 16949 7389 16952
rect 7423 16949 7435 16983
rect 7377 16943 7435 16949
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 13096 16980 13124 17020
rect 13725 17017 13737 17020
rect 13771 17017 13783 17051
rect 13725 17011 13783 17017
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 13998 17048 14004 17060
rect 13872 17020 14004 17048
rect 13872 17008 13878 17020
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 11940 16952 13124 16980
rect 14108 16980 14136 17088
rect 15580 17088 16160 17116
rect 16485 17119 16543 17125
rect 14458 17048 14464 17060
rect 14419 17020 14464 17048
rect 14458 17008 14464 17020
rect 14516 17008 14522 17060
rect 15580 16980 15608 17088
rect 16485 17085 16497 17119
rect 16531 17116 16543 17119
rect 16942 17116 16948 17128
rect 16531 17088 16948 17116
rect 16531 17085 16543 17088
rect 16485 17079 16543 17085
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 15654 17008 15660 17060
rect 15712 17048 15718 17060
rect 17052 17048 17080 17156
rect 17972 17116 18000 17156
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18138 17184 18144 17196
rect 18095 17156 18144 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 18322 17184 18328 17196
rect 18283 17156 18328 17184
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17153 18475 17187
rect 18417 17147 18475 17153
rect 18432 17116 18460 17147
rect 19794 17144 19800 17196
rect 19852 17193 19858 17196
rect 19852 17184 19864 17193
rect 19852 17156 19897 17184
rect 19852 17147 19864 17156
rect 19852 17144 19858 17147
rect 19978 17144 19984 17196
rect 20036 17184 20042 17196
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20036 17156 20637 17184
rect 20036 17144 20042 17156
rect 20625 17153 20637 17156
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 22112 17184 22140 17212
rect 21048 17156 22140 17184
rect 22281 17187 22339 17193
rect 21048 17144 21054 17156
rect 22281 17153 22293 17187
rect 22327 17184 22339 17187
rect 22554 17184 22560 17196
rect 22327 17156 22560 17184
rect 22327 17153 22339 17156
rect 22281 17147 22339 17153
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 22741 17187 22799 17193
rect 22741 17153 22753 17187
rect 22787 17184 22799 17187
rect 23290 17184 23296 17196
rect 22787 17156 23296 17184
rect 22787 17153 22799 17156
rect 22741 17147 22799 17153
rect 23290 17144 23296 17156
rect 23348 17144 23354 17196
rect 19058 17116 19064 17128
rect 17972 17088 19064 17116
rect 19058 17076 19064 17088
rect 19116 17076 19122 17128
rect 20070 17116 20076 17128
rect 20031 17088 20076 17116
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 21358 17116 21364 17128
rect 20487 17088 21364 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 22152 17088 22197 17116
rect 22152 17076 22158 17088
rect 15712 17020 17080 17048
rect 15712 17008 15718 17020
rect 18322 17008 18328 17060
rect 18380 17048 18386 17060
rect 18506 17048 18512 17060
rect 18380 17020 18512 17048
rect 18380 17008 18386 17020
rect 18506 17008 18512 17020
rect 18564 17008 18570 17060
rect 20898 17008 20904 17060
rect 20956 17048 20962 17060
rect 21634 17048 21640 17060
rect 20956 17020 21640 17048
rect 20956 17008 20962 17020
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 22922 17048 22928 17060
rect 22883 17020 22928 17048
rect 22922 17008 22928 17020
rect 22980 17008 22986 17060
rect 15930 16980 15936 16992
rect 14108 16952 15608 16980
rect 15891 16952 15936 16980
rect 11940 16940 11946 16952
rect 15930 16940 15936 16952
rect 15988 16940 15994 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16390 16980 16396 16992
rect 16080 16952 16396 16980
rect 16080 16940 16086 16952
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 21082 16980 21088 16992
rect 16724 16952 21088 16980
rect 16724 16940 16730 16952
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21358 16980 21364 16992
rect 21315 16952 21364 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21358 16940 21364 16952
rect 21416 16980 21422 16992
rect 22002 16980 22008 16992
rect 21416 16952 22008 16980
rect 21416 16940 21422 16952
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22649 16983 22707 16989
rect 22649 16949 22661 16983
rect 22695 16980 22707 16983
rect 22738 16980 22744 16992
rect 22695 16952 22744 16980
rect 22695 16949 22707 16952
rect 22649 16943 22707 16949
rect 22738 16940 22744 16952
rect 22796 16940 22802 16992
rect 1104 16890 23460 16912
rect 1104 16838 3749 16890
rect 3801 16838 3813 16890
rect 3865 16838 3877 16890
rect 3929 16838 3941 16890
rect 3993 16838 4005 16890
rect 4057 16838 9347 16890
rect 9399 16838 9411 16890
rect 9463 16838 9475 16890
rect 9527 16838 9539 16890
rect 9591 16838 9603 16890
rect 9655 16838 14945 16890
rect 14997 16838 15009 16890
rect 15061 16838 15073 16890
rect 15125 16838 15137 16890
rect 15189 16838 15201 16890
rect 15253 16838 20543 16890
rect 20595 16838 20607 16890
rect 20659 16838 20671 16890
rect 20723 16838 20735 16890
rect 20787 16838 20799 16890
rect 20851 16838 23460 16890
rect 1104 16816 23460 16838
rect 4154 16776 4160 16788
rect 4115 16748 4160 16776
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 4985 16779 5043 16785
rect 4985 16776 4997 16779
rect 4856 16748 4997 16776
rect 4856 16736 4862 16748
rect 4985 16745 4997 16748
rect 5031 16776 5043 16779
rect 6546 16776 6552 16788
rect 5031 16748 6552 16776
rect 5031 16745 5043 16748
rect 4985 16739 5043 16745
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 12529 16779 12587 16785
rect 12529 16776 12541 16779
rect 9732 16748 12541 16776
rect 9732 16736 9738 16748
rect 12529 16745 12541 16748
rect 12575 16776 12587 16779
rect 12710 16776 12716 16788
rect 12575 16748 12716 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 16206 16776 16212 16788
rect 13004 16748 16212 16776
rect 5166 16708 5172 16720
rect 5127 16680 5172 16708
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 4706 16640 4712 16652
rect 4667 16612 4712 16640
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 6564 16649 6592 16736
rect 11606 16668 11612 16720
rect 11664 16708 11670 16720
rect 13004 16708 13032 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 17770 16736 17776 16788
rect 17828 16776 17834 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 17828 16748 18429 16776
rect 17828 16736 17834 16748
rect 18417 16745 18429 16748
rect 18463 16776 18475 16779
rect 18598 16776 18604 16788
rect 18463 16748 18604 16776
rect 18463 16745 18475 16748
rect 18417 16739 18475 16745
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 20438 16776 20444 16788
rect 18708 16748 20444 16776
rect 14090 16708 14096 16720
rect 11664 16680 13032 16708
rect 14051 16680 14096 16708
rect 11664 16668 11670 16680
rect 14090 16668 14096 16680
rect 14148 16668 14154 16720
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 6595 16612 6653 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 6641 16609 6653 16612
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 8996 16612 9781 16640
rect 8996 16600 9002 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 12360 16612 12868 16640
rect 6270 16532 6276 16584
rect 6328 16581 6334 16584
rect 6328 16572 6340 16581
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 6328 16544 6373 16572
rect 8312 16544 10149 16572
rect 6328 16535 6340 16544
rect 6328 16532 6334 16535
rect 6454 16464 6460 16516
rect 6512 16504 6518 16516
rect 6822 16504 6828 16516
rect 6512 16476 6828 16504
rect 6512 16464 6518 16476
rect 6822 16464 6828 16476
rect 6880 16513 6886 16516
rect 6880 16507 6944 16513
rect 6880 16473 6898 16507
rect 6932 16473 6944 16507
rect 6880 16467 6944 16473
rect 6880 16464 6886 16467
rect 4522 16436 4528 16448
rect 4483 16408 4528 16436
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 4614 16396 4620 16448
rect 4672 16436 4678 16448
rect 8110 16436 8116 16448
rect 4672 16408 4717 16436
rect 8071 16408 8116 16436
rect 4672 16396 4678 16408
rect 8110 16396 8116 16408
rect 8168 16436 8174 16448
rect 8312 16445 8340 16544
rect 10137 16541 10149 16544
rect 10183 16572 10195 16575
rect 11609 16575 11667 16581
rect 11609 16572 11621 16575
rect 10183 16544 11621 16572
rect 10183 16541 10195 16544
rect 10137 16535 10195 16541
rect 11609 16541 11621 16544
rect 11655 16572 11667 16575
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11655 16544 11805 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 11793 16541 11805 16544
rect 11839 16572 11851 16575
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11839 16544 11989 16572
rect 11839 16541 11851 16544
rect 11793 16535 11851 16541
rect 11977 16541 11989 16544
rect 12023 16572 12035 16575
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 12023 16544 12173 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 12161 16541 12173 16544
rect 12207 16572 12219 16575
rect 12360 16572 12388 16612
rect 12207 16544 12388 16572
rect 12840 16572 12868 16612
rect 13909 16575 13967 16581
rect 13909 16572 13921 16575
rect 12840 16544 13921 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 9585 16507 9643 16513
rect 9585 16473 9597 16507
rect 9631 16504 9643 16507
rect 10226 16504 10232 16516
rect 9631 16476 10232 16504
rect 9631 16473 9643 16476
rect 9585 16467 9643 16473
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 10404 16507 10462 16513
rect 10404 16473 10416 16507
rect 10450 16504 10462 16507
rect 10686 16504 10692 16516
rect 10450 16476 10692 16504
rect 10450 16473 10462 16476
rect 10404 16467 10462 16473
rect 10686 16464 10692 16476
rect 10744 16464 10750 16516
rect 12360 16513 12388 16544
rect 13909 16541 13921 16544
rect 13955 16572 13967 16575
rect 15473 16575 15531 16581
rect 15473 16572 15485 16575
rect 13955 16544 15485 16572
rect 13955 16541 13967 16544
rect 13909 16535 13967 16541
rect 15473 16541 15485 16544
rect 15519 16541 15531 16575
rect 15473 16535 15531 16541
rect 12345 16507 12403 16513
rect 12345 16473 12357 16507
rect 12391 16473 12403 16507
rect 12345 16467 12403 16473
rect 13630 16464 13636 16516
rect 13688 16513 13694 16516
rect 13688 16504 13700 16513
rect 14090 16504 14096 16516
rect 13688 16476 14096 16504
rect 13688 16467 13700 16476
rect 13688 16464 13694 16467
rect 14090 16464 14096 16476
rect 14148 16464 14154 16516
rect 14274 16464 14280 16516
rect 14332 16504 14338 16516
rect 15206 16507 15264 16513
rect 15206 16504 15218 16507
rect 14332 16476 15218 16504
rect 14332 16464 14338 16476
rect 15206 16473 15218 16476
rect 15252 16473 15264 16507
rect 15488 16504 15516 16535
rect 16666 16532 16672 16584
rect 16724 16581 16730 16584
rect 16724 16572 16736 16581
rect 16945 16575 17003 16581
rect 16724 16544 16769 16572
rect 16724 16535 16736 16544
rect 16945 16541 16957 16575
rect 16991 16572 17003 16575
rect 17037 16575 17095 16581
rect 17037 16572 17049 16575
rect 16991 16544 17049 16572
rect 16991 16541 17003 16544
rect 16945 16535 17003 16541
rect 17037 16541 17049 16544
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 17304 16575 17362 16581
rect 17304 16541 17316 16575
rect 17350 16572 17362 16575
rect 17586 16572 17592 16584
rect 17350 16544 17592 16572
rect 17350 16541 17362 16544
rect 17304 16535 17362 16541
rect 16724 16532 16730 16535
rect 16574 16504 16580 16516
rect 15488 16476 16580 16504
rect 15206 16467 15264 16473
rect 16574 16464 16580 16476
rect 16632 16504 16638 16516
rect 16960 16504 16988 16535
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16572 18659 16575
rect 18708 16572 18736 16748
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 20625 16779 20683 16785
rect 20625 16745 20637 16779
rect 20671 16776 20683 16779
rect 20898 16776 20904 16788
rect 20671 16748 20904 16776
rect 20671 16745 20683 16748
rect 20625 16739 20683 16745
rect 18785 16711 18843 16717
rect 18785 16677 18797 16711
rect 18831 16677 18843 16711
rect 18785 16671 18843 16677
rect 18647 16544 18736 16572
rect 18800 16572 18828 16671
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18800 16544 18889 16572
rect 18647 16541 18659 16544
rect 18601 16535 18659 16541
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 19242 16572 19248 16584
rect 19203 16544 19248 16572
rect 18877 16535 18935 16541
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 19518 16581 19524 16584
rect 19512 16572 19524 16581
rect 19479 16544 19524 16572
rect 19512 16535 19524 16544
rect 19518 16532 19524 16535
rect 19576 16532 19582 16584
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 20640 16572 20668 16739
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 21545 16779 21603 16785
rect 21545 16745 21557 16779
rect 21591 16745 21603 16779
rect 21545 16739 21603 16745
rect 20993 16643 21051 16649
rect 20993 16609 21005 16643
rect 21039 16640 21051 16643
rect 21358 16640 21364 16652
rect 21039 16612 21364 16640
rect 21039 16609 21051 16612
rect 20993 16603 21051 16609
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 19852 16544 20668 16572
rect 21085 16575 21143 16581
rect 19852 16532 19858 16544
rect 21085 16541 21097 16575
rect 21131 16572 21143 16575
rect 21266 16572 21272 16584
rect 21131 16544 21272 16572
rect 21131 16541 21143 16544
rect 21085 16535 21143 16541
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 21560 16572 21588 16739
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 22244 16748 22477 16776
rect 22244 16736 22250 16748
rect 22465 16745 22477 16748
rect 22511 16745 22523 16779
rect 23014 16776 23020 16788
rect 22975 16748 23020 16776
rect 22465 16739 22523 16745
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 22554 16668 22560 16720
rect 22612 16668 22618 16720
rect 22002 16600 22008 16652
rect 22060 16640 22066 16652
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 22060 16612 22201 16640
rect 22060 16600 22066 16612
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 22572 16640 22600 16668
rect 22572 16612 22968 16640
rect 22189 16603 22247 16609
rect 21560 16544 21956 16572
rect 21928 16516 21956 16544
rect 22554 16532 22560 16584
rect 22612 16572 22618 16584
rect 22940 16581 22968 16612
rect 22649 16575 22707 16581
rect 22649 16572 22661 16575
rect 22612 16544 22661 16572
rect 22612 16532 22618 16544
rect 22649 16541 22661 16544
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 22925 16575 22983 16581
rect 22925 16541 22937 16575
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 20622 16504 20628 16516
rect 16632 16476 16988 16504
rect 17512 16476 20628 16504
rect 16632 16464 16638 16476
rect 8297 16439 8355 16445
rect 8297 16436 8309 16439
rect 8168 16408 8309 16436
rect 8168 16396 8174 16408
rect 8297 16405 8309 16408
rect 8343 16405 8355 16439
rect 9214 16436 9220 16448
rect 9175 16408 9220 16436
rect 8297 16399 8355 16405
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 9674 16436 9680 16448
rect 9635 16408 9680 16436
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 11517 16439 11575 16445
rect 11517 16405 11529 16439
rect 11563 16436 11575 16439
rect 15378 16436 15384 16448
rect 11563 16408 15384 16436
rect 11563 16405 11575 16408
rect 11517 16399 11575 16405
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 15562 16396 15568 16448
rect 15620 16436 15626 16448
rect 17512 16436 17540 16476
rect 20622 16464 20628 16476
rect 20680 16464 20686 16516
rect 21910 16464 21916 16516
rect 21968 16464 21974 16516
rect 15620 16408 17540 16436
rect 19061 16439 19119 16445
rect 15620 16396 15626 16408
rect 19061 16405 19073 16439
rect 19107 16436 19119 16439
rect 20990 16436 20996 16448
rect 19107 16408 20996 16436
rect 19107 16405 19119 16408
rect 19061 16399 19119 16405
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 21177 16439 21235 16445
rect 21177 16405 21189 16439
rect 21223 16436 21235 16439
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 21223 16408 21649 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21637 16405 21649 16408
rect 21683 16405 21695 16439
rect 21637 16399 21695 16405
rect 21726 16396 21732 16448
rect 21784 16436 21790 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 21784 16408 22017 16436
rect 21784 16396 21790 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 22097 16439 22155 16445
rect 22097 16405 22109 16439
rect 22143 16436 22155 16439
rect 22370 16436 22376 16448
rect 22143 16408 22376 16436
rect 22143 16405 22155 16408
rect 22097 16399 22155 16405
rect 22370 16396 22376 16408
rect 22428 16396 22434 16448
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 22741 16439 22799 16445
rect 22741 16436 22753 16439
rect 22704 16408 22753 16436
rect 22704 16396 22710 16408
rect 22741 16405 22753 16408
rect 22787 16405 22799 16439
rect 22741 16399 22799 16405
rect 1104 16346 23460 16368
rect 1104 16294 6548 16346
rect 6600 16294 6612 16346
rect 6664 16294 6676 16346
rect 6728 16294 6740 16346
rect 6792 16294 6804 16346
rect 6856 16294 12146 16346
rect 12198 16294 12210 16346
rect 12262 16294 12274 16346
rect 12326 16294 12338 16346
rect 12390 16294 12402 16346
rect 12454 16294 17744 16346
rect 17796 16294 17808 16346
rect 17860 16294 17872 16346
rect 17924 16294 17936 16346
rect 17988 16294 18000 16346
rect 18052 16294 23460 16346
rect 1104 16272 23460 16294
rect 3602 16192 3608 16244
rect 3660 16232 3666 16244
rect 3973 16235 4031 16241
rect 3973 16232 3985 16235
rect 3660 16204 3985 16232
rect 3660 16192 3666 16204
rect 3973 16201 3985 16204
rect 4019 16201 4031 16235
rect 3973 16195 4031 16201
rect 4341 16235 4399 16241
rect 4341 16201 4353 16235
rect 4387 16232 4399 16235
rect 8481 16235 8539 16241
rect 8481 16232 8493 16235
rect 4387 16204 8493 16232
rect 4387 16201 4399 16204
rect 4341 16195 4399 16201
rect 8481 16201 8493 16204
rect 8527 16201 8539 16235
rect 8481 16195 8539 16201
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 12434 16232 12440 16244
rect 8895 16204 12440 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 12434 16192 12440 16204
rect 12492 16192 12498 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16758 16232 16764 16244
rect 16163 16204 16764 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16758 16192 16764 16204
rect 16816 16232 16822 16244
rect 18049 16235 18107 16241
rect 16816 16204 18000 16232
rect 16816 16192 16822 16204
rect 4522 16164 4528 16176
rect 3712 16136 4528 16164
rect 3712 16105 3740 16136
rect 4522 16124 4528 16136
rect 4580 16124 4586 16176
rect 4798 16124 4804 16176
rect 4856 16164 4862 16176
rect 6914 16164 6920 16176
rect 4856 16136 6920 16164
rect 4856 16124 4862 16136
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 5534 16096 5540 16108
rect 4479 16068 5540 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 3436 16028 3464 16059
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 5902 16056 5908 16108
rect 5960 16105 5966 16108
rect 6196 16105 6224 16136
rect 6914 16124 6920 16136
rect 6972 16164 6978 16176
rect 10781 16167 10839 16173
rect 10781 16164 10793 16167
rect 6972 16136 7880 16164
rect 6972 16124 6978 16136
rect 7852 16105 7880 16136
rect 8128 16136 10793 16164
rect 8128 16108 8156 16136
rect 5960 16096 5972 16105
rect 6181 16099 6239 16105
rect 5960 16068 6005 16096
rect 5960 16059 5972 16068
rect 6181 16065 6193 16099
rect 6227 16065 6239 16099
rect 6181 16059 6239 16065
rect 7581 16099 7639 16105
rect 7581 16065 7593 16099
rect 7627 16096 7639 16099
rect 7837 16099 7895 16105
rect 7627 16068 7788 16096
rect 7627 16065 7639 16068
rect 7581 16059 7639 16065
rect 5960 16056 5966 16059
rect 3436 16000 3740 16028
rect 3510 15920 3516 15972
rect 3568 15960 3574 15972
rect 3605 15963 3663 15969
rect 3605 15960 3617 15963
rect 3568 15932 3617 15960
rect 3568 15920 3574 15932
rect 3605 15929 3617 15932
rect 3651 15929 3663 15963
rect 3712 15960 3740 16000
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 4396 16000 4537 16028
rect 4396 15988 4402 16000
rect 4525 15997 4537 16000
rect 4571 15997 4583 16031
rect 7760 16028 7788 16068
rect 7837 16065 7849 16099
rect 7883 16096 7895 16099
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7883 16068 7941 16096
rect 7883 16065 7895 16068
rect 7837 16059 7895 16065
rect 7929 16065 7941 16068
rect 7975 16096 7987 16099
rect 8110 16096 8116 16108
rect 7975 16068 8116 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 8202 16056 8208 16108
rect 8260 16096 8266 16108
rect 9324 16105 9352 16136
rect 10781 16133 10793 16136
rect 10827 16164 10839 16167
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 10827 16136 11805 16164
rect 10827 16133 10839 16136
rect 10781 16127 10839 16133
rect 11793 16133 11805 16136
rect 11839 16164 11851 16167
rect 11977 16167 12035 16173
rect 11977 16164 11989 16167
rect 11839 16136 11989 16164
rect 11839 16133 11851 16136
rect 11793 16127 11851 16133
rect 11977 16133 11989 16136
rect 12023 16164 12035 16167
rect 12345 16167 12403 16173
rect 12345 16164 12357 16167
rect 12023 16136 12357 16164
rect 12023 16133 12035 16136
rect 11977 16127 12035 16133
rect 12345 16133 12357 16136
rect 12391 16164 12403 16167
rect 12529 16167 12587 16173
rect 12529 16164 12541 16167
rect 12391 16136 12541 16164
rect 12391 16133 12403 16136
rect 12345 16127 12403 16133
rect 12529 16133 12541 16136
rect 12575 16164 12587 16167
rect 14185 16167 14243 16173
rect 14185 16164 14197 16167
rect 12575 16136 14197 16164
rect 12575 16133 12587 16136
rect 12529 16127 12587 16133
rect 9309 16099 9367 16105
rect 8260 16068 9260 16096
rect 8260 16056 8266 16068
rect 8846 16028 8852 16040
rect 7760 16000 8852 16028
rect 4525 15991 4583 15997
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 8941 16031 8999 16037
rect 8941 15997 8953 16031
rect 8987 15997 8999 16031
rect 8941 15991 8999 15997
rect 4614 15960 4620 15972
rect 3712 15932 4620 15960
rect 3605 15923 3663 15929
rect 4614 15920 4620 15932
rect 4672 15920 4678 15972
rect 4801 15963 4859 15969
rect 4801 15929 4813 15963
rect 4847 15960 4859 15963
rect 4890 15960 4896 15972
rect 4847 15932 4896 15960
rect 4847 15929 4859 15932
rect 4801 15923 4859 15929
rect 4890 15920 4896 15932
rect 4948 15920 4954 15972
rect 6362 15920 6368 15972
rect 6420 15960 6426 15972
rect 6457 15963 6515 15969
rect 6457 15960 6469 15963
rect 6420 15932 6469 15960
rect 6420 15920 6426 15932
rect 6457 15929 6469 15932
rect 6503 15929 6515 15963
rect 6457 15923 6515 15929
rect 3881 15895 3939 15901
rect 3881 15861 3893 15895
rect 3927 15892 3939 15895
rect 7650 15892 7656 15904
rect 3927 15864 7656 15892
rect 3927 15861 3939 15864
rect 3881 15855 3939 15861
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 8956 15892 8984 15991
rect 9030 15988 9036 16040
rect 9088 16028 9094 16040
rect 9232 16028 9260 16068
rect 9309 16065 9321 16099
rect 9355 16065 9367 16099
rect 9565 16099 9623 16105
rect 9565 16096 9577 16099
rect 9309 16059 9367 16065
rect 9416 16068 9577 16096
rect 9416 16028 9444 16068
rect 9565 16065 9577 16068
rect 9611 16065 9623 16099
rect 11146 16096 11152 16108
rect 11107 16068 11152 16096
rect 9565 16059 9623 16065
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 11330 16096 11336 16108
rect 11291 16068 11336 16096
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 11422 16056 11428 16108
rect 11480 16096 11486 16108
rect 12728 16105 12756 16136
rect 14185 16133 14197 16136
rect 14231 16164 14243 16167
rect 14369 16167 14427 16173
rect 14369 16164 14381 16167
rect 14231 16136 14381 16164
rect 14231 16133 14243 16136
rect 14185 16127 14243 16133
rect 14369 16133 14381 16136
rect 14415 16133 14427 16167
rect 14369 16127 14427 16133
rect 15004 16167 15062 16173
rect 15004 16133 15016 16167
rect 15050 16164 15062 16167
rect 15562 16164 15568 16176
rect 15050 16136 15568 16164
rect 15050 16133 15062 16136
rect 15004 16127 15062 16133
rect 11609 16099 11667 16105
rect 11609 16096 11621 16099
rect 11480 16068 11621 16096
rect 11480 16056 11486 16068
rect 11609 16065 11621 16068
rect 11655 16065 11667 16099
rect 11609 16059 11667 16065
rect 12713 16099 12771 16105
rect 12713 16065 12725 16099
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 12969 16099 13027 16105
rect 12969 16096 12981 16099
rect 12860 16068 12981 16096
rect 12860 16056 12866 16068
rect 12969 16065 12981 16068
rect 13015 16065 13027 16099
rect 14384 16096 14412 16127
rect 15562 16124 15568 16136
rect 15620 16124 15626 16176
rect 16022 16124 16028 16176
rect 16080 16164 16086 16176
rect 16482 16164 16488 16176
rect 16080 16136 16488 16164
rect 16080 16124 16086 16136
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 16936 16167 16994 16173
rect 16936 16133 16948 16167
rect 16982 16164 16994 16167
rect 17034 16164 17040 16176
rect 16982 16136 17040 16164
rect 16982 16133 16994 16136
rect 16936 16127 16994 16133
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 17972 16164 18000 16204
rect 18049 16201 18061 16235
rect 18095 16232 18107 16235
rect 18230 16232 18236 16244
rect 18095 16204 18236 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 18506 16192 18512 16244
rect 18564 16232 18570 16244
rect 18693 16235 18751 16241
rect 18693 16232 18705 16235
rect 18564 16204 18705 16232
rect 18564 16192 18570 16204
rect 18693 16201 18705 16204
rect 18739 16232 18751 16235
rect 19978 16232 19984 16244
rect 18739 16204 19984 16232
rect 18739 16201 18751 16204
rect 18693 16195 18751 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 20625 16235 20683 16241
rect 20625 16232 20637 16235
rect 20404 16204 20637 16232
rect 20404 16192 20410 16204
rect 20625 16201 20637 16204
rect 20671 16201 20683 16235
rect 20625 16195 20683 16201
rect 20993 16235 21051 16241
rect 20993 16201 21005 16235
rect 21039 16201 21051 16235
rect 20993 16195 21051 16201
rect 19828 16167 19886 16173
rect 17972 16136 18552 16164
rect 14737 16099 14795 16105
rect 14737 16096 14749 16099
rect 14384 16068 14749 16096
rect 12969 16059 13027 16065
rect 14737 16065 14749 16068
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 16301 16099 16359 16105
rect 16301 16096 16313 16099
rect 15804 16068 16313 16096
rect 15804 16056 15810 16068
rect 16301 16065 16313 16068
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16632 16068 16681 16096
rect 16632 16056 16638 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16065 18475 16099
rect 18524 16096 18552 16136
rect 19828 16133 19840 16167
rect 19874 16164 19886 16167
rect 20162 16164 20168 16176
rect 19874 16136 20168 16164
rect 19874 16133 19886 16136
rect 19828 16127 19886 16133
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 21008 16164 21036 16195
rect 21082 16192 21088 16244
rect 21140 16232 21146 16244
rect 21361 16235 21419 16241
rect 21361 16232 21373 16235
rect 21140 16204 21373 16232
rect 21140 16192 21146 16204
rect 21361 16201 21373 16204
rect 21407 16201 21419 16235
rect 21361 16195 21419 16201
rect 21637 16235 21695 16241
rect 21637 16201 21649 16235
rect 21683 16232 21695 16235
rect 22278 16232 22284 16244
rect 21683 16204 22284 16232
rect 21683 16201 21695 16204
rect 21637 16195 21695 16201
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 22554 16232 22560 16244
rect 22515 16204 22560 16232
rect 22554 16192 22560 16204
rect 22612 16192 22618 16244
rect 22189 16167 22247 16173
rect 22189 16164 22201 16167
rect 21008 16136 22201 16164
rect 22189 16133 22201 16136
rect 22235 16133 22247 16167
rect 22370 16164 22376 16176
rect 22189 16127 22247 16133
rect 22296 16136 22376 16164
rect 18524 16068 20668 16096
rect 18417 16059 18475 16065
rect 9088 16000 9133 16028
rect 9232 16000 9444 16028
rect 18325 16031 18383 16037
rect 9088 15988 9094 16000
rect 18325 15997 18337 16031
rect 18371 15997 18383 16031
rect 18432 16028 18460 16059
rect 19058 16028 19064 16040
rect 18432 16000 19064 16028
rect 18325 15991 18383 15997
rect 16482 15960 16488 15972
rect 16443 15932 16488 15960
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 18340 15960 18368 15991
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 20070 16028 20076 16040
rect 20031 16000 20076 16028
rect 20070 15988 20076 16000
rect 20128 15988 20134 16040
rect 20349 16031 20407 16037
rect 20349 15997 20361 16031
rect 20395 15997 20407 16031
rect 20349 15991 20407 15997
rect 18690 15960 18696 15972
rect 18340 15932 18696 15960
rect 18690 15920 18696 15932
rect 18748 15920 18754 15972
rect 20364 15960 20392 15991
rect 20438 15988 20444 16040
rect 20496 16028 20502 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20496 16000 20545 16028
rect 20496 15988 20502 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20640 16028 20668 16068
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21177 16099 21235 16105
rect 21177 16096 21189 16099
rect 20956 16068 21189 16096
rect 20956 16056 20962 16068
rect 21177 16065 21189 16068
rect 21223 16096 21235 16099
rect 21266 16096 21272 16108
rect 21223 16068 21272 16096
rect 21223 16065 21235 16068
rect 21177 16059 21235 16065
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16096 21511 16099
rect 21910 16096 21916 16108
rect 21499 16068 21916 16096
rect 21499 16065 21511 16068
rect 21453 16059 21511 16065
rect 21910 16056 21916 16068
rect 21968 16056 21974 16108
rect 22296 16096 22324 16136
rect 22370 16124 22376 16136
rect 22428 16164 22434 16176
rect 23198 16164 23204 16176
rect 22428 16136 23204 16164
rect 22428 16124 22434 16136
rect 23198 16124 23204 16136
rect 23256 16124 23262 16176
rect 22020 16068 22324 16096
rect 21726 16028 21732 16040
rect 20640 16000 21732 16028
rect 20533 15991 20591 15997
rect 21726 15988 21732 16000
rect 21784 15988 21790 16040
rect 22020 16037 22048 16068
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22520 16068 22845 16096
rect 22520 16056 22526 16068
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 22922 16056 22928 16108
rect 22980 16096 22986 16108
rect 22980 16068 23025 16096
rect 22980 16056 22986 16068
rect 22005 16031 22063 16037
rect 22005 15997 22017 16031
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 22097 16031 22155 16037
rect 22097 15997 22109 16031
rect 22143 16028 22155 16031
rect 22370 16028 22376 16040
rect 22143 16000 22376 16028
rect 22143 15997 22155 16000
rect 22097 15991 22155 15997
rect 22370 15988 22376 16000
rect 22428 15988 22434 16040
rect 21910 15960 21916 15972
rect 20364 15932 21916 15960
rect 21910 15920 21916 15932
rect 21968 15920 21974 15972
rect 22922 15960 22928 15972
rect 22066 15932 22928 15960
rect 10686 15892 10692 15904
rect 8956 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 12250 15892 12256 15904
rect 12211 15864 12256 15892
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 14093 15895 14151 15901
rect 14093 15892 14105 15895
rect 12676 15864 14105 15892
rect 12676 15852 12682 15864
rect 14093 15861 14105 15864
rect 14139 15892 14151 15895
rect 14274 15892 14280 15904
rect 14139 15864 14280 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 14550 15892 14556 15904
rect 14511 15864 14556 15892
rect 14550 15852 14556 15864
rect 14608 15852 14614 15904
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 16666 15892 16672 15904
rect 15160 15864 16672 15892
rect 15160 15852 15166 15864
rect 16666 15852 16672 15864
rect 16724 15892 16730 15904
rect 17310 15892 17316 15904
rect 16724 15864 17316 15892
rect 16724 15852 16730 15864
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 18601 15895 18659 15901
rect 18601 15861 18613 15895
rect 18647 15892 18659 15895
rect 19150 15892 19156 15904
rect 18647 15864 19156 15892
rect 18647 15861 18659 15864
rect 18601 15855 18659 15861
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 22066 15892 22094 15932
rect 22922 15920 22928 15932
rect 22980 15920 22986 15972
rect 19392 15864 22094 15892
rect 19392 15852 19398 15864
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 22649 15895 22707 15901
rect 22649 15892 22661 15895
rect 22520 15864 22661 15892
rect 22520 15852 22526 15864
rect 22649 15861 22661 15864
rect 22695 15861 22707 15895
rect 23106 15892 23112 15904
rect 23067 15864 23112 15892
rect 22649 15855 22707 15861
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 1104 15802 23460 15824
rect 1104 15750 3749 15802
rect 3801 15750 3813 15802
rect 3865 15750 3877 15802
rect 3929 15750 3941 15802
rect 3993 15750 4005 15802
rect 4057 15750 9347 15802
rect 9399 15750 9411 15802
rect 9463 15750 9475 15802
rect 9527 15750 9539 15802
rect 9591 15750 9603 15802
rect 9655 15750 14945 15802
rect 14997 15750 15009 15802
rect 15061 15750 15073 15802
rect 15125 15750 15137 15802
rect 15189 15750 15201 15802
rect 15253 15750 20543 15802
rect 20595 15750 20607 15802
rect 20659 15750 20671 15802
rect 20723 15750 20735 15802
rect 20787 15750 20799 15802
rect 20851 15750 23460 15802
rect 1104 15728 23460 15750
rect 4249 15691 4307 15697
rect 4249 15657 4261 15691
rect 4295 15688 4307 15691
rect 4430 15688 4436 15700
rect 4295 15660 4436 15688
rect 4295 15657 4307 15660
rect 4249 15651 4307 15657
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 5077 15691 5135 15697
rect 5077 15688 5089 15691
rect 4856 15660 5089 15688
rect 4856 15648 4862 15660
rect 5077 15657 5089 15660
rect 5123 15657 5135 15691
rect 5077 15651 5135 15657
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 4801 15555 4859 15561
rect 4801 15552 4813 15555
rect 4396 15524 4813 15552
rect 4396 15512 4402 15524
rect 4801 15521 4813 15524
rect 4847 15521 4859 15555
rect 5092 15552 5120 15651
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 6641 15691 6699 15697
rect 6641 15688 6653 15691
rect 6512 15660 6653 15688
rect 6512 15648 6518 15660
rect 6641 15657 6653 15660
rect 6687 15657 6699 15691
rect 6641 15651 6699 15657
rect 9122 15648 9128 15700
rect 9180 15688 9186 15700
rect 11790 15688 11796 15700
rect 9180 15660 11796 15688
rect 9180 15648 9186 15660
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12802 15688 12808 15700
rect 12492 15660 12808 15688
rect 12492 15648 12498 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 14642 15688 14648 15700
rect 13127 15660 14648 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 15470 15648 15476 15700
rect 15528 15688 15534 15700
rect 15933 15691 15991 15697
rect 15933 15688 15945 15691
rect 15528 15660 15945 15688
rect 15528 15648 15534 15660
rect 15933 15657 15945 15660
rect 15979 15657 15991 15691
rect 16206 15688 16212 15700
rect 16167 15660 16212 15688
rect 15933 15651 15991 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17402 15648 17408 15700
rect 17460 15688 17466 15700
rect 18233 15691 18291 15697
rect 17460 15660 18184 15688
rect 17460 15648 17466 15660
rect 6270 15580 6276 15632
rect 6328 15620 6334 15632
rect 6733 15623 6791 15629
rect 6733 15620 6745 15623
rect 6328 15592 6745 15620
rect 6328 15580 6334 15592
rect 6733 15589 6745 15592
rect 6779 15589 6791 15623
rect 6733 15583 6791 15589
rect 14553 15623 14611 15629
rect 14553 15589 14565 15623
rect 14599 15620 14611 15623
rect 15654 15620 15660 15632
rect 14599 15592 15660 15620
rect 14599 15589 14611 15592
rect 14553 15583 14611 15589
rect 15654 15580 15660 15592
rect 15712 15580 15718 15632
rect 15838 15580 15844 15632
rect 15896 15620 15902 15632
rect 16025 15623 16083 15629
rect 16025 15620 16037 15623
rect 15896 15592 16037 15620
rect 15896 15580 15902 15592
rect 16025 15589 16037 15592
rect 16071 15589 16083 15623
rect 18156 15620 18184 15660
rect 18233 15657 18245 15691
rect 18279 15688 18291 15691
rect 18322 15688 18328 15700
rect 18279 15660 18328 15688
rect 18279 15657 18291 15660
rect 18233 15651 18291 15657
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 19576 15660 20208 15688
rect 19576 15648 19582 15660
rect 20180 15620 20208 15660
rect 20346 15648 20352 15700
rect 20404 15688 20410 15700
rect 20625 15691 20683 15697
rect 20625 15688 20637 15691
rect 20404 15660 20637 15688
rect 20404 15648 20410 15660
rect 20625 15657 20637 15660
rect 20671 15657 20683 15691
rect 21818 15688 21824 15700
rect 20625 15651 20683 15657
rect 21376 15660 21824 15688
rect 20530 15620 20536 15632
rect 18156 15592 18828 15620
rect 20180 15592 20536 15620
rect 16025 15583 16083 15589
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 5092 15524 5273 15552
rect 4801 15515 4859 15521
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 8110 15552 8116 15564
rect 8071 15524 8116 15552
rect 5261 15515 5319 15521
rect 8110 15512 8116 15524
rect 8168 15552 8174 15564
rect 8297 15555 8355 15561
rect 8297 15552 8309 15555
rect 8168 15524 8309 15552
rect 8168 15512 8174 15524
rect 8297 15521 8309 15524
rect 8343 15552 8355 15555
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 8343 15524 8493 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 8481 15521 8493 15524
rect 8527 15552 8539 15555
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 8527 15524 9597 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 8202 15484 8208 15496
rect 4755 15456 8208 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 9600 15484 9628 15515
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 14826 15552 14832 15564
rect 10744 15524 11560 15552
rect 10744 15512 10750 15524
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 9600 15456 11069 15484
rect 11057 15453 11069 15456
rect 11103 15484 11115 15487
rect 11330 15484 11336 15496
rect 11103 15456 11336 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 11330 15444 11336 15456
rect 11388 15484 11394 15496
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11388 15456 11437 15484
rect 11388 15444 11394 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11532 15484 11560 15524
rect 12912 15524 14832 15552
rect 12912 15493 12940 15524
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 15470 15512 15476 15564
rect 15528 15552 15534 15564
rect 15930 15552 15936 15564
rect 15528 15524 15936 15552
rect 15528 15512 15534 15524
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 11681 15487 11739 15493
rect 11681 15484 11693 15487
rect 11532 15456 11693 15484
rect 11425 15447 11483 15453
rect 11681 15453 11693 15456
rect 11727 15453 11739 15487
rect 11681 15447 11739 15453
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 16040 15484 16068 15583
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 18800 15561 18828 15592
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 18288 15524 18705 15552
rect 18288 15512 18294 15524
rect 18693 15521 18705 15524
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15521 18843 15555
rect 19242 15552 19248 15564
rect 19203 15524 19248 15552
rect 18785 15515 18843 15521
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 20993 15555 21051 15561
rect 20993 15521 21005 15555
rect 21039 15552 21051 15555
rect 21266 15552 21272 15564
rect 21039 15524 21272 15552
rect 21039 15521 21051 15524
rect 20993 15515 21051 15521
rect 21266 15512 21272 15524
rect 21324 15512 21330 15564
rect 16393 15487 16451 15493
rect 16393 15484 16405 15487
rect 13587 15456 15976 15484
rect 16040 15456 16405 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 5506 15419 5564 15425
rect 5506 15416 5518 15419
rect 5408 15388 5518 15416
rect 5408 15376 5414 15388
rect 5506 15385 5518 15388
rect 5552 15385 5564 15419
rect 5506 15379 5564 15385
rect 6656 15388 6960 15416
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15348 4675 15351
rect 6656 15348 6684 15388
rect 4663 15320 6684 15348
rect 6932 15348 6960 15388
rect 7742 15376 7748 15428
rect 7800 15416 7806 15428
rect 7846 15419 7904 15425
rect 7846 15416 7858 15419
rect 7800 15388 7858 15416
rect 7800 15376 7806 15388
rect 7846 15385 7858 15388
rect 7892 15385 7904 15419
rect 7846 15379 7904 15385
rect 9306 15376 9312 15428
rect 9364 15416 9370 15428
rect 9830 15419 9888 15425
rect 9830 15416 9842 15419
rect 9364 15388 9842 15416
rect 9364 15376 9370 15388
rect 9830 15385 9842 15388
rect 9876 15385 9888 15419
rect 9830 15379 9888 15385
rect 13265 15419 13323 15425
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13446 15416 13452 15428
rect 13311 15388 13452 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13446 15376 13452 15388
rect 13504 15416 13510 15428
rect 13725 15419 13783 15425
rect 13725 15416 13737 15419
rect 13504 15388 13737 15416
rect 13504 15376 13510 15388
rect 13725 15385 13737 15388
rect 13771 15416 13783 15419
rect 13909 15419 13967 15425
rect 13909 15416 13921 15419
rect 13771 15388 13921 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 13909 15385 13921 15388
rect 13955 15416 13967 15419
rect 14185 15419 14243 15425
rect 14185 15416 14197 15419
rect 13955 15388 14197 15416
rect 13955 15385 13967 15388
rect 13909 15379 13967 15385
rect 14185 15385 14197 15388
rect 14231 15416 14243 15419
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 14231 15388 14381 15416
rect 14231 15385 14243 15388
rect 14185 15379 14243 15385
rect 14369 15385 14381 15388
rect 14415 15416 14427 15419
rect 14737 15419 14795 15425
rect 14737 15416 14749 15419
rect 14415 15388 14749 15416
rect 14415 15385 14427 15388
rect 14369 15379 14427 15385
rect 14737 15385 14749 15388
rect 14783 15416 14795 15419
rect 14921 15419 14979 15425
rect 14921 15416 14933 15419
rect 14783 15388 14933 15416
rect 14783 15385 14795 15388
rect 14737 15379 14795 15385
rect 14921 15385 14933 15388
rect 14967 15416 14979 15419
rect 15105 15419 15163 15425
rect 15105 15416 15117 15419
rect 14967 15388 15117 15416
rect 14967 15385 14979 15388
rect 14921 15379 14979 15385
rect 15105 15385 15117 15388
rect 15151 15416 15163 15419
rect 15654 15416 15660 15428
rect 15151 15388 15660 15416
rect 15151 15385 15163 15388
rect 15105 15379 15163 15385
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 15948 15416 15976 15456
rect 16393 15453 16405 15456
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 16482 15444 16488 15496
rect 16540 15484 16546 15496
rect 16540 15456 16585 15484
rect 16868 15456 18000 15484
rect 16540 15444 16546 15456
rect 16868 15416 16896 15456
rect 15948 15388 16896 15416
rect 16942 15376 16948 15428
rect 17000 15416 17006 15428
rect 17874 15419 17932 15425
rect 17874 15416 17886 15419
rect 17000 15388 17886 15416
rect 17000 15376 17006 15388
rect 17874 15385 17886 15388
rect 17920 15385 17932 15419
rect 17874 15379 17932 15385
rect 9214 15348 9220 15360
rect 6932 15320 9220 15348
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 10778 15308 10784 15360
rect 10836 15348 10842 15360
rect 10965 15351 11023 15357
rect 10965 15348 10977 15351
rect 10836 15320 10977 15348
rect 10836 15308 10842 15320
rect 10965 15317 10977 15320
rect 11011 15317 11023 15351
rect 15562 15348 15568 15360
rect 15523 15320 15568 15348
rect 10965 15311 11023 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 16666 15348 16672 15360
rect 16627 15320 16672 15348
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 16761 15351 16819 15357
rect 16761 15317 16773 15351
rect 16807 15348 16819 15351
rect 17034 15348 17040 15360
rect 16807 15320 17040 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17972 15348 18000 15456
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 19260 15484 19288 15512
rect 21376 15484 21404 15660
rect 21818 15648 21824 15660
rect 21876 15648 21882 15700
rect 22370 15688 22376 15700
rect 22331 15660 22376 15688
rect 22370 15648 22376 15660
rect 22428 15648 22434 15700
rect 22002 15620 22008 15632
rect 21744 15592 22008 15620
rect 21744 15561 21772 15592
rect 22002 15580 22008 15592
rect 22060 15580 22066 15632
rect 22094 15580 22100 15632
rect 22152 15620 22158 15632
rect 22465 15623 22523 15629
rect 22465 15620 22477 15623
rect 22152 15592 22477 15620
rect 22152 15580 22158 15592
rect 22465 15589 22477 15592
rect 22511 15589 22523 15623
rect 22465 15583 22523 15589
rect 21729 15555 21787 15561
rect 21729 15521 21741 15555
rect 21775 15521 21787 15555
rect 21729 15515 21787 15521
rect 21818 15512 21824 15564
rect 21876 15552 21882 15564
rect 23017 15555 23075 15561
rect 23017 15552 23029 15555
rect 21876 15524 23029 15552
rect 21876 15512 21882 15524
rect 23017 15521 23029 15524
rect 23063 15521 23075 15555
rect 23017 15515 23075 15521
rect 18196 15456 19288 15484
rect 19444 15456 21404 15484
rect 18196 15444 18202 15456
rect 18598 15416 18604 15428
rect 18559 15388 18604 15416
rect 18598 15376 18604 15388
rect 18656 15376 18662 15428
rect 19058 15376 19064 15428
rect 19116 15416 19122 15428
rect 19444 15416 19472 15456
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 22649 15487 22707 15493
rect 22649 15484 22661 15487
rect 21692 15456 22661 15484
rect 21692 15444 21698 15456
rect 22649 15453 22661 15456
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 22738 15444 22744 15496
rect 22796 15484 22802 15496
rect 22925 15487 22983 15493
rect 22925 15484 22937 15487
rect 22796 15456 22937 15484
rect 22796 15444 22802 15456
rect 22925 15453 22937 15456
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 19116 15388 19472 15416
rect 19512 15419 19570 15425
rect 19116 15376 19122 15388
rect 19512 15385 19524 15419
rect 19558 15416 19570 15419
rect 20438 15416 20444 15428
rect 19558 15388 20444 15416
rect 19558 15385 19570 15388
rect 19512 15379 19570 15385
rect 20438 15376 20444 15388
rect 20496 15376 20502 15428
rect 20530 15376 20536 15428
rect 20588 15416 20594 15428
rect 22005 15419 22063 15425
rect 22005 15416 22017 15419
rect 20588 15388 22017 15416
rect 20588 15376 20594 15388
rect 22005 15385 22017 15388
rect 22051 15385 22063 15419
rect 22005 15379 22063 15385
rect 20898 15348 20904 15360
rect 17972 15320 20904 15348
rect 20898 15308 20904 15320
rect 20956 15308 20962 15360
rect 21082 15348 21088 15360
rect 21043 15320 21088 15348
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 21545 15351 21603 15357
rect 21232 15320 21277 15348
rect 21232 15308 21238 15320
rect 21545 15317 21557 15351
rect 21591 15348 21603 15351
rect 21818 15348 21824 15360
rect 21591 15320 21824 15348
rect 21591 15317 21603 15320
rect 21545 15311 21603 15317
rect 21818 15308 21824 15320
rect 21876 15308 21882 15360
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22738 15348 22744 15360
rect 21968 15320 22013 15348
rect 22699 15320 22744 15348
rect 21968 15308 21974 15320
rect 22738 15308 22744 15320
rect 22796 15308 22802 15360
rect 1104 15258 23460 15280
rect 1104 15206 6548 15258
rect 6600 15206 6612 15258
rect 6664 15206 6676 15258
rect 6728 15206 6740 15258
rect 6792 15206 6804 15258
rect 6856 15206 12146 15258
rect 12198 15206 12210 15258
rect 12262 15206 12274 15258
rect 12326 15206 12338 15258
rect 12390 15206 12402 15258
rect 12454 15206 17744 15258
rect 17796 15206 17808 15258
rect 17860 15206 17872 15258
rect 17924 15206 17936 15258
rect 17988 15206 18000 15258
rect 18052 15206 23460 15258
rect 1104 15184 23460 15206
rect 5074 15104 5080 15156
rect 5132 15144 5138 15156
rect 5132 15116 8156 15144
rect 5132 15104 5138 15116
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 7092 15079 7150 15085
rect 7092 15076 7104 15079
rect 5776 15048 7104 15076
rect 5776 15036 5782 15048
rect 7092 15045 7104 15048
rect 7138 15076 7150 15079
rect 7374 15076 7380 15088
rect 7138 15048 7380 15076
rect 7138 15045 7150 15048
rect 7092 15039 7150 15045
rect 7374 15036 7380 15048
rect 7432 15036 7438 15088
rect 4890 15008 4896 15020
rect 4851 14980 4896 15008
rect 4890 14968 4896 14980
rect 4948 14968 4954 15020
rect 5626 15008 5632 15020
rect 5539 14980 5632 15008
rect 5626 14968 5632 14980
rect 5684 15008 5690 15020
rect 6270 15008 6276 15020
rect 5684 14980 6276 15008
rect 5684 14968 5690 14980
rect 6270 14968 6276 14980
rect 6328 15008 6334 15020
rect 6457 15011 6515 15017
rect 6457 15008 6469 15011
rect 6328 14980 6469 15008
rect 6328 14968 6334 14980
rect 6457 14977 6469 14980
rect 6503 14977 6515 15011
rect 6457 14971 6515 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 6914 15008 6920 15020
rect 6871 14980 6920 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 8128 15008 8156 15116
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 8260 15116 8401 15144
rect 8260 15104 8266 15116
rect 8389 15113 8401 15116
rect 8435 15113 8447 15147
rect 8389 15107 8447 15113
rect 8757 15147 8815 15153
rect 8757 15113 8769 15147
rect 8803 15144 8815 15147
rect 8803 15116 11753 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 8849 15079 8907 15085
rect 8849 15045 8861 15079
rect 8895 15076 8907 15079
rect 11725 15076 11753 15116
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 11848 15116 12909 15144
rect 11848 15104 11854 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 12897 15107 12955 15113
rect 13173 15147 13231 15153
rect 13173 15113 13185 15147
rect 13219 15144 13231 15147
rect 13446 15144 13452 15156
rect 13219 15116 13452 15144
rect 13219 15113 13231 15116
rect 13173 15107 13231 15113
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 14369 15147 14427 15153
rect 14369 15113 14381 15147
rect 14415 15144 14427 15147
rect 15562 15144 15568 15156
rect 14415 15116 15568 15144
rect 14415 15113 14427 15116
rect 14369 15107 14427 15113
rect 13630 15076 13636 15088
rect 8895 15048 11652 15076
rect 11725 15048 13636 15076
rect 8895 15045 8907 15048
rect 8849 15039 8907 15045
rect 10778 15008 10784 15020
rect 8128 14980 10784 15008
rect 10778 14968 10784 14980
rect 10836 15008 10842 15020
rect 11066 15011 11124 15017
rect 11066 15008 11078 15011
rect 10836 14980 11078 15008
rect 10836 14968 10842 14980
rect 11066 14977 11078 14980
rect 11112 14977 11124 15011
rect 11330 15008 11336 15020
rect 11291 14980 11336 15008
rect 11066 14971 11124 14977
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5534 14940 5540 14952
rect 5399 14912 5540 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 5534 14900 5540 14912
rect 5592 14940 5598 14952
rect 5902 14940 5908 14952
rect 5592 14912 5908 14940
rect 5592 14900 5598 14912
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 9030 14940 9036 14952
rect 8991 14912 9036 14940
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9953 14875 10011 14881
rect 9953 14872 9965 14875
rect 7760 14844 9965 14872
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 5077 14807 5135 14813
rect 5077 14804 5089 14807
rect 4764 14776 5089 14804
rect 4764 14764 4770 14776
rect 5077 14773 5089 14776
rect 5123 14773 5135 14807
rect 5077 14767 5135 14773
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6420 14776 6561 14804
rect 6420 14764 6426 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 7760 14804 7788 14844
rect 9953 14841 9965 14844
rect 9999 14841 10011 14875
rect 9953 14835 10011 14841
rect 8202 14804 8208 14816
rect 6696 14776 7788 14804
rect 8163 14776 8208 14804
rect 6696 14764 6702 14776
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 11112 14776 11529 14804
rect 11112 14764 11118 14776
rect 11517 14773 11529 14776
rect 11563 14773 11575 14807
rect 11624 14804 11652 15048
rect 13630 15036 13636 15048
rect 13688 15036 13694 15088
rect 11882 15008 11888 15020
rect 11843 14980 11888 15008
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 14384 15008 14412 15107
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 19334 15144 19340 15156
rect 17276 15116 19340 15144
rect 17276 15104 17282 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 21634 15144 21640 15156
rect 19444 15116 21404 15144
rect 21595 15116 21640 15144
rect 16684 15048 18184 15076
rect 14323 14980 14412 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 15470 14968 15476 15020
rect 15528 15017 15534 15020
rect 15528 15008 15540 15017
rect 15528 14980 15573 15008
rect 15528 14971 15540 14980
rect 15528 14968 15534 14971
rect 15654 14968 15660 15020
rect 15712 15008 15718 15020
rect 15749 15011 15807 15017
rect 15749 15008 15761 15011
rect 15712 14980 15761 15008
rect 15712 14968 15718 14980
rect 15749 14977 15761 14980
rect 15795 15008 15807 15011
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 15795 14980 15945 15008
rect 15795 14977 15807 14980
rect 15749 14971 15807 14977
rect 15933 14977 15945 14980
rect 15979 15008 15991 15011
rect 16206 15008 16212 15020
rect 15979 14980 16212 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16206 14968 16212 14980
rect 16264 15008 16270 15020
rect 16684 15017 16712 15048
rect 18156 15020 18184 15048
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 16264 14980 16313 15008
rect 16264 14968 16270 14980
rect 16301 14977 16313 14980
rect 16347 15008 16359 15011
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16347 14980 16681 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16925 15011 16983 15017
rect 16925 15008 16937 15011
rect 16816 14980 16937 15008
rect 16816 14968 16822 14980
rect 16925 14977 16937 14980
rect 16971 14977 16983 15011
rect 18138 15008 18144 15020
rect 18099 14980 18144 15008
rect 16925 14971 16983 14977
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18408 15011 18466 15017
rect 18408 15008 18420 15011
rect 18248 14980 18420 15008
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11848 14912 11989 14940
rect 11848 14900 11854 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12434 14940 12440 14952
rect 12207 14912 12440 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 18248 14940 18276 14980
rect 18408 14977 18420 14980
rect 18454 15008 18466 15011
rect 19444 15008 19472 15116
rect 21269 15079 21327 15085
rect 21269 15076 21281 15079
rect 18454 14980 19472 15008
rect 19536 15048 21281 15076
rect 18454 14977 18466 14980
rect 18408 14971 18466 14977
rect 18064 14912 18276 14940
rect 15838 14832 15844 14884
rect 15896 14872 15902 14884
rect 16393 14875 16451 14881
rect 16393 14872 16405 14875
rect 15896 14844 16405 14872
rect 15896 14832 15902 14844
rect 16393 14841 16405 14844
rect 16439 14872 16451 14875
rect 16482 14872 16488 14884
rect 16439 14844 16488 14872
rect 16439 14841 16451 14844
rect 16393 14835 16451 14841
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 18064 14881 18092 14912
rect 19150 14900 19156 14952
rect 19208 14940 19214 14952
rect 19536 14940 19564 15048
rect 21269 15045 21281 15048
rect 21315 15045 21327 15079
rect 21376 15076 21404 15116
rect 21634 15104 21640 15116
rect 21692 15104 21698 15156
rect 22462 15144 22468 15156
rect 22423 15116 22468 15144
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 22557 15147 22615 15153
rect 22557 15113 22569 15147
rect 22603 15144 22615 15147
rect 22738 15144 22744 15156
rect 22603 15116 22744 15144
rect 22603 15113 22615 15116
rect 22557 15107 22615 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 21910 15076 21916 15088
rect 21376 15048 21916 15076
rect 21269 15039 21327 15045
rect 21910 15036 21916 15048
rect 21968 15036 21974 15088
rect 19610 14968 19616 15020
rect 19668 15008 19674 15020
rect 20726 15011 20784 15017
rect 20726 15008 20738 15011
rect 19668 14980 20738 15008
rect 19668 14968 19674 14980
rect 20726 14977 20738 14980
rect 20772 15008 20784 15011
rect 21453 15011 21511 15017
rect 21453 15008 21465 15011
rect 20772 14980 21465 15008
rect 20772 14977 20784 14980
rect 20726 14971 20784 14977
rect 21453 14977 21465 14980
rect 21499 14977 21511 15011
rect 21453 14971 21511 14977
rect 21726 14968 21732 15020
rect 21784 15008 21790 15020
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21784 14980 21833 15008
rect 21784 14968 21790 14980
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 23198 15008 23204 15020
rect 23155 14980 23204 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 19208 14912 19564 14940
rect 20993 14943 21051 14949
rect 19208 14900 19214 14912
rect 20993 14909 21005 14943
rect 21039 14909 21051 14943
rect 20993 14903 21051 14909
rect 18049 14875 18107 14881
rect 18049 14841 18061 14875
rect 18095 14841 18107 14875
rect 19518 14872 19524 14884
rect 19479 14844 19524 14872
rect 18049 14835 18107 14841
rect 19518 14832 19524 14844
rect 19576 14832 19582 14884
rect 12618 14804 12624 14816
rect 11624 14776 12624 14804
rect 11517 14767 11575 14773
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 12802 14804 12808 14816
rect 12763 14776 12808 14804
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 13262 14804 13268 14816
rect 13223 14776 13268 14804
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 13412 14776 13645 14804
rect 13412 14764 13418 14776
rect 13633 14773 13645 14776
rect 13679 14773 13691 14807
rect 13633 14767 13691 14773
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 15804 14776 16037 14804
rect 15804 14764 15810 14776
rect 16025 14773 16037 14776
rect 16071 14773 16083 14807
rect 16025 14767 16083 14773
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 19334 14804 19340 14816
rect 16172 14776 19340 14804
rect 16172 14764 16178 14776
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19613 14807 19671 14813
rect 19613 14804 19625 14807
rect 19484 14776 19625 14804
rect 19484 14764 19490 14776
rect 19613 14773 19625 14776
rect 19659 14773 19671 14807
rect 19613 14767 19671 14773
rect 20070 14764 20076 14816
rect 20128 14804 20134 14816
rect 21008 14804 21036 14903
rect 21082 14900 21088 14952
rect 21140 14940 21146 14952
rect 22649 14943 22707 14949
rect 21140 14912 22094 14940
rect 21140 14900 21146 14912
rect 22066 14872 22094 14912
rect 22649 14909 22661 14943
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 22664 14872 22692 14903
rect 22066 14844 22692 14872
rect 21085 14807 21143 14813
rect 21085 14804 21097 14807
rect 20128 14776 21097 14804
rect 20128 14764 20134 14776
rect 21085 14773 21097 14776
rect 21131 14804 21143 14807
rect 21542 14804 21548 14816
rect 21131 14776 21548 14804
rect 21131 14773 21143 14776
rect 21085 14767 21143 14773
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 22002 14804 22008 14816
rect 21963 14776 22008 14804
rect 22002 14764 22008 14776
rect 22060 14764 22066 14816
rect 22097 14807 22155 14813
rect 22097 14773 22109 14807
rect 22143 14804 22155 14807
rect 22462 14804 22468 14816
rect 22143 14776 22468 14804
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 22925 14807 22983 14813
rect 22925 14773 22937 14807
rect 22971 14804 22983 14807
rect 23014 14804 23020 14816
rect 22971 14776 23020 14804
rect 22971 14773 22983 14776
rect 22925 14767 22983 14773
rect 23014 14764 23020 14776
rect 23072 14764 23078 14816
rect 1104 14714 23460 14736
rect 1104 14662 3749 14714
rect 3801 14662 3813 14714
rect 3865 14662 3877 14714
rect 3929 14662 3941 14714
rect 3993 14662 4005 14714
rect 4057 14662 9347 14714
rect 9399 14662 9411 14714
rect 9463 14662 9475 14714
rect 9527 14662 9539 14714
rect 9591 14662 9603 14714
rect 9655 14662 14945 14714
rect 14997 14662 15009 14714
rect 15061 14662 15073 14714
rect 15125 14662 15137 14714
rect 15189 14662 15201 14714
rect 15253 14662 20543 14714
rect 20595 14662 20607 14714
rect 20659 14662 20671 14714
rect 20723 14662 20735 14714
rect 20787 14662 20799 14714
rect 20851 14662 23460 14714
rect 1104 14640 23460 14662
rect 5626 14600 5632 14612
rect 5276 14572 5632 14600
rect 5074 14464 5080 14476
rect 5035 14436 5080 14464
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5276 14473 5304 14572
rect 5626 14560 5632 14572
rect 5684 14560 5690 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 6917 14603 6975 14609
rect 6917 14600 6929 14603
rect 5868 14572 6929 14600
rect 5868 14560 5874 14572
rect 6917 14569 6929 14572
rect 6963 14600 6975 14603
rect 7006 14600 7012 14612
rect 6963 14572 7012 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8168 14572 8401 14600
rect 8168 14560 8174 14572
rect 8312 14473 8340 14572
rect 8389 14569 8401 14572
rect 8435 14600 8447 14603
rect 8573 14603 8631 14609
rect 8573 14600 8585 14603
rect 8435 14572 8585 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 8573 14569 8585 14572
rect 8619 14569 8631 14603
rect 11330 14600 11336 14612
rect 11291 14572 11336 14600
rect 8573 14563 8631 14569
rect 8588 14532 8616 14563
rect 11330 14560 11336 14572
rect 11388 14600 11394 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 11388 14572 11437 14600
rect 11388 14560 11394 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11606 14600 11612 14612
rect 11567 14572 11612 14600
rect 11425 14563 11483 14569
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 16942 14600 16948 14612
rect 12860 14572 16804 14600
rect 16903 14572 16948 14600
rect 12860 14560 12866 14572
rect 9674 14532 9680 14544
rect 8588 14504 9680 14532
rect 9674 14492 9680 14504
rect 9732 14532 9738 14544
rect 11149 14535 11207 14541
rect 9732 14504 9812 14532
rect 9732 14492 9738 14504
rect 9784 14473 9812 14504
rect 11149 14501 11161 14535
rect 11195 14532 11207 14535
rect 11882 14532 11888 14544
rect 11195 14504 11888 14532
rect 11195 14501 11207 14504
rect 11149 14495 11207 14501
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 16206 14532 16212 14544
rect 16132 14504 16212 14532
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14433 5319 14467
rect 5261 14427 5319 14433
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14433 9827 14467
rect 13354 14464 13360 14476
rect 9769 14427 9827 14433
rect 12912 14436 13360 14464
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 6914 14396 6920 14408
rect 5491 14368 6920 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 6914 14356 6920 14368
rect 6972 14356 6978 14408
rect 9600 14396 9628 14427
rect 10318 14396 10324 14408
rect 9600 14368 10324 14396
rect 10318 14356 10324 14368
rect 10376 14396 10382 14408
rect 12434 14396 12440 14408
rect 10376 14368 12020 14396
rect 10376 14356 10382 14368
rect 4985 14331 5043 14337
rect 4985 14297 4997 14331
rect 5031 14328 5043 14331
rect 5712 14331 5770 14337
rect 5712 14328 5724 14331
rect 5031 14300 5724 14328
rect 5031 14297 5043 14300
rect 4985 14291 5043 14297
rect 5712 14297 5724 14300
rect 5758 14328 5770 14331
rect 6638 14328 6644 14340
rect 5758 14300 6644 14328
rect 5758 14297 5770 14300
rect 5712 14291 5770 14297
rect 6638 14288 6644 14300
rect 6696 14288 6702 14340
rect 8030 14331 8088 14337
rect 8030 14328 8042 14331
rect 6840 14300 8042 14328
rect 4617 14263 4675 14269
rect 4617 14229 4629 14263
rect 4663 14260 4675 14263
rect 4890 14260 4896 14272
rect 4663 14232 4896 14260
rect 4663 14229 4675 14232
rect 4617 14223 4675 14229
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 5810 14260 5816 14272
rect 5132 14232 5816 14260
rect 5132 14220 5138 14232
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6454 14220 6460 14272
rect 6512 14260 6518 14272
rect 6840 14269 6868 14300
rect 8030 14297 8042 14300
rect 8076 14297 8088 14331
rect 8030 14291 8088 14297
rect 9309 14331 9367 14337
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 9766 14328 9772 14340
rect 9355 14300 9772 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 10036 14331 10094 14337
rect 10036 14297 10048 14331
rect 10082 14328 10094 14331
rect 10082 14300 11284 14328
rect 10082 14297 10094 14300
rect 10036 14291 10094 14297
rect 11256 14272 11284 14300
rect 11422 14288 11428 14340
rect 11480 14328 11486 14340
rect 11992 14328 12020 14368
rect 12360 14368 12440 14396
rect 12360 14328 12388 14368
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 12733 14399 12791 14405
rect 12733 14365 12745 14399
rect 12779 14396 12791 14399
rect 12912 14396 12940 14436
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13722 14464 13728 14476
rect 13683 14436 13728 14464
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 16132 14473 16160 14504
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 16776 14532 16804 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 17586 14600 17592 14612
rect 17420 14572 17592 14600
rect 17420 14532 17448 14572
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 18196 14572 18429 14600
rect 18196 14560 18202 14572
rect 16776 14504 17448 14532
rect 18340 14473 18368 14572
rect 18417 14569 18429 14572
rect 18463 14569 18475 14603
rect 18782 14600 18788 14612
rect 18743 14572 18788 14600
rect 18417 14563 18475 14569
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 19484 14572 20392 14600
rect 19484 14560 19490 14572
rect 18874 14532 18880 14544
rect 18835 14504 18880 14532
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 20364 14532 20392 14572
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 20625 14603 20683 14609
rect 20625 14600 20637 14603
rect 20496 14572 20637 14600
rect 20496 14560 20502 14572
rect 20625 14569 20637 14572
rect 20671 14569 20683 14603
rect 20625 14563 20683 14569
rect 21082 14532 21088 14544
rect 20364 14504 21088 14532
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 21821 14535 21879 14541
rect 21821 14501 21833 14535
rect 21867 14532 21879 14535
rect 22738 14532 22744 14544
rect 21867 14504 22744 14532
rect 21867 14501 21879 14504
rect 21821 14495 21879 14501
rect 22738 14492 22744 14504
rect 22796 14492 22802 14544
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 18325 14467 18383 14473
rect 18325 14433 18337 14467
rect 18371 14464 18383 14467
rect 19245 14467 19303 14473
rect 19245 14464 19257 14467
rect 18371 14436 19257 14464
rect 18371 14433 18383 14436
rect 18325 14427 18383 14433
rect 19245 14433 19257 14436
rect 19291 14433 19303 14467
rect 21266 14464 21272 14476
rect 21227 14436 21272 14464
rect 19245 14427 19303 14433
rect 21266 14424 21272 14436
rect 21324 14424 21330 14476
rect 22462 14464 22468 14476
rect 22423 14436 22468 14464
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 22557 14467 22615 14473
rect 22557 14433 22569 14467
rect 22603 14433 22615 14467
rect 22557 14427 22615 14433
rect 12779 14368 12940 14396
rect 12989 14399 13047 14405
rect 12779 14365 12791 14368
rect 12733 14359 12791 14365
rect 12989 14365 13001 14399
rect 13035 14396 13047 14399
rect 14274 14396 14280 14408
rect 13035 14368 14280 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 14274 14356 14280 14368
rect 14332 14396 14338 14408
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 14332 14368 14381 14396
rect 14332 14356 14338 14368
rect 14369 14365 14381 14368
rect 14415 14396 14427 14399
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14415 14368 14565 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17310 14396 17316 14408
rect 16807 14368 17316 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 18601 14399 18659 14405
rect 18601 14365 18613 14399
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14396 19119 14399
rect 19150 14396 19156 14408
rect 19107 14368 19156 14396
rect 19107 14365 19119 14368
rect 19061 14359 19119 14365
rect 12894 14328 12900 14340
rect 11480 14300 11928 14328
rect 11992 14300 12900 14328
rect 11480 14288 11486 14300
rect 6825 14263 6883 14269
rect 6825 14260 6837 14263
rect 6512 14232 6837 14260
rect 6512 14220 6518 14232
rect 6825 14229 6837 14232
rect 6871 14229 6883 14263
rect 8938 14260 8944 14272
rect 8899 14232 8944 14260
rect 6825 14223 6883 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9401 14263 9459 14269
rect 9401 14229 9413 14263
rect 9447 14260 9459 14263
rect 10962 14260 10968 14272
rect 9447 14232 10968 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11790 14260 11796 14272
rect 11296 14232 11796 14260
rect 11296 14220 11302 14232
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 11900 14260 11928 14300
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13630 14328 13636 14340
rect 13543 14300 13636 14328
rect 13630 14288 13636 14300
rect 13688 14328 13694 14340
rect 15470 14328 15476 14340
rect 13688 14300 15476 14328
rect 13688 14288 13694 14300
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 15850 14331 15908 14337
rect 15850 14297 15862 14331
rect 15896 14328 15908 14331
rect 15896 14300 17172 14328
rect 15896 14297 15908 14300
rect 15850 14291 15908 14297
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 11900 14232 13185 14260
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 13173 14223 13231 14229
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14260 13599 14263
rect 14642 14260 14648 14272
rect 13587 14232 14648 14260
rect 13587 14229 13599 14232
rect 13541 14223 13599 14229
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 14737 14263 14795 14269
rect 14737 14229 14749 14263
rect 14783 14260 14795 14263
rect 15194 14260 15200 14272
rect 14783 14232 15200 14260
rect 14783 14229 14795 14232
rect 14737 14223 14795 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 15378 14220 15384 14272
rect 15436 14260 15442 14272
rect 15856 14260 15884 14291
rect 16482 14260 16488 14272
rect 15436 14232 15884 14260
rect 16443 14232 16488 14260
rect 15436 14220 15442 14232
rect 16482 14220 16488 14232
rect 16540 14220 16546 14272
rect 16666 14260 16672 14272
rect 16627 14232 16672 14260
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 17144 14260 17172 14300
rect 17218 14288 17224 14340
rect 17276 14328 17282 14340
rect 18058 14331 18116 14337
rect 18058 14328 18070 14331
rect 17276 14300 18070 14328
rect 17276 14288 17282 14300
rect 18058 14297 18070 14300
rect 18104 14297 18116 14331
rect 18616 14328 18644 14359
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 19518 14405 19524 14408
rect 19512 14396 19524 14405
rect 19479 14368 19524 14396
rect 19512 14359 19524 14368
rect 19518 14356 19524 14359
rect 19576 14356 19582 14408
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 21545 14399 21603 14405
rect 21545 14396 21557 14399
rect 21508 14368 21557 14396
rect 21508 14356 21514 14368
rect 21545 14365 21557 14368
rect 21591 14365 21603 14399
rect 21545 14359 21603 14365
rect 21634 14356 21640 14408
rect 21692 14396 21698 14408
rect 21692 14368 21737 14396
rect 21692 14356 21698 14368
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22572 14396 22600 14427
rect 23014 14396 23020 14408
rect 22152 14368 22600 14396
rect 22975 14368 23020 14396
rect 22152 14356 22158 14368
rect 23014 14356 23020 14368
rect 23072 14356 23078 14408
rect 19886 14328 19892 14340
rect 18616 14300 19892 14328
rect 18058 14291 18116 14297
rect 19886 14288 19892 14300
rect 19944 14288 19950 14340
rect 22462 14328 22468 14340
rect 22020 14300 22468 14328
rect 21174 14260 21180 14272
rect 17144 14232 21180 14260
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 22020 14269 22048 14300
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 22005 14263 22063 14269
rect 22005 14229 22017 14263
rect 22051 14229 22063 14263
rect 22370 14260 22376 14272
rect 22331 14232 22376 14260
rect 22005 14223 22063 14229
rect 22370 14220 22376 14232
rect 22428 14220 22434 14272
rect 22922 14260 22928 14272
rect 22883 14232 22928 14260
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 1104 14170 23460 14192
rect 1104 14118 6548 14170
rect 6600 14118 6612 14170
rect 6664 14118 6676 14170
rect 6728 14118 6740 14170
rect 6792 14118 6804 14170
rect 6856 14118 12146 14170
rect 12198 14118 12210 14170
rect 12262 14118 12274 14170
rect 12326 14118 12338 14170
rect 12390 14118 12402 14170
rect 12454 14118 17744 14170
rect 17796 14118 17808 14170
rect 17860 14118 17872 14170
rect 17924 14118 17936 14170
rect 17988 14118 18000 14170
rect 18052 14118 23460 14170
rect 1104 14096 23460 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1728 14028 1869 14056
rect 1728 14016 1734 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 1857 14019 1915 14025
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 6454 14056 6460 14068
rect 4755 14028 6460 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 6454 14016 6460 14028
rect 6512 14016 6518 14068
rect 6914 14016 6920 14068
rect 6972 14016 6978 14068
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 11238 14056 11244 14068
rect 11199 14028 11244 14056
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11388 14028 11529 14056
rect 11388 14016 11394 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 13630 14056 13636 14068
rect 13219 14028 13636 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 4801 13991 4859 13997
rect 4801 13957 4813 13991
rect 4847 13988 4859 13991
rect 5074 13988 5080 14000
rect 4847 13960 5080 13988
rect 4847 13957 4859 13960
rect 4801 13951 4859 13957
rect 5074 13948 5080 13960
rect 5132 13948 5138 14000
rect 6932 13988 6960 14016
rect 6656 13960 6960 13988
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13889 2099 13923
rect 4338 13920 4344 13932
rect 4299 13892 4344 13920
rect 2041 13883 2099 13889
rect 2056 13852 2084 13883
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 6656 13929 6684 13960
rect 6914 13929 6920 13932
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13920 5687 13923
rect 6641 13923 6699 13929
rect 5675 13892 6592 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 2130 13852 2136 13864
rect 2056 13824 2136 13852
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5534 13852 5540 13864
rect 4663 13824 5540 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5718 13852 5724 13864
rect 5679 13824 5724 13852
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 5902 13852 5908 13864
rect 5863 13824 5908 13852
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 6564 13852 6592 13892
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6908 13883 6920 13929
rect 6972 13920 6978 13932
rect 8110 13920 8116 13932
rect 6972 13892 7008 13920
rect 8071 13892 8116 13920
rect 6914 13880 6920 13883
rect 6972 13880 6978 13892
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8386 13929 8392 13932
rect 8380 13920 8392 13929
rect 8347 13892 8392 13920
rect 8380 13883 8392 13892
rect 8386 13880 8392 13883
rect 8444 13880 8450 13932
rect 9692 13920 9720 14016
rect 9766 13948 9772 14000
rect 9824 13988 9830 14000
rect 10106 13991 10164 13997
rect 10106 13988 10118 13991
rect 9824 13960 10118 13988
rect 9824 13948 9830 13960
rect 10106 13957 10118 13960
rect 10152 13988 10164 13991
rect 10870 13988 10876 14000
rect 10152 13960 10876 13988
rect 10152 13957 10164 13960
rect 10106 13951 10164 13957
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9692 13892 9873 13920
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 11532 13920 11560 14019
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 14642 14056 14648 14068
rect 14603 14028 14648 14056
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 14829 14059 14887 14065
rect 14829 14025 14841 14059
rect 14875 14056 14887 14059
rect 15378 14056 15384 14068
rect 14875 14028 15384 14056
rect 14875 14025 14887 14028
rect 14829 14019 14887 14025
rect 15378 14016 15384 14028
rect 15436 14056 15442 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15436 14028 15945 14056
rect 15436 14016 15442 14028
rect 15933 14025 15945 14028
rect 15979 14056 15991 14059
rect 16025 14059 16083 14065
rect 16025 14056 16037 14059
rect 15979 14028 16037 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 16025 14025 16037 14028
rect 16071 14056 16083 14059
rect 16206 14056 16212 14068
rect 16071 14028 16212 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16206 14016 16212 14028
rect 16264 14056 16270 14068
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 16264 14028 16405 14056
rect 16264 14016 16270 14028
rect 16393 14025 16405 14028
rect 16439 14025 16451 14059
rect 17034 14056 17040 14068
rect 16995 14028 17040 14056
rect 16393 14019 16451 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 19610 14056 19616 14068
rect 18064 14028 18828 14056
rect 19571 14028 19616 14056
rect 11882 13948 11888 14000
rect 11940 13988 11946 14000
rect 12038 13991 12096 13997
rect 12038 13988 12050 13991
rect 11940 13960 12050 13988
rect 11940 13948 11946 13960
rect 12038 13957 12050 13960
rect 12084 13957 12096 13991
rect 14274 13988 14280 14000
rect 12038 13951 12096 13957
rect 13280 13960 14280 13988
rect 13280 13929 13308 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 15010 13988 15016 14000
rect 14971 13960 15016 13988
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 15565 13991 15623 13997
rect 15565 13957 15577 13991
rect 15611 13988 15623 13991
rect 18064 13988 18092 14028
rect 15611 13960 18092 13988
rect 15611 13957 15623 13960
rect 15565 13951 15623 13957
rect 18138 13948 18144 14000
rect 18196 13948 18202 14000
rect 18800 13988 18828 14028
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 20898 14016 20904 14068
rect 20956 14056 20962 14068
rect 21085 14059 21143 14065
rect 21085 14056 21097 14059
rect 20956 14028 21097 14056
rect 20956 14016 20962 14028
rect 21085 14025 21097 14028
rect 21131 14056 21143 14059
rect 22189 14059 22247 14065
rect 22189 14056 22201 14059
rect 21131 14028 22201 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 22189 14025 22201 14028
rect 22235 14025 22247 14059
rect 22830 14056 22836 14068
rect 22791 14028 22836 14056
rect 22189 14019 22247 14025
rect 22830 14016 22836 14028
rect 22888 14016 22894 14068
rect 19794 13988 19800 14000
rect 18800 13960 19800 13988
rect 19794 13948 19800 13960
rect 19852 13948 19858 14000
rect 21266 13948 21272 14000
rect 21324 13988 21330 14000
rect 21361 13991 21419 13997
rect 21361 13988 21373 13991
rect 21324 13960 21373 13988
rect 21324 13948 21330 13960
rect 21361 13957 21373 13960
rect 21407 13988 21419 13991
rect 21910 13988 21916 14000
rect 21407 13960 21916 13988
rect 21407 13957 21419 13960
rect 21361 13951 21419 13957
rect 21910 13948 21916 13960
rect 21968 13948 21974 14000
rect 22002 13948 22008 14000
rect 22060 13988 22066 14000
rect 22060 13960 23152 13988
rect 22060 13948 22066 13960
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11532 13892 11805 13920
rect 9861 13883 9919 13889
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 13532 13923 13590 13929
rect 13532 13889 13544 13923
rect 13578 13920 13590 13923
rect 15194 13920 15200 13932
rect 13578 13892 15200 13920
rect 13578 13889 13590 13892
rect 13532 13883 13590 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15749 13923 15807 13929
rect 15749 13889 15761 13923
rect 15795 13920 15807 13923
rect 16114 13920 16120 13932
rect 15795 13892 16120 13920
rect 15795 13889 15807 13892
rect 15749 13883 15807 13889
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 18156 13920 18184 13948
rect 18506 13929 18512 13932
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 16347 13892 18092 13920
rect 18156 13892 18245 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 6564 13824 6684 13852
rect 4154 13716 4160 13728
rect 4115 13688 4160 13716
rect 4154 13676 4160 13688
rect 4212 13676 4218 13728
rect 5166 13716 5172 13728
rect 5127 13688 5172 13716
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 6656 13716 6684 13824
rect 14918 13812 14924 13864
rect 14976 13852 14982 13864
rect 16482 13852 16488 13864
rect 14976 13824 16488 13852
rect 14976 13812 14982 13824
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 16850 13852 16856 13864
rect 16684 13824 16856 13852
rect 15197 13787 15255 13793
rect 15197 13753 15209 13787
rect 15243 13784 15255 13787
rect 15286 13784 15292 13796
rect 15243 13756 15292 13784
rect 15243 13753 15255 13756
rect 15197 13747 15255 13753
rect 15286 13744 15292 13756
rect 15344 13784 15350 13796
rect 16022 13784 16028 13796
rect 15344 13756 16028 13784
rect 15344 13744 15350 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 16684 13793 16712 13824
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 16942 13812 16948 13864
rect 17000 13852 17006 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 17000 13824 17141 13852
rect 17000 13812 17006 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 17310 13852 17316 13864
rect 17271 13824 17316 13852
rect 17129 13815 17187 13821
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 18064 13852 18092 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18500 13920 18512 13929
rect 18467 13892 18512 13920
rect 18233 13883 18291 13889
rect 18500 13883 18512 13892
rect 18138 13852 18144 13864
rect 17696 13824 18000 13852
rect 18064 13824 18144 13852
rect 17696 13793 17724 13824
rect 17972 13793 18000 13824
rect 18138 13812 18144 13824
rect 18196 13812 18202 13864
rect 16669 13787 16727 13793
rect 16669 13753 16681 13787
rect 16715 13753 16727 13787
rect 16669 13747 16727 13753
rect 17589 13787 17647 13793
rect 17589 13753 17601 13787
rect 17635 13784 17647 13787
rect 17681 13787 17739 13793
rect 17681 13784 17693 13787
rect 17635 13756 17693 13784
rect 17635 13753 17647 13756
rect 17589 13747 17647 13753
rect 17681 13753 17693 13756
rect 17727 13753 17739 13787
rect 17681 13747 17739 13753
rect 17957 13787 18015 13793
rect 17957 13753 17969 13787
rect 18003 13784 18015 13787
rect 18049 13787 18107 13793
rect 18049 13784 18061 13787
rect 18003 13756 18061 13784
rect 18003 13753 18015 13756
rect 17957 13747 18015 13753
rect 18049 13753 18061 13756
rect 18095 13784 18107 13787
rect 18248 13784 18276 13883
rect 18506 13880 18512 13883
rect 18564 13880 18570 13932
rect 19978 13929 19984 13932
rect 19972 13920 19984 13929
rect 19891 13892 19984 13920
rect 19972 13883 19984 13892
rect 20036 13920 20042 13932
rect 20036 13892 20760 13920
rect 19978 13880 19984 13883
rect 20036 13880 20042 13892
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13821 19763 13855
rect 20732 13852 20760 13892
rect 21450 13880 21456 13932
rect 21508 13920 21514 13932
rect 23124 13929 23152 13960
rect 22649 13923 22707 13929
rect 21508 13892 22508 13920
rect 21508 13880 21514 13892
rect 21910 13852 21916 13864
rect 20732 13824 21772 13852
rect 21871 13824 21916 13852
rect 19705 13815 19763 13821
rect 18095 13756 18276 13784
rect 18095 13753 18107 13756
rect 18049 13747 18107 13753
rect 7006 13716 7012 13728
rect 5316 13688 5361 13716
rect 6656 13688 7012 13716
rect 5316 13676 5322 13688
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 8018 13716 8024 13728
rect 7979 13688 8024 13716
rect 8018 13676 8024 13688
rect 8076 13676 8082 13728
rect 9214 13676 9220 13728
rect 9272 13716 9278 13728
rect 9493 13719 9551 13725
rect 9493 13716 9505 13719
rect 9272 13688 9505 13716
rect 9272 13676 9278 13688
rect 9493 13685 9505 13688
rect 9539 13685 9551 13719
rect 18248 13716 18276 13756
rect 18598 13716 18604 13728
rect 18248 13688 18604 13716
rect 9493 13679 9551 13685
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 19720 13716 19748 13815
rect 21542 13784 21548 13796
rect 21503 13756 21548 13784
rect 21542 13744 21548 13756
rect 21600 13744 21606 13796
rect 21744 13784 21772 13824
rect 21910 13812 21916 13824
rect 21968 13812 21974 13864
rect 22097 13855 22155 13861
rect 22097 13852 22109 13855
rect 22020 13824 22109 13852
rect 22020 13784 22048 13824
rect 22097 13821 22109 13824
rect 22143 13821 22155 13855
rect 22480 13852 22508 13892
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 23109 13923 23167 13929
rect 22695 13892 23060 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 23032 13852 23060 13892
rect 23109 13889 23121 13923
rect 23155 13889 23167 13923
rect 23109 13883 23167 13889
rect 23842 13852 23848 13864
rect 22480 13824 22968 13852
rect 23032 13824 23848 13852
rect 22097 13815 22155 13821
rect 22940 13793 22968 13824
rect 23842 13812 23848 13824
rect 23900 13812 23906 13864
rect 21744 13756 22048 13784
rect 22925 13787 22983 13793
rect 22925 13753 22937 13787
rect 22971 13753 22983 13787
rect 22925 13747 22983 13753
rect 20070 13716 20076 13728
rect 19720 13688 20076 13716
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 21269 13719 21327 13725
rect 21269 13685 21281 13719
rect 21315 13716 21327 13719
rect 22002 13716 22008 13728
rect 21315 13688 22008 13716
rect 21315 13685 21327 13688
rect 21269 13679 21327 13685
rect 22002 13676 22008 13688
rect 22060 13676 22066 13728
rect 22554 13716 22560 13728
rect 22515 13688 22560 13716
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 1104 13626 23460 13648
rect 1104 13574 3749 13626
rect 3801 13574 3813 13626
rect 3865 13574 3877 13626
rect 3929 13574 3941 13626
rect 3993 13574 4005 13626
rect 4057 13574 9347 13626
rect 9399 13574 9411 13626
rect 9463 13574 9475 13626
rect 9527 13574 9539 13626
rect 9591 13574 9603 13626
rect 9655 13574 14945 13626
rect 14997 13574 15009 13626
rect 15061 13574 15073 13626
rect 15125 13574 15137 13626
rect 15189 13574 15201 13626
rect 15253 13574 20543 13626
rect 20595 13574 20607 13626
rect 20659 13574 20671 13626
rect 20723 13574 20735 13626
rect 20787 13574 20799 13626
rect 20851 13574 23460 13626
rect 1104 13552 23460 13574
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3476 13484 3801 13512
rect 3476 13472 3482 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4396 13484 4629 13512
rect 4396 13472 4402 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 4617 13475 4675 13481
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 6914 13512 6920 13524
rect 6595 13484 6920 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 6564 13444 6592 13475
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8110 13512 8116 13524
rect 8071 13484 8116 13512
rect 8110 13472 8116 13484
rect 8168 13512 8174 13524
rect 8294 13512 8300 13524
rect 8168 13484 8300 13512
rect 8168 13472 8174 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 14185 13515 14243 13521
rect 10928 13484 10973 13512
rect 10928 13472 10934 13484
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 14274 13512 14280 13524
rect 14231 13484 14280 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 14274 13472 14280 13484
rect 14332 13512 14338 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 14332 13484 15301 13512
rect 14332 13472 14338 13484
rect 15289 13481 15301 13484
rect 15335 13512 15347 13515
rect 15378 13512 15384 13524
rect 15335 13484 15384 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 17218 13512 17224 13524
rect 17179 13484 17224 13512
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 18414 13472 18420 13524
rect 18472 13512 18478 13524
rect 21545 13515 21603 13521
rect 18472 13484 20668 13512
rect 18472 13472 18478 13484
rect 6196 13416 6592 13444
rect 4338 13376 4344 13388
rect 4251 13348 4344 13376
rect 4338 13336 4344 13348
rect 4396 13376 4402 13388
rect 4982 13376 4988 13388
rect 4396 13348 4988 13376
rect 4396 13336 4402 13348
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5169 13379 5227 13385
rect 5169 13345 5181 13379
rect 5215 13376 5227 13379
rect 5350 13376 5356 13388
rect 5215 13348 5356 13376
rect 5215 13345 5227 13348
rect 5169 13339 5227 13345
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 6196 13385 6224 13416
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 6270 13336 6276 13388
rect 6328 13376 6334 13388
rect 7929 13379 7987 13385
rect 6328 13348 6373 13376
rect 6328 13336 6334 13348
rect 7929 13345 7941 13379
rect 7975 13376 7987 13379
rect 8128 13376 8156 13472
rect 15102 13444 15108 13456
rect 15063 13416 15108 13444
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 7975 13348 8156 13376
rect 15396 13376 15424 13472
rect 20640 13444 20668 13484
rect 21545 13481 21557 13515
rect 21591 13512 21603 13515
rect 21634 13512 21640 13524
rect 21591 13484 21640 13512
rect 21591 13481 21603 13484
rect 21545 13475 21603 13481
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 22373 13447 22431 13453
rect 22373 13444 22385 13447
rect 20640 13416 22385 13444
rect 22373 13413 22385 13416
rect 22419 13413 22431 13447
rect 22373 13407 22431 13413
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15396 13348 15761 13376
rect 7975 13345 7987 13348
rect 7929 13339 7987 13345
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 18598 13376 18604 13388
rect 18559 13348 18604 13376
rect 15749 13339 15807 13345
rect 18598 13336 18604 13348
rect 18656 13336 18662 13388
rect 20901 13379 20959 13385
rect 20901 13345 20913 13379
rect 20947 13376 20959 13379
rect 21450 13376 21456 13388
rect 20947 13348 21456 13376
rect 20947 13345 20959 13348
rect 20901 13339 20959 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 21818 13336 21824 13388
rect 21876 13376 21882 13388
rect 22005 13379 22063 13385
rect 22005 13376 22017 13379
rect 21876 13348 22017 13376
rect 21876 13336 21882 13348
rect 22005 13345 22017 13348
rect 22051 13345 22063 13379
rect 22005 13339 22063 13345
rect 22097 13379 22155 13385
rect 22097 13345 22109 13379
rect 22143 13345 22155 13379
rect 22097 13339 22155 13345
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 4430 13308 4436 13320
rect 3467 13280 4436 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 5258 13308 5264 13320
rect 5123 13280 5264 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 8018 13308 8024 13320
rect 6135 13280 8024 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 8018 13268 8024 13280
rect 8076 13308 8082 13320
rect 10514 13311 10572 13317
rect 10514 13308 10526 13311
rect 8076 13280 10526 13308
rect 8076 13268 8082 13280
rect 10514 13277 10526 13280
rect 10560 13277 10572 13311
rect 10514 13271 10572 13277
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13308 10839 13311
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 10827 13280 12265 13308
rect 10827 13277 10839 13280
rect 10781 13271 10839 13277
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 13170 13308 13176 13320
rect 13131 13280 13176 13308
rect 12253 13271 12311 13277
rect 4157 13243 4215 13249
rect 4157 13240 4169 13243
rect 3620 13212 4169 13240
rect 3620 13181 3648 13212
rect 4157 13209 4169 13212
rect 4203 13209 4215 13243
rect 4157 13203 4215 13209
rect 4985 13243 5043 13249
rect 4985 13209 4997 13243
rect 5031 13240 5043 13243
rect 5031 13212 5764 13240
rect 5031 13209 5043 13212
rect 4985 13203 5043 13209
rect 3605 13175 3663 13181
rect 3605 13141 3617 13175
rect 3651 13141 3663 13175
rect 3605 13135 3663 13141
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 5736 13181 5764 13212
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 7684 13243 7742 13249
rect 7684 13240 7696 13243
rect 7064 13212 7696 13240
rect 7064 13200 7070 13212
rect 7684 13209 7696 13212
rect 7730 13240 7742 13243
rect 8202 13240 8208 13252
rect 7730 13212 8208 13240
rect 7730 13209 7742 13212
rect 7684 13203 7742 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 8294 13200 8300 13252
rect 8352 13240 8358 13252
rect 8389 13243 8447 13249
rect 8389 13240 8401 13243
rect 8352 13212 8401 13240
rect 8352 13200 8358 13212
rect 8389 13209 8401 13212
rect 8435 13240 8447 13243
rect 9030 13240 9036 13252
rect 8435 13212 9036 13240
rect 8435 13209 8447 13212
rect 8389 13203 8447 13209
rect 9030 13200 9036 13212
rect 9088 13200 9094 13252
rect 10962 13240 10968 13252
rect 10520 13212 10968 13240
rect 10520 13184 10548 13212
rect 10962 13200 10968 13212
rect 11020 13240 11026 13252
rect 11986 13243 12044 13249
rect 11986 13240 11998 13243
rect 11020 13212 11998 13240
rect 11020 13200 11026 13212
rect 11986 13209 11998 13212
rect 12032 13209 12044 13243
rect 11986 13203 12044 13209
rect 5721 13175 5779 13181
rect 4304 13144 4349 13172
rect 4304 13132 4310 13144
rect 5721 13141 5733 13175
rect 5767 13141 5779 13175
rect 5721 13135 5779 13141
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 9214 13172 9220 13184
rect 5868 13144 9220 13172
rect 5868 13132 5874 13144
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9398 13172 9404 13184
rect 9359 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 10502 13132 10508 13184
rect 10560 13132 10566 13184
rect 12268 13172 12296 13271
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 15703 13280 18889 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 18877 13277 18889 13280
rect 18923 13308 18935 13311
rect 19334 13308 19340 13320
rect 18923 13280 19340 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 20070 13268 20076 13320
rect 20128 13308 20134 13320
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 20128 13280 20637 13308
rect 20128 13268 20134 13280
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 22112 13308 22140 13339
rect 22554 13336 22560 13388
rect 22612 13376 22618 13388
rect 22833 13379 22891 13385
rect 22833 13376 22845 13379
rect 22612 13348 22845 13376
rect 22612 13336 22618 13348
rect 22833 13345 22845 13348
rect 22879 13345 22891 13379
rect 22833 13339 22891 13345
rect 22922 13336 22928 13388
rect 22980 13376 22986 13388
rect 22980 13348 23025 13376
rect 22980 13336 22986 13348
rect 22186 13308 22192 13320
rect 22112 13280 22192 13308
rect 20625 13271 20683 13277
rect 22186 13268 22192 13280
rect 22244 13308 22250 13320
rect 22940 13308 22968 13336
rect 22244 13280 22968 13308
rect 22244 13268 22250 13280
rect 16022 13249 16028 13252
rect 16016 13203 16028 13249
rect 16080 13240 16086 13252
rect 18334 13243 18392 13249
rect 18334 13240 18346 13243
rect 16080 13212 16116 13240
rect 17144 13212 18346 13240
rect 16022 13200 16028 13203
rect 16080 13200 16086 13212
rect 12437 13175 12495 13181
rect 12437 13172 12449 13175
rect 12268 13144 12449 13172
rect 12437 13141 12449 13144
rect 12483 13172 12495 13175
rect 12802 13172 12808 13184
rect 12483 13144 12808 13172
rect 12483 13141 12495 13144
rect 12437 13135 12495 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13814 13172 13820 13184
rect 13775 13144 13820 13172
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 17034 13132 17040 13184
rect 17092 13172 17098 13184
rect 17144 13181 17172 13212
rect 18334 13209 18346 13212
rect 18380 13209 18392 13243
rect 18334 13203 18392 13209
rect 18785 13243 18843 13249
rect 18785 13209 18797 13243
rect 18831 13240 18843 13243
rect 19150 13240 19156 13252
rect 18831 13212 19156 13240
rect 18831 13209 18843 13212
rect 18785 13203 18843 13209
rect 19150 13200 19156 13212
rect 19208 13240 19214 13252
rect 19426 13240 19432 13252
rect 19208 13212 19432 13240
rect 19208 13200 19214 13212
rect 19426 13200 19432 13212
rect 19484 13200 19490 13252
rect 20380 13243 20438 13249
rect 20380 13209 20392 13243
rect 20426 13240 20438 13243
rect 20898 13240 20904 13252
rect 20426 13212 20904 13240
rect 20426 13209 20438 13212
rect 20380 13203 20438 13209
rect 20898 13200 20904 13212
rect 20956 13200 20962 13252
rect 21082 13240 21088 13252
rect 21043 13212 21088 13240
rect 21082 13200 21088 13212
rect 21140 13200 21146 13252
rect 21913 13243 21971 13249
rect 21913 13240 21925 13243
rect 21468 13212 21925 13240
rect 17129 13175 17187 13181
rect 17129 13172 17141 13175
rect 17092 13144 17141 13172
rect 17092 13132 17098 13144
rect 17129 13141 17141 13144
rect 17175 13141 17187 13175
rect 19058 13172 19064 13184
rect 19019 13144 19064 13172
rect 17129 13135 17187 13141
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 19245 13175 19303 13181
rect 19245 13141 19257 13175
rect 19291 13172 19303 13175
rect 19610 13172 19616 13184
rect 19291 13144 19616 13172
rect 19291 13141 19303 13144
rect 19245 13135 19303 13141
rect 19610 13132 19616 13144
rect 19668 13132 19674 13184
rect 19702 13132 19708 13184
rect 19760 13172 19766 13184
rect 21468 13181 21496 13212
rect 21913 13209 21925 13212
rect 21959 13209 21971 13243
rect 21913 13203 21971 13209
rect 20993 13175 21051 13181
rect 20993 13172 21005 13175
rect 19760 13144 21005 13172
rect 19760 13132 19766 13144
rect 20993 13141 21005 13144
rect 21039 13141 21051 13175
rect 20993 13135 21051 13141
rect 21453 13175 21511 13181
rect 21453 13141 21465 13175
rect 21499 13141 21511 13175
rect 21453 13135 21511 13141
rect 21542 13132 21548 13184
rect 21600 13172 21606 13184
rect 22741 13175 22799 13181
rect 22741 13172 22753 13175
rect 21600 13144 22753 13172
rect 21600 13132 21606 13144
rect 22741 13141 22753 13144
rect 22787 13141 22799 13175
rect 22741 13135 22799 13141
rect 1104 13082 23460 13104
rect 1104 13030 6548 13082
rect 6600 13030 6612 13082
rect 6664 13030 6676 13082
rect 6728 13030 6740 13082
rect 6792 13030 6804 13082
rect 6856 13030 12146 13082
rect 12198 13030 12210 13082
rect 12262 13030 12274 13082
rect 12326 13030 12338 13082
rect 12390 13030 12402 13082
rect 12454 13030 17744 13082
rect 17796 13030 17808 13082
rect 17860 13030 17872 13082
rect 17924 13030 17936 13082
rect 17988 13030 18000 13082
rect 18052 13030 23460 13082
rect 1104 13008 23460 13030
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 3605 12971 3663 12977
rect 3605 12968 3617 12971
rect 3292 12940 3617 12968
rect 3292 12928 3298 12940
rect 3605 12937 3617 12940
rect 3651 12937 3663 12971
rect 3605 12931 3663 12937
rect 4065 12971 4123 12977
rect 4065 12937 4077 12971
rect 4111 12968 4123 12971
rect 4154 12968 4160 12980
rect 4111 12940 4160 12968
rect 4111 12937 4123 12940
rect 4065 12931 4123 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4430 12968 4436 12980
rect 4391 12940 4436 12968
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 4801 12971 4859 12977
rect 4801 12937 4813 12971
rect 4847 12968 4859 12971
rect 5166 12968 5172 12980
rect 4847 12940 5172 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5810 12968 5816 12980
rect 5771 12940 5816 12968
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 6825 12971 6883 12977
rect 6825 12937 6837 12971
rect 6871 12968 6883 12971
rect 9398 12968 9404 12980
rect 6871 12940 9404 12968
rect 6871 12937 6883 12940
rect 6825 12931 6883 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10597 12971 10655 12977
rect 10597 12937 10609 12971
rect 10643 12968 10655 12971
rect 11054 12968 11060 12980
rect 10643 12940 11060 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 11606 12968 11612 12980
rect 11388 12940 11612 12968
rect 11388 12928 11394 12940
rect 11606 12928 11612 12940
rect 11664 12968 11670 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 11664 12940 12633 12968
rect 11664 12928 11670 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 12621 12931 12679 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 16206 12968 16212 12980
rect 13127 12940 14780 12968
rect 16167 12940 16212 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 4890 12900 4896 12912
rect 4851 12872 4896 12900
rect 4890 12860 4896 12872
rect 4948 12860 4954 12912
rect 7285 12903 7343 12909
rect 7285 12869 7297 12903
rect 7331 12900 7343 12903
rect 9030 12900 9036 12912
rect 7331 12872 9036 12900
rect 7331 12869 7343 12872
rect 7285 12863 7343 12869
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 8772 12841 8800 12872
rect 9030 12860 9036 12872
rect 9088 12900 9094 12912
rect 9088 12872 11284 12900
rect 9088 12860 9094 12872
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3384 12804 3985 12832
rect 3384 12792 3390 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12832 6791 12835
rect 8490 12835 8548 12841
rect 8490 12832 8502 12835
rect 6779 12804 8502 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 8490 12801 8502 12804
rect 8536 12832 8548 12835
rect 8757 12835 8815 12841
rect 8536 12804 8708 12832
rect 8536 12801 8548 12804
rect 8490 12795 8548 12801
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12764 4307 12767
rect 4338 12764 4344 12776
rect 4295 12736 4344 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 5077 12767 5135 12773
rect 5077 12764 5089 12767
rect 5040 12736 5089 12764
rect 5040 12724 5046 12736
rect 5077 12733 5089 12736
rect 5123 12764 5135 12767
rect 5350 12764 5356 12776
rect 5123 12736 5356 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 5920 12696 5948 12727
rect 6086 12724 6092 12776
rect 6144 12764 6150 12776
rect 6362 12764 6368 12776
rect 6144 12736 6368 12764
rect 6144 12724 6150 12736
rect 6362 12724 6368 12736
rect 6420 12764 6426 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6420 12736 6929 12764
rect 6420 12724 6426 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 8680 12764 8708 12804
rect 8757 12801 8769 12835
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 10244 12841 10272 12872
rect 9962 12835 10020 12841
rect 9962 12832 9974 12835
rect 9456 12804 9974 12832
rect 9456 12792 9462 12804
rect 9962 12801 9974 12804
rect 10008 12801 10020 12835
rect 9962 12795 10020 12801
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12801 10287 12835
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10229 12795 10287 12801
rect 10428 12804 10701 12832
rect 8680 12736 8892 12764
rect 6917 12727 6975 12733
rect 8864 12705 8892 12736
rect 8849 12699 8907 12705
rect 5920 12668 7880 12696
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 5445 12631 5503 12637
rect 5445 12628 5457 12631
rect 4948 12600 5457 12628
rect 4948 12588 4954 12600
rect 5445 12597 5457 12600
rect 5491 12597 5503 12631
rect 6362 12628 6368 12640
rect 6323 12600 6368 12628
rect 5445 12591 5503 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 7374 12628 7380 12640
rect 7335 12600 7380 12628
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 7852 12628 7880 12668
rect 8849 12665 8861 12699
rect 8895 12665 8907 12699
rect 8849 12659 8907 12665
rect 8386 12628 8392 12640
rect 7852 12600 8392 12628
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 10428 12628 10456 12804
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 10520 12696 10548 12727
rect 10778 12696 10784 12708
rect 10520 12668 10784 12696
rect 10778 12656 10784 12668
rect 10836 12656 10842 12708
rect 11054 12696 11060 12708
rect 11015 12668 11060 12696
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 11256 12705 11284 12872
rect 12802 12860 12808 12912
rect 12860 12900 12866 12912
rect 14752 12900 14780 12940
rect 16206 12928 16212 12940
rect 16264 12968 16270 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 16264 12940 16405 12968
rect 16264 12928 16270 12940
rect 16393 12937 16405 12940
rect 16439 12968 16451 12971
rect 17310 12968 17316 12980
rect 16439 12940 17316 12968
rect 16439 12937 16451 12940
rect 16393 12931 16451 12937
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 18322 12968 18328 12980
rect 18283 12940 18328 12968
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 20165 12971 20223 12977
rect 20165 12968 20177 12971
rect 19996 12940 20177 12968
rect 16298 12900 16304 12912
rect 12860 12872 14320 12900
rect 14752 12872 16304 12900
rect 12860 12860 12866 12872
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 13188 12841 13216 12872
rect 14292 12844 14320 12872
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 17782 12903 17840 12909
rect 17782 12900 17794 12903
rect 16540 12872 17794 12900
rect 16540 12860 16546 12872
rect 17782 12869 17794 12872
rect 17828 12869 17840 12903
rect 18960 12903 19018 12909
rect 17782 12863 17840 12869
rect 18156 12872 18920 12900
rect 18156 12844 18184 12872
rect 12713 12835 12771 12841
rect 12713 12832 12725 12835
rect 11848 12804 12725 12832
rect 11848 12792 11854 12804
rect 12713 12801 12725 12804
rect 12759 12801 12771 12835
rect 12713 12795 12771 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 13440 12835 13498 12841
rect 13440 12801 13452 12835
rect 13486 12832 13498 12835
rect 13814 12832 13820 12844
rect 13486 12804 13820 12832
rect 13486 12801 13498 12804
rect 13440 12795 13498 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 14332 12804 14657 12832
rect 14332 12792 14338 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14912 12835 14970 12841
rect 14912 12801 14924 12835
rect 14958 12832 14970 12835
rect 15378 12832 15384 12844
rect 14958 12804 15384 12832
rect 14958 12801 14970 12804
rect 14912 12795 14970 12801
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 18138 12832 18144 12844
rect 18099 12804 18144 12832
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 18414 12832 18420 12844
rect 18375 12804 18420 12832
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18892 12832 18920 12872
rect 18960 12869 18972 12903
rect 19006 12900 19018 12903
rect 19996 12900 20024 12940
rect 20165 12937 20177 12940
rect 20211 12968 20223 12971
rect 22189 12971 22247 12977
rect 22189 12968 22201 12971
rect 20211 12940 22201 12968
rect 20211 12937 20223 12940
rect 20165 12931 20223 12937
rect 22189 12937 22201 12940
rect 22235 12937 22247 12971
rect 22189 12931 22247 12937
rect 22370 12928 22376 12980
rect 22428 12968 22434 12980
rect 22649 12971 22707 12977
rect 22649 12968 22661 12971
rect 22428 12940 22661 12968
rect 22428 12928 22434 12940
rect 22649 12937 22661 12940
rect 22695 12937 22707 12971
rect 22649 12931 22707 12937
rect 19006 12872 20024 12900
rect 19006 12869 19018 12872
rect 18960 12863 19018 12869
rect 19334 12832 19340 12844
rect 18892 12804 19340 12832
rect 19334 12792 19340 12804
rect 19392 12792 19398 12844
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 21278 12835 21336 12841
rect 21278 12832 21290 12835
rect 20404 12804 21290 12832
rect 20404 12792 20410 12804
rect 21278 12801 21290 12804
rect 21324 12832 21336 12835
rect 21545 12835 21603 12841
rect 21324 12804 21496 12832
rect 21324 12801 21336 12804
rect 21278 12795 21336 12801
rect 12529 12767 12587 12773
rect 12529 12733 12541 12767
rect 12575 12733 12587 12767
rect 12529 12727 12587 12733
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18598 12764 18604 12776
rect 18095 12736 18604 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 11241 12699 11299 12705
rect 11241 12665 11253 12699
rect 11287 12696 11299 12699
rect 12544 12696 12572 12727
rect 18598 12724 18604 12736
rect 18656 12764 18662 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18656 12736 18705 12764
rect 18656 12724 18662 12736
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 21468 12764 21496 12804
rect 21545 12801 21557 12835
rect 21591 12832 21603 12835
rect 21634 12832 21640 12844
rect 21591 12804 21640 12832
rect 21591 12801 21603 12804
rect 21545 12795 21603 12801
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 22002 12792 22008 12844
rect 22060 12832 22066 12844
rect 23106 12832 23112 12844
rect 22060 12804 22416 12832
rect 23067 12804 23112 12832
rect 22060 12792 22066 12804
rect 22388 12773 22416 12804
rect 23106 12792 23112 12804
rect 23164 12792 23170 12844
rect 22281 12767 22339 12773
rect 22281 12764 22293 12767
rect 21468 12736 22293 12764
rect 18693 12727 18751 12733
rect 22281 12733 22293 12736
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12733 22431 12767
rect 22373 12727 22431 12733
rect 12710 12696 12716 12708
rect 11287 12668 11652 12696
rect 12544 12668 12716 12696
rect 11287 12665 11299 12668
rect 11241 12659 11299 12665
rect 11422 12628 11428 12640
rect 10428 12600 11428 12628
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 11624 12637 11652 12668
rect 12710 12656 12716 12668
rect 12768 12656 12774 12708
rect 16022 12696 16028 12708
rect 15983 12668 16028 12696
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 19978 12656 19984 12708
rect 20036 12696 20042 12708
rect 20073 12699 20131 12705
rect 20073 12696 20085 12699
rect 20036 12668 20085 12696
rect 20036 12656 20042 12668
rect 20073 12665 20085 12668
rect 20119 12665 20131 12699
rect 20073 12659 20131 12665
rect 11609 12631 11667 12637
rect 11609 12597 11621 12631
rect 11655 12628 11667 12631
rect 12158 12628 12164 12640
rect 11655 12600 12164 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 14553 12631 14611 12637
rect 14553 12597 14565 12631
rect 14599 12628 14611 12631
rect 15378 12628 15384 12640
rect 14599 12600 15384 12628
rect 14599 12597 14611 12600
rect 14553 12591 14611 12597
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 16666 12628 16672 12640
rect 16627 12600 16672 12628
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 18414 12628 18420 12640
rect 17184 12600 18420 12628
rect 17184 12588 17190 12600
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18601 12631 18659 12637
rect 18601 12597 18613 12631
rect 18647 12628 18659 12631
rect 19058 12628 19064 12640
rect 18647 12600 19064 12628
rect 18647 12597 18659 12600
rect 18601 12591 18659 12597
rect 19058 12588 19064 12600
rect 19116 12588 19122 12640
rect 21821 12631 21879 12637
rect 21821 12597 21833 12631
rect 21867 12628 21879 12631
rect 22002 12628 22008 12640
rect 21867 12600 22008 12628
rect 21867 12597 21879 12600
rect 21821 12591 21879 12597
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 22922 12628 22928 12640
rect 22883 12600 22928 12628
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 1104 12538 23460 12560
rect 1104 12486 3749 12538
rect 3801 12486 3813 12538
rect 3865 12486 3877 12538
rect 3929 12486 3941 12538
rect 3993 12486 4005 12538
rect 4057 12486 9347 12538
rect 9399 12486 9411 12538
rect 9463 12486 9475 12538
rect 9527 12486 9539 12538
rect 9591 12486 9603 12538
rect 9655 12486 14945 12538
rect 14997 12486 15009 12538
rect 15061 12486 15073 12538
rect 15125 12486 15137 12538
rect 15189 12486 15201 12538
rect 15253 12486 20543 12538
rect 20595 12486 20607 12538
rect 20659 12486 20671 12538
rect 20723 12486 20735 12538
rect 20787 12486 20799 12538
rect 20851 12486 23460 12538
rect 1104 12464 23460 12486
rect 6362 12424 6368 12436
rect 4448 12396 6368 12424
rect 4448 12297 4476 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8481 12427 8539 12433
rect 8481 12424 8493 12427
rect 8444 12396 8493 12424
rect 8444 12384 8450 12396
rect 8481 12393 8493 12396
rect 8527 12393 8539 12427
rect 8481 12387 8539 12393
rect 9140 12396 10456 12424
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12288 4675 12291
rect 5074 12288 5080 12300
rect 4663 12260 5080 12288
rect 4663 12257 4675 12260
rect 4617 12251 4675 12257
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 5994 12288 6000 12300
rect 5491 12260 6000 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 9140 12297 9168 12396
rect 9677 12359 9735 12365
rect 9677 12325 9689 12359
rect 9723 12325 9735 12359
rect 10428 12356 10456 12396
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 10560 12396 10609 12424
rect 10560 12384 10566 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 11606 12424 11612 12436
rect 10597 12387 10655 12393
rect 10796 12396 11612 12424
rect 10796 12368 10824 12396
rect 11606 12384 11612 12396
rect 11664 12424 11670 12436
rect 12158 12424 12164 12436
rect 11664 12396 12020 12424
rect 12071 12396 12164 12424
rect 11664 12384 11670 12396
rect 10778 12356 10784 12368
rect 10428 12328 10784 12356
rect 9677 12319 9735 12325
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12257 9183 12291
rect 9125 12251 9183 12257
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12220 5227 12223
rect 7009 12223 7067 12229
rect 5215 12192 6868 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12152 4399 12155
rect 5442 12152 5448 12164
rect 4387 12124 5448 12152
rect 4387 12121 4399 12124
rect 4341 12115 4399 12121
rect 5442 12112 5448 12124
rect 5500 12112 5506 12164
rect 6454 12112 6460 12164
rect 6512 12152 6518 12164
rect 6742 12155 6800 12161
rect 6742 12152 6754 12155
rect 6512 12124 6754 12152
rect 6512 12112 6518 12124
rect 6742 12121 6754 12124
rect 6788 12121 6800 12155
rect 6840 12152 6868 12192
rect 7009 12189 7021 12223
rect 7055 12220 7067 12223
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 7055 12192 7113 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 7101 12189 7113 12192
rect 7147 12220 7159 12223
rect 7147 12192 8064 12220
rect 7147 12189 7159 12192
rect 7101 12183 7159 12189
rect 8036 12164 8064 12192
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 8996 12192 9321 12220
rect 8996 12180 9002 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9692 12220 9720 12319
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11992 12356 12020 12396
rect 12158 12384 12164 12396
rect 12216 12424 12222 12436
rect 12802 12424 12808 12436
rect 12216 12396 12808 12424
rect 12216 12384 12222 12396
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 13265 12427 13323 12433
rect 13265 12393 13277 12427
rect 13311 12424 13323 12427
rect 13906 12424 13912 12436
rect 13311 12396 13912 12424
rect 13311 12393 13323 12396
rect 13265 12387 13323 12393
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 16574 12424 16580 12436
rect 14016 12396 16160 12424
rect 16535 12396 16580 12424
rect 12250 12356 12256 12368
rect 11992 12328 12256 12356
rect 12250 12316 12256 12328
rect 12308 12316 12314 12368
rect 14016 12356 14044 12396
rect 12406 12328 14044 12356
rect 10318 12288 10324 12300
rect 10279 12260 10324 12288
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 12158 12288 12164 12300
rect 12023 12260 12164 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12406 12220 12434 12328
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 14461 12359 14519 12365
rect 14461 12356 14473 12359
rect 14332 12328 14473 12356
rect 14332 12316 14338 12328
rect 14461 12325 14473 12328
rect 14507 12356 14519 12359
rect 14645 12359 14703 12365
rect 14645 12356 14657 12359
rect 14507 12328 14657 12356
rect 14507 12325 14519 12328
rect 14461 12319 14519 12325
rect 14645 12325 14657 12328
rect 14691 12356 14703 12359
rect 15102 12356 15108 12368
rect 14691 12328 15108 12356
rect 14691 12325 14703 12328
rect 14645 12319 14703 12325
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 12710 12288 12716 12300
rect 12671 12260 12716 12288
rect 12710 12248 12716 12260
rect 12768 12288 12774 12300
rect 13722 12288 13728 12300
rect 12768 12260 13728 12288
rect 12768 12248 12774 12260
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 16132 12288 16160 12396
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 18506 12424 18512 12436
rect 16684 12396 18512 12424
rect 16482 12356 16488 12368
rect 16443 12328 16488 12356
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 16684 12288 16712 12396
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 21450 12424 21456 12436
rect 18892 12396 20208 12424
rect 21411 12396 21456 12424
rect 14568 12260 15240 12288
rect 16132 12260 16712 12288
rect 16776 12328 17632 12356
rect 9692 12192 12434 12220
rect 12897 12223 12955 12229
rect 9309 12183 9367 12189
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 13170 12220 13176 12232
rect 12943 12192 13176 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 7190 12152 7196 12164
rect 6840 12124 7196 12152
rect 6742 12115 6800 12121
rect 7190 12112 7196 12124
rect 7248 12152 7254 12164
rect 7346 12155 7404 12161
rect 7346 12152 7358 12155
rect 7248 12124 7358 12152
rect 7248 12112 7254 12124
rect 7346 12121 7358 12124
rect 7392 12121 7404 12155
rect 7346 12115 7404 12121
rect 8018 12112 8024 12164
rect 8076 12152 8082 12164
rect 8573 12155 8631 12161
rect 8573 12152 8585 12155
rect 8076 12124 8585 12152
rect 8076 12112 8082 12124
rect 8573 12121 8585 12124
rect 8619 12121 8631 12155
rect 8573 12115 8631 12121
rect 9217 12155 9275 12161
rect 9217 12121 9229 12155
rect 9263 12152 9275 12155
rect 10137 12155 10195 12161
rect 9263 12124 9812 12152
rect 9263 12121 9275 12124
rect 9217 12115 9275 12121
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 3973 12087 4031 12093
rect 3973 12084 3985 12087
rect 3200 12056 3985 12084
rect 3200 12044 3206 12056
rect 3973 12053 3985 12056
rect 4019 12053 4031 12087
rect 3973 12047 4031 12053
rect 4801 12087 4859 12093
rect 4801 12053 4813 12087
rect 4847 12084 4859 12087
rect 4982 12084 4988 12096
rect 4847 12056 4988 12084
rect 4847 12053 4859 12056
rect 4801 12047 4859 12053
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 5629 12087 5687 12093
rect 5629 12084 5641 12087
rect 5307 12056 5641 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 5629 12053 5641 12056
rect 5675 12084 5687 12087
rect 7006 12084 7012 12096
rect 5675 12056 7012 12084
rect 5675 12053 5687 12056
rect 5629 12047 5687 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 9784 12093 9812 12124
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10410 12152 10416 12164
rect 10183 12124 10416 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10410 12112 10416 12124
rect 10468 12152 10474 12164
rect 11710 12155 11768 12161
rect 11710 12152 11722 12155
rect 10468 12124 11722 12152
rect 10468 12112 10474 12124
rect 11710 12121 11722 12124
rect 11756 12121 11768 12155
rect 11710 12115 11768 12121
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 14568 12152 14596 12260
rect 15102 12220 15108 12232
rect 15063 12192 15108 12220
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 15212 12220 15240 12260
rect 16776 12220 16804 12328
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 17604 12297 17632 12328
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 16908 12260 17141 12288
rect 16908 12248 16914 12260
rect 17129 12257 17141 12260
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 17954 12288 17960 12300
rect 17635 12260 17960 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 15212 12192 16804 12220
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12220 17003 12223
rect 17218 12220 17224 12232
rect 16991 12192 17224 12220
rect 16991 12189 17003 12192
rect 16945 12183 17003 12189
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 18322 12180 18328 12232
rect 18380 12220 18386 12232
rect 18509 12223 18567 12229
rect 18509 12220 18521 12223
rect 18380 12192 18521 12220
rect 18380 12180 18386 12192
rect 18509 12189 18521 12192
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 18892 12229 18920 12396
rect 20180 12356 20208 12396
rect 21450 12384 21456 12396
rect 21508 12384 21514 12436
rect 21910 12384 21916 12436
rect 21968 12384 21974 12436
rect 21928 12356 21956 12384
rect 20180 12328 21588 12356
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12288 20959 12291
rect 21358 12288 21364 12300
rect 20947 12260 21364 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 21358 12248 21364 12260
rect 21416 12248 21422 12300
rect 18877 12223 18935 12229
rect 18656 12192 18701 12220
rect 18656 12180 18662 12192
rect 18877 12189 18889 12223
rect 18923 12189 18935 12223
rect 18877 12183 18935 12189
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19334 12220 19340 12232
rect 19291 12192 19340 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 12308 12124 14596 12152
rect 15372 12155 15430 12161
rect 12308 12112 12314 12124
rect 15372 12121 15384 12155
rect 15418 12152 15430 12155
rect 15470 12152 15476 12164
rect 15418 12124 15476 12152
rect 15418 12121 15430 12124
rect 15372 12115 15430 12121
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 16482 12112 16488 12164
rect 16540 12152 16546 12164
rect 17773 12155 17831 12161
rect 17773 12152 17785 12155
rect 16540 12124 17785 12152
rect 16540 12112 16546 12124
rect 17773 12121 17785 12124
rect 17819 12121 17831 12155
rect 17773 12115 17831 12121
rect 18690 12112 18696 12164
rect 18748 12152 18754 12164
rect 19260 12152 19288 12183
rect 19334 12180 19340 12192
rect 19392 12220 19398 12232
rect 19978 12220 19984 12232
rect 19392 12192 19984 12220
rect 19392 12180 19398 12192
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20993 12223 21051 12229
rect 20993 12220 21005 12223
rect 20180 12192 21005 12220
rect 18748 12124 19288 12152
rect 19512 12155 19570 12161
rect 18748 12112 18754 12124
rect 19512 12121 19524 12155
rect 19558 12152 19570 12155
rect 19610 12152 19616 12164
rect 19558 12124 19616 12152
rect 19558 12121 19570 12124
rect 19512 12115 19570 12121
rect 19610 12112 19616 12124
rect 19668 12152 19674 12164
rect 20180 12152 20208 12192
rect 20993 12189 21005 12192
rect 21039 12189 21051 12223
rect 20993 12183 21051 12189
rect 21085 12155 21143 12161
rect 21085 12152 21097 12155
rect 19668 12124 20208 12152
rect 20824 12124 21097 12152
rect 19668 12112 19674 12124
rect 9769 12087 9827 12093
rect 9769 12053 9781 12087
rect 9815 12053 9827 12087
rect 9769 12047 9827 12053
rect 10229 12087 10287 12093
rect 10229 12053 10241 12087
rect 10275 12084 10287 12087
rect 11974 12084 11980 12096
rect 10275 12056 11980 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12802 12084 12808 12096
rect 12763 12056 12808 12084
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 15013 12087 15071 12093
rect 15013 12053 15025 12087
rect 15059 12084 15071 12087
rect 16942 12084 16948 12096
rect 15059 12056 16948 12084
rect 15059 12053 15071 12056
rect 15013 12047 15071 12053
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 17034 12044 17040 12096
rect 17092 12084 17098 12096
rect 17092 12056 17137 12084
rect 17092 12044 17098 12056
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 17681 12087 17739 12093
rect 17681 12084 17693 12087
rect 17460 12056 17693 12084
rect 17460 12044 17466 12056
rect 17681 12053 17693 12056
rect 17727 12053 17739 12087
rect 18138 12084 18144 12096
rect 18099 12056 18144 12084
rect 17681 12047 17739 12053
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 18288 12056 18337 12084
rect 18288 12044 18294 12056
rect 18325 12053 18337 12056
rect 18371 12053 18383 12087
rect 18782 12084 18788 12096
rect 18743 12056 18788 12084
rect 18325 12047 18383 12053
rect 18782 12044 18788 12056
rect 18840 12044 18846 12096
rect 19061 12087 19119 12093
rect 19061 12053 19073 12087
rect 19107 12084 19119 12087
rect 19794 12084 19800 12096
rect 19107 12056 19800 12084
rect 19107 12053 19119 12056
rect 19061 12047 19119 12053
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 20254 12044 20260 12096
rect 20312 12084 20318 12096
rect 20625 12087 20683 12093
rect 20625 12084 20637 12087
rect 20312 12056 20637 12084
rect 20312 12044 20318 12056
rect 20625 12053 20637 12056
rect 20671 12084 20683 12087
rect 20824 12084 20852 12124
rect 21085 12121 21097 12124
rect 21131 12121 21143 12155
rect 21085 12115 21143 12121
rect 21560 12093 21588 12328
rect 21836 12328 21956 12356
rect 21726 12180 21732 12232
rect 21784 12220 21790 12232
rect 21836 12220 21864 12328
rect 22646 12316 22652 12368
rect 22704 12356 22710 12368
rect 22922 12356 22928 12368
rect 22704 12328 22928 12356
rect 22704 12316 22710 12328
rect 22922 12316 22928 12328
rect 22980 12316 22986 12368
rect 22186 12248 22192 12300
rect 22244 12288 22250 12300
rect 22370 12288 22376 12300
rect 22244 12260 22376 12288
rect 22244 12248 22250 12260
rect 22370 12248 22376 12260
rect 22428 12248 22434 12300
rect 23014 12288 23020 12300
rect 22975 12260 23020 12288
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 21784 12192 21864 12220
rect 21913 12223 21971 12229
rect 21784 12180 21790 12192
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22002 12220 22008 12232
rect 21959 12192 22008 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22796 12192 22845 12220
rect 22796 12180 22802 12192
rect 22833 12189 22845 12192
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 21634 12112 21640 12164
rect 21692 12152 21698 12164
rect 21692 12124 22416 12152
rect 21692 12112 21698 12124
rect 20671 12056 20852 12084
rect 21545 12087 21603 12093
rect 20671 12053 20683 12056
rect 20625 12047 20683 12053
rect 21545 12053 21557 12087
rect 21591 12053 21603 12087
rect 22002 12084 22008 12096
rect 21963 12056 22008 12084
rect 21545 12047 21603 12053
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 22388 12093 22416 12124
rect 22373 12087 22431 12093
rect 22373 12053 22385 12087
rect 22419 12084 22431 12087
rect 22554 12084 22560 12096
rect 22419 12056 22560 12084
rect 22419 12053 22431 12056
rect 22373 12047 22431 12053
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 22738 12084 22744 12096
rect 22699 12056 22744 12084
rect 22738 12044 22744 12056
rect 22796 12044 22802 12096
rect 1104 11994 23460 12016
rect 1104 11942 6548 11994
rect 6600 11942 6612 11994
rect 6664 11942 6676 11994
rect 6728 11942 6740 11994
rect 6792 11942 6804 11994
rect 6856 11942 12146 11994
rect 12198 11942 12210 11994
rect 12262 11942 12274 11994
rect 12326 11942 12338 11994
rect 12390 11942 12402 11994
rect 12454 11942 17744 11994
rect 17796 11942 17808 11994
rect 17860 11942 17872 11994
rect 17924 11942 17936 11994
rect 17988 11942 18000 11994
rect 18052 11942 23460 11994
rect 1104 11920 23460 11942
rect 3326 11880 3332 11892
rect 3287 11852 3332 11880
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 3605 11883 3663 11889
rect 3605 11849 3617 11883
rect 3651 11880 3663 11883
rect 4246 11880 4252 11892
rect 3651 11852 4252 11880
rect 3651 11849 3663 11852
rect 3605 11843 3663 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 4522 11880 4528 11892
rect 4479 11852 4528 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 4890 11880 4896 11892
rect 4851 11852 4896 11880
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 5442 11880 5448 11892
rect 5040 11852 5085 11880
rect 5403 11852 5448 11880
rect 5040 11840 5046 11852
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 6454 11880 6460 11892
rect 5859 11852 6460 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 6454 11840 6460 11852
rect 6512 11880 6518 11892
rect 6825 11883 6883 11889
rect 6825 11880 6837 11883
rect 6512 11852 6837 11880
rect 6512 11840 6518 11852
rect 6825 11849 6837 11852
rect 6871 11849 6883 11883
rect 6825 11843 6883 11849
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 11790 11880 11796 11892
rect 9732 11852 11796 11880
rect 9732 11840 9738 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12897 11883 12955 11889
rect 12897 11849 12909 11883
rect 12943 11880 12955 11883
rect 13170 11880 13176 11892
rect 12943 11852 13176 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13596 11852 13921 11880
rect 13596 11840 13602 11852
rect 13909 11849 13921 11852
rect 13955 11880 13967 11883
rect 14274 11880 14280 11892
rect 13955 11852 14280 11880
rect 13955 11849 13967 11852
rect 13909 11843 13967 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 14424 11852 14933 11880
rect 14424 11840 14430 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 15378 11880 15384 11892
rect 15339 11852 15384 11880
rect 14921 11843 14979 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 16025 11883 16083 11889
rect 16025 11880 16037 11883
rect 15712 11852 16037 11880
rect 15712 11840 15718 11852
rect 16025 11849 16037 11852
rect 16071 11849 16083 11883
rect 16482 11880 16488 11892
rect 16443 11852 16488 11880
rect 16025 11843 16083 11849
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 16945 11883 17003 11889
rect 16945 11880 16957 11883
rect 16724 11852 16957 11880
rect 16724 11840 16730 11852
rect 16945 11849 16957 11852
rect 16991 11849 17003 11883
rect 17402 11880 17408 11892
rect 17363 11852 17408 11880
rect 16945 11843 17003 11849
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 18322 11880 18328 11892
rect 18283 11852 18328 11880
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 19978 11880 19984 11892
rect 18656 11852 19984 11880
rect 18656 11840 18662 11852
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20073 11883 20131 11889
rect 20073 11849 20085 11883
rect 20119 11880 20131 11883
rect 20346 11880 20352 11892
rect 20119 11852 20352 11880
rect 20119 11849 20131 11852
rect 20073 11843 20131 11849
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 21082 11840 21088 11892
rect 21140 11880 21146 11892
rect 21140 11852 22876 11880
rect 21140 11840 21146 11852
rect 4154 11772 4160 11824
rect 4212 11812 4218 11824
rect 4338 11812 4344 11824
rect 4212 11784 4344 11812
rect 4212 11772 4218 11784
rect 4338 11772 4344 11784
rect 4396 11772 4402 11824
rect 5905 11815 5963 11821
rect 5905 11781 5917 11815
rect 5951 11812 5963 11815
rect 7374 11812 7380 11824
rect 5951 11784 7380 11812
rect 5951 11781 5963 11784
rect 5905 11775 5963 11781
rect 7374 11772 7380 11784
rect 7432 11812 7438 11824
rect 7938 11815 7996 11821
rect 7938 11812 7950 11815
rect 7432 11784 7950 11812
rect 7432 11772 7438 11784
rect 7938 11781 7950 11784
rect 7984 11781 7996 11815
rect 7938 11775 7996 11781
rect 10812 11815 10870 11821
rect 10812 11781 10824 11815
rect 10858 11812 10870 11815
rect 11330 11812 11336 11824
rect 10858 11784 11336 11812
rect 10858 11781 10870 11784
rect 10812 11775 10870 11781
rect 11330 11772 11336 11784
rect 11388 11772 11394 11824
rect 12986 11772 12992 11824
rect 13044 11812 13050 11824
rect 13262 11812 13268 11824
rect 13044 11784 13268 11812
rect 13044 11772 13050 11784
rect 13262 11772 13268 11784
rect 13320 11812 13326 11824
rect 14292 11812 14320 11840
rect 14461 11815 14519 11821
rect 14461 11812 14473 11815
rect 13320 11784 13584 11812
rect 14292 11784 14473 11812
rect 13320 11772 13326 11784
rect 3142 11744 3148 11756
rect 3103 11716 3148 11744
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 3436 11608 3464 11707
rect 3602 11704 3608 11756
rect 3660 11744 3666 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3660 11716 3985 11744
rect 3660 11704 3666 11716
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 4246 11744 4252 11756
rect 4111 11716 4252 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 11773 11747 11831 11753
rect 11773 11744 11785 11747
rect 10376 11716 11785 11744
rect 10376 11704 10382 11716
rect 11773 11713 11785 11716
rect 11819 11744 11831 11747
rect 12802 11744 12808 11756
rect 11819 11716 12808 11744
rect 11819 11713 11831 11716
rect 11773 11707 11831 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 13136 11716 13369 11744
rect 13136 11704 13142 11716
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11676 3942 11688
rect 4154 11676 4160 11688
rect 3936 11648 4160 11676
rect 3936 11636 3942 11648
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 5074 11676 5080 11688
rect 5035 11648 5080 11676
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 6086 11676 6092 11688
rect 6047 11648 6092 11676
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 11103 11648 11253 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 11241 11645 11253 11648
rect 11287 11676 11299 11679
rect 11514 11676 11520 11688
rect 11287 11648 11520 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 4525 11611 4583 11617
rect 4525 11608 4537 11611
rect 3436 11580 4537 11608
rect 4525 11577 4537 11580
rect 4571 11577 4583 11611
rect 4525 11571 4583 11577
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8220 11540 8248 11639
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 13556 11685 13584 11784
rect 14461 11781 14473 11784
rect 14507 11812 14519 11815
rect 14553 11815 14611 11821
rect 14553 11812 14565 11815
rect 14507 11784 14565 11812
rect 14507 11781 14519 11784
rect 14461 11775 14519 11781
rect 14553 11781 14565 11784
rect 14599 11812 14611 11815
rect 14737 11815 14795 11821
rect 14737 11812 14749 11815
rect 14599 11784 14749 11812
rect 14599 11781 14611 11784
rect 14553 11775 14611 11781
rect 14737 11781 14749 11784
rect 14783 11781 14795 11815
rect 14737 11775 14795 11781
rect 15289 11815 15347 11821
rect 15289 11781 15301 11815
rect 15335 11812 15347 11815
rect 15930 11812 15936 11824
rect 15335 11784 15936 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 15930 11772 15936 11784
rect 15988 11772 15994 11824
rect 17681 11815 17739 11821
rect 17681 11812 17693 11815
rect 16868 11784 17693 11812
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 16117 11747 16175 11753
rect 13688 11716 15976 11744
rect 13688 11704 13694 11716
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 13464 11608 13492 11639
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 15948 11685 15976 11716
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16206 11744 16212 11756
rect 16163 11716 16212 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 16868 11685 16896 11784
rect 17681 11781 17693 11784
rect 17727 11812 17739 11815
rect 18230 11812 18236 11824
rect 17727 11784 18236 11812
rect 17727 11781 17739 11784
rect 17681 11775 17739 11781
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 18782 11772 18788 11824
rect 18840 11812 18846 11824
rect 20990 11812 20996 11824
rect 18840 11784 20996 11812
rect 18840 11772 18846 11784
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 21634 11812 21640 11824
rect 21192 11784 21640 11812
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11744 17923 11747
rect 17954 11744 17960 11756
rect 17911 11716 17960 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11744 18199 11747
rect 18322 11744 18328 11756
rect 18187 11716 18328 11744
rect 18187 11713 18199 11716
rect 18141 11707 18199 11713
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 13780 11648 15485 11676
rect 13780 11636 13786 11648
rect 15473 11645 15485 11648
rect 15519 11645 15531 11679
rect 15473 11639 15531 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 12820 11580 13492 11608
rect 8297 11543 8355 11549
rect 8297 11540 8309 11543
rect 8076 11512 8309 11540
rect 8076 11500 8082 11512
rect 8297 11509 8309 11512
rect 8343 11509 8355 11543
rect 8297 11503 8355 11509
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 12820 11540 12848 11580
rect 12986 11540 12992 11552
rect 11848 11512 12848 11540
rect 12947 11512 12992 11540
rect 11848 11500 11854 11512
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 15488 11540 15516 11639
rect 15948 11608 15976 11639
rect 16942 11636 16948 11688
rect 17000 11676 17006 11688
rect 18156 11676 18184 11707
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11713 18475 11747
rect 18690 11744 18696 11756
rect 18651 11716 18696 11744
rect 18417 11707 18475 11713
rect 17000 11648 18184 11676
rect 17000 11636 17006 11648
rect 17497 11611 17555 11617
rect 17497 11608 17509 11611
rect 15948 11580 17509 11608
rect 17497 11577 17509 11580
rect 17543 11577 17555 11611
rect 18432 11608 18460 11707
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 18960 11747 19018 11753
rect 18960 11713 18972 11747
rect 19006 11744 19018 11747
rect 19242 11744 19248 11756
rect 19006 11716 19248 11744
rect 19006 11713 19018 11716
rect 18960 11707 19018 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 21192 11744 21220 11784
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 22189 11815 22247 11821
rect 22189 11781 22201 11815
rect 22235 11812 22247 11815
rect 22278 11812 22284 11824
rect 22235 11784 22284 11812
rect 22235 11781 22247 11784
rect 22189 11775 22247 11781
rect 22278 11772 22284 11784
rect 22336 11772 22342 11824
rect 22646 11812 22652 11824
rect 22607 11784 22652 11812
rect 22646 11772 22652 11784
rect 22704 11772 22710 11824
rect 22848 11821 22876 11852
rect 22833 11815 22891 11821
rect 22833 11781 22845 11815
rect 22879 11781 22891 11815
rect 22833 11775 22891 11781
rect 20005 11716 21220 11744
rect 18432 11580 18736 11608
rect 17497 11571 17555 11577
rect 16758 11540 16764 11552
rect 15488 11512 16764 11540
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18598 11540 18604 11552
rect 18559 11512 18604 11540
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 18708 11540 18736 11580
rect 20005 11540 20033 11716
rect 21266 11704 21272 11756
rect 21324 11753 21330 11756
rect 21324 11744 21336 11753
rect 21542 11744 21548 11756
rect 21324 11716 21369 11744
rect 21503 11716 21548 11744
rect 21324 11707 21336 11716
rect 21324 11704 21330 11707
rect 21542 11704 21548 11716
rect 21600 11744 21606 11756
rect 23017 11747 23075 11753
rect 23017 11744 23029 11747
rect 21600 11716 23029 11744
rect 21600 11704 21606 11716
rect 23017 11713 23029 11716
rect 23063 11713 23075 11747
rect 23017 11707 23075 11713
rect 22281 11679 22339 11685
rect 22281 11645 22293 11679
rect 22327 11645 22339 11679
rect 22281 11639 22339 11645
rect 18708 11512 20033 11540
rect 20165 11543 20223 11549
rect 20165 11509 20177 11543
rect 20211 11540 20223 11543
rect 20346 11540 20352 11552
rect 20211 11512 20352 11540
rect 20211 11509 20223 11512
rect 20165 11503 20223 11509
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 21634 11500 21640 11552
rect 21692 11540 21698 11552
rect 21821 11543 21879 11549
rect 21821 11540 21833 11543
rect 21692 11512 21833 11540
rect 21692 11500 21698 11512
rect 21821 11509 21833 11512
rect 21867 11509 21879 11543
rect 22296 11540 22324 11639
rect 22370 11636 22376 11688
rect 22428 11676 22434 11688
rect 22428 11648 22473 11676
rect 22428 11636 22434 11648
rect 22554 11540 22560 11552
rect 22296 11512 22560 11540
rect 21821 11503 21879 11509
rect 22554 11500 22560 11512
rect 22612 11500 22618 11552
rect 1104 11450 23460 11472
rect 1104 11398 3749 11450
rect 3801 11398 3813 11450
rect 3865 11398 3877 11450
rect 3929 11398 3941 11450
rect 3993 11398 4005 11450
rect 4057 11398 9347 11450
rect 9399 11398 9411 11450
rect 9463 11398 9475 11450
rect 9527 11398 9539 11450
rect 9591 11398 9603 11450
rect 9655 11398 14945 11450
rect 14997 11398 15009 11450
rect 15061 11398 15073 11450
rect 15125 11398 15137 11450
rect 15189 11398 15201 11450
rect 15253 11398 20543 11450
rect 20595 11398 20607 11450
rect 20659 11398 20671 11450
rect 20723 11398 20735 11450
rect 20787 11398 20799 11450
rect 20851 11398 23460 11450
rect 1104 11376 23460 11398
rect 7190 11336 7196 11348
rect 7151 11308 7196 11336
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 10410 11336 10416 11348
rect 10371 11308 10416 11336
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 11974 11336 11980 11348
rect 11935 11308 11980 11336
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 13538 11336 13544 11348
rect 13499 11308 13544 11336
rect 13538 11296 13544 11308
rect 13596 11336 13602 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 13596 11308 13645 11336
rect 13596 11296 13602 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 16850 11336 16856 11348
rect 15703 11308 16856 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 16850 11296 16856 11308
rect 16908 11336 16914 11348
rect 17034 11336 17040 11348
rect 16908 11308 17040 11336
rect 16908 11296 16914 11308
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 19242 11336 19248 11348
rect 18012 11308 18644 11336
rect 19155 11308 19248 11336
rect 18012 11296 18018 11308
rect 5718 11268 5724 11280
rect 5679 11240 5724 11268
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 10318 11268 10324 11280
rect 10279 11240 10324 11268
rect 10318 11228 10324 11240
rect 10376 11228 10382 11280
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 4338 11200 4344 11212
rect 4203 11172 4344 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 4801 11203 4859 11209
rect 4801 11200 4813 11203
rect 4764 11172 4813 11200
rect 4764 11160 4770 11172
rect 4801 11169 4813 11172
rect 4847 11169 4859 11203
rect 4801 11163 4859 11169
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 13446 11200 13452 11212
rect 13403 11172 13452 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 5074 11132 5080 11144
rect 5035 11104 5080 11132
rect 5074 11092 5080 11104
rect 5132 11092 5138 11144
rect 7098 11132 7104 11144
rect 7059 11104 7104 11132
rect 7098 11092 7104 11104
rect 7156 11132 7162 11144
rect 8018 11132 8024 11144
rect 7156 11104 8024 11132
rect 7156 11092 7162 11104
rect 8018 11092 8024 11104
rect 8076 11132 8082 11144
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8076 11104 8585 11132
rect 8076 11092 8082 11104
rect 8573 11101 8585 11104
rect 8619 11132 8631 11135
rect 8665 11135 8723 11141
rect 8665 11132 8677 11135
rect 8619 11104 8677 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 8665 11101 8677 11104
rect 8711 11132 8723 11135
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8711 11104 8953 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9208 11135 9266 11141
rect 9208 11101 9220 11135
rect 9254 11132 9266 11135
rect 9674 11132 9680 11144
rect 9254 11104 9680 11132
rect 9254 11101 9266 11104
rect 9208 11095 9266 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 12066 11132 12072 11144
rect 11839 11104 12072 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 12066 11092 12072 11104
rect 12124 11132 12130 11144
rect 13372 11132 13400 11163
rect 13446 11160 13452 11172
rect 13504 11200 13510 11212
rect 13556 11200 13584 11296
rect 15470 11268 15476 11280
rect 15431 11240 15476 11268
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 18616 11268 18644 11308
rect 19242 11296 19248 11308
rect 19300 11336 19306 11348
rect 21453 11339 21511 11345
rect 19300 11308 20760 11336
rect 19300 11296 19306 11308
rect 19058 11268 19064 11280
rect 18616 11240 19064 11268
rect 19058 11228 19064 11240
rect 19116 11268 19122 11280
rect 19334 11268 19340 11280
rect 19116 11240 19340 11268
rect 19116 11228 19122 11240
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 13504 11172 14105 11200
rect 13504 11160 13510 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15654 11200 15660 11212
rect 15160 11172 15660 11200
rect 15160 11160 15166 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 17037 11203 17095 11209
rect 17037 11169 17049 11203
rect 17083 11200 17095 11203
rect 17310 11200 17316 11212
rect 17083 11172 17316 11200
rect 17083 11169 17095 11172
rect 17037 11163 17095 11169
rect 17310 11160 17316 11172
rect 17368 11200 17374 11212
rect 17681 11203 17739 11209
rect 17681 11200 17693 11203
rect 17368 11172 17693 11200
rect 17368 11160 17374 11172
rect 17681 11169 17693 11172
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 12124 11104 13400 11132
rect 14360 11135 14418 11141
rect 12124 11092 12130 11104
rect 14360 11101 14372 11135
rect 14406 11132 14418 11135
rect 14642 11132 14648 11144
rect 14406 11104 14648 11132
rect 14406 11101 14418 11104
rect 14360 11095 14418 11101
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 17129 11135 17187 11141
rect 16592 11104 16896 11132
rect 4249 11067 4307 11073
rect 4249 11033 4261 11067
rect 4295 11064 4307 11067
rect 5442 11064 5448 11076
rect 4295 11036 5448 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 6454 11024 6460 11076
rect 6512 11064 6518 11076
rect 6834 11067 6892 11073
rect 6834 11064 6846 11067
rect 6512 11036 6846 11064
rect 6512 11024 6518 11036
rect 6834 11033 6846 11036
rect 6880 11033 6892 11067
rect 6834 11027 6892 11033
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 8306 11067 8364 11073
rect 8306 11064 8318 11067
rect 7064 11036 8318 11064
rect 7064 11024 7070 11036
rect 8306 11033 8318 11036
rect 8352 11033 8364 11067
rect 8306 11027 8364 11033
rect 11548 11067 11606 11073
rect 11548 11033 11560 11067
rect 11594 11064 11606 11067
rect 11974 11064 11980 11076
rect 11594 11036 11980 11064
rect 11594 11033 11606 11036
rect 11548 11027 11606 11033
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 13078 11024 13084 11076
rect 13136 11073 13142 11076
rect 13136 11064 13148 11073
rect 13909 11067 13967 11073
rect 13136 11036 13181 11064
rect 13136 11027 13148 11036
rect 13909 11033 13921 11067
rect 13955 11064 13967 11067
rect 16592 11064 16620 11104
rect 13955 11036 16620 11064
rect 13955 11033 13967 11036
rect 13909 11027 13967 11033
rect 13136 11024 13142 11027
rect 16666 11024 16672 11076
rect 16724 11064 16730 11076
rect 16770 11067 16828 11073
rect 16770 11064 16782 11067
rect 16724 11036 16782 11064
rect 16724 11024 16730 11036
rect 16770 11033 16782 11036
rect 16816 11033 16828 11067
rect 16868 11064 16896 11104
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 19334 11132 19340 11144
rect 17175 11104 19340 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 17144 11064 17172 11095
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 20346 11092 20352 11144
rect 20404 11141 20410 11144
rect 20404 11132 20416 11141
rect 20622 11132 20628 11144
rect 20404 11104 20484 11132
rect 20583 11104 20628 11132
rect 20404 11095 20416 11104
rect 20404 11092 20410 11095
rect 17586 11064 17592 11076
rect 16868 11036 17172 11064
rect 17547 11036 17592 11064
rect 16770 11027 16828 11033
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 17948 11067 18006 11073
rect 17948 11033 17960 11067
rect 17994 11064 18006 11067
rect 19242 11064 19248 11076
rect 17994 11036 19248 11064
rect 17994 11033 18006 11036
rect 17948 11027 18006 11033
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 20456 11064 20484 11104
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 20732 11132 20760 11308
rect 21453 11305 21465 11339
rect 21499 11336 21511 11339
rect 22002 11336 22008 11348
rect 21499 11308 22008 11336
rect 21499 11305 21511 11308
rect 21453 11299 21511 11305
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22278 11228 22284 11280
rect 22336 11268 22342 11280
rect 22336 11240 22381 11268
rect 22336 11228 22342 11240
rect 20901 11203 20959 11209
rect 20901 11169 20913 11203
rect 20947 11200 20959 11203
rect 21726 11200 21732 11212
rect 20947 11172 21732 11200
rect 20947 11169 20959 11172
rect 20901 11163 20959 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 22830 11200 22836 11212
rect 22791 11172 22836 11200
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 23014 11200 23020 11212
rect 22975 11172 23020 11200
rect 23014 11160 23020 11172
rect 23072 11160 23078 11212
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 20732 11104 21097 11132
rect 21085 11101 21097 11104
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 21358 11092 21364 11144
rect 21416 11132 21422 11144
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 21416 11104 22753 11132
rect 21416 11092 21422 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 20993 11067 21051 11073
rect 20993 11064 21005 11067
rect 20456 11036 21005 11064
rect 20993 11033 21005 11036
rect 21039 11033 21051 11067
rect 20993 11027 21051 11033
rect 21266 11024 21272 11076
rect 21324 11064 21330 11076
rect 21913 11067 21971 11073
rect 21913 11064 21925 11067
rect 21324 11036 21925 11064
rect 21324 11024 21330 11036
rect 21913 11033 21925 11036
rect 21959 11033 21971 11067
rect 21913 11027 21971 11033
rect 4338 10956 4344 11008
rect 4396 10996 4402 11008
rect 4396 10968 4441 10996
rect 4396 10956 4402 10968
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4709 10999 4767 11005
rect 4709 10996 4721 10999
rect 4580 10968 4721 10996
rect 4580 10956 4586 10968
rect 4709 10965 4721 10968
rect 4755 10965 4767 10999
rect 4709 10959 4767 10965
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 7742 10996 7748 11008
rect 5040 10968 7748 10996
rect 5040 10956 5046 10968
rect 7742 10956 7748 10968
rect 7800 10996 7806 11008
rect 10318 10996 10324 11008
rect 7800 10968 10324 10996
rect 7800 10956 7806 10968
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10996 17371 10999
rect 18506 10996 18512 11008
rect 17359 10968 18512 10996
rect 17359 10965 17371 10968
rect 17313 10959 17371 10965
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 18966 10956 18972 11008
rect 19024 10996 19030 11008
rect 19061 10999 19119 11005
rect 19061 10996 19073 10999
rect 19024 10968 19073 10996
rect 19024 10956 19030 10968
rect 19061 10965 19073 10968
rect 19107 10965 19119 10999
rect 19061 10959 19119 10965
rect 19150 10956 19156 11008
rect 19208 10996 19214 11008
rect 21821 10999 21879 11005
rect 21821 10996 21833 10999
rect 19208 10968 21833 10996
rect 19208 10956 19214 10968
rect 21821 10965 21833 10968
rect 21867 10965 21879 10999
rect 22370 10996 22376 11008
rect 22331 10968 22376 10996
rect 21821 10959 21879 10965
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 1104 10906 23460 10928
rect 1104 10854 6548 10906
rect 6600 10854 6612 10906
rect 6664 10854 6676 10906
rect 6728 10854 6740 10906
rect 6792 10854 6804 10906
rect 6856 10854 12146 10906
rect 12198 10854 12210 10906
rect 12262 10854 12274 10906
rect 12326 10854 12338 10906
rect 12390 10854 12402 10906
rect 12454 10854 17744 10906
rect 17796 10854 17808 10906
rect 17860 10854 17872 10906
rect 17924 10854 17936 10906
rect 17988 10854 18000 10906
rect 18052 10854 23460 10906
rect 1104 10832 23460 10854
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4396 10764 4629 10792
rect 4396 10752 4402 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 4982 10792 4988 10804
rect 4943 10764 4988 10792
rect 4617 10755 4675 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 12897 10795 12955 10801
rect 5828 10764 12434 10792
rect 5077 10727 5135 10733
rect 5077 10693 5089 10727
rect 5123 10724 5135 10727
rect 5828 10724 5856 10764
rect 5123 10696 5856 10724
rect 5905 10727 5963 10733
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 5905 10693 5917 10727
rect 5951 10724 5963 10727
rect 6822 10724 6828 10736
rect 5951 10696 6828 10724
rect 5951 10693 5963 10696
rect 5905 10687 5963 10693
rect 6822 10684 6828 10696
rect 6880 10684 6886 10736
rect 7033 10696 7788 10724
rect 4522 10656 4528 10668
rect 4483 10628 4528 10656
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 7033 10656 7061 10696
rect 5859 10628 7061 10656
rect 7760 10656 7788 10696
rect 7926 10684 7932 10736
rect 7984 10733 7990 10736
rect 7984 10724 7996 10733
rect 7984 10696 8029 10724
rect 7984 10687 7996 10696
rect 7984 10684 7990 10687
rect 8110 10684 8116 10736
rect 8168 10724 8174 10736
rect 11790 10733 11796 10736
rect 9094 10727 9152 10733
rect 9094 10724 9106 10727
rect 8168 10696 9106 10724
rect 8168 10684 8174 10696
rect 9094 10693 9106 10696
rect 9140 10693 9152 10727
rect 11784 10724 11796 10733
rect 11751 10696 11796 10724
rect 9094 10687 9152 10693
rect 11784 10687 11796 10696
rect 11790 10684 11796 10687
rect 11848 10684 11854 10736
rect 12406 10724 12434 10764
rect 12897 10761 12909 10795
rect 12943 10792 12955 10795
rect 13078 10792 13084 10804
rect 12943 10764 13084 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 13262 10792 13268 10804
rect 13223 10764 13268 10792
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 14826 10752 14832 10804
rect 14884 10792 14890 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 14884 10764 15025 10792
rect 14884 10752 14890 10764
rect 15013 10761 15025 10764
rect 15059 10792 15071 10795
rect 15102 10792 15108 10804
rect 15059 10764 15108 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 22554 10792 22560 10804
rect 18156 10764 21956 10792
rect 22515 10764 22560 10792
rect 14654 10727 14712 10733
rect 14654 10724 14666 10727
rect 12406 10696 14666 10724
rect 14654 10693 14666 10696
rect 14700 10724 14712 10727
rect 15378 10724 15384 10736
rect 14700 10696 15384 10724
rect 14700 10693 14712 10696
rect 14654 10687 14712 10693
rect 15378 10684 15384 10696
rect 15436 10684 15442 10736
rect 15948 10696 16436 10724
rect 10502 10656 10508 10668
rect 7760 10628 10272 10656
rect 10415 10628 10508 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 5169 10591 5227 10597
rect 5169 10588 5181 10591
rect 4764 10560 5181 10588
rect 4764 10548 4770 10560
rect 5169 10557 5181 10560
rect 5215 10557 5227 10591
rect 5169 10551 5227 10557
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 8251 10560 8861 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 8849 10557 8861 10560
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 4246 10480 4252 10532
rect 4304 10520 4310 10532
rect 4341 10523 4399 10529
rect 4341 10520 4353 10523
rect 4304 10492 4353 10520
rect 4304 10480 4310 10492
rect 4341 10489 4353 10492
rect 4387 10489 4399 10523
rect 4341 10483 4399 10489
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 6012 10520 6040 10551
rect 6822 10520 6828 10532
rect 5132 10492 6040 10520
rect 6783 10492 6828 10520
rect 5132 10480 5138 10492
rect 6822 10480 6828 10492
rect 6880 10480 6886 10532
rect 8220 10464 8248 10551
rect 5902 10412 5908 10464
rect 5960 10452 5966 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 5960 10424 6653 10452
rect 5960 10412 5966 10424
rect 6641 10421 6653 10424
rect 6687 10452 6699 10455
rect 7098 10452 7104 10464
rect 6687 10424 7104 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 7098 10412 7104 10424
rect 7156 10452 7162 10464
rect 8202 10452 8208 10464
rect 7156 10424 8208 10452
rect 7156 10412 7162 10424
rect 8202 10412 8208 10424
rect 8260 10452 8266 10464
rect 8297 10455 8355 10461
rect 8297 10452 8309 10455
rect 8260 10424 8309 10452
rect 8260 10412 8266 10424
rect 8297 10421 8309 10424
rect 8343 10421 8355 10455
rect 8864 10452 8892 10551
rect 10244 10529 10272 10628
rect 10502 10616 10508 10628
rect 10560 10656 10566 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10560 10628 10701 10656
rect 10560 10616 10566 10628
rect 10689 10625 10701 10628
rect 10735 10656 10747 10659
rect 11514 10656 11520 10668
rect 10735 10628 11520 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 11514 10616 11520 10628
rect 11572 10656 11578 10668
rect 12066 10656 12072 10668
rect 11572 10628 12072 10656
rect 11572 10616 11578 10628
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 13630 10656 13636 10668
rect 13403 10628 13636 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 13814 10656 13820 10668
rect 13740 10628 13820 10656
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10588 13139 10591
rect 13446 10588 13452 10600
rect 13127 10560 13452 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13446 10548 13452 10560
rect 13504 10588 13510 10600
rect 13740 10588 13768 10628
rect 13814 10616 13820 10628
rect 13872 10656 13878 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 13872 10628 14933 10656
rect 13872 10616 13878 10628
rect 14921 10625 14933 10628
rect 14967 10656 14979 10659
rect 15654 10656 15660 10668
rect 14967 10628 15660 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 15654 10616 15660 10628
rect 15712 10656 15718 10668
rect 15948 10656 15976 10696
rect 16114 10656 16120 10668
rect 16172 10665 16178 10668
rect 16408 10665 16436 10696
rect 15712 10628 15976 10656
rect 16084 10628 16120 10656
rect 15712 10616 15718 10628
rect 16114 10616 16120 10628
rect 16172 10619 16184 10665
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10656 16451 10659
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16439 10628 16681 10656
rect 16439 10625 16451 10628
rect 16393 10619 16451 10625
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 16936 10659 16994 10665
rect 16936 10625 16948 10659
rect 16982 10656 16994 10659
rect 17218 10656 17224 10668
rect 16982 10628 17224 10656
rect 16982 10625 16994 10628
rect 16936 10619 16994 10625
rect 16172 10616 16178 10619
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 18156 10656 18184 10764
rect 18233 10727 18291 10733
rect 18233 10693 18245 10727
rect 18279 10724 18291 10727
rect 19426 10724 19432 10736
rect 18279 10696 19432 10724
rect 18279 10693 18291 10696
rect 18233 10687 18291 10693
rect 18616 10665 18644 10696
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 20622 10684 20628 10736
rect 20680 10724 20686 10736
rect 21542 10724 21548 10736
rect 20680 10696 21548 10724
rect 20680 10684 20686 10696
rect 21542 10684 21548 10696
rect 21600 10684 21606 10736
rect 18325 10659 18383 10665
rect 18325 10656 18337 10659
rect 18156 10628 18337 10656
rect 18325 10625 18337 10628
rect 18371 10625 18383 10659
rect 18325 10619 18383 10625
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18868 10659 18926 10665
rect 18868 10656 18880 10659
rect 18601 10619 18659 10625
rect 18708 10628 18880 10656
rect 18708 10588 18736 10628
rect 18868 10625 18880 10628
rect 18914 10656 18926 10659
rect 19150 10656 19156 10668
rect 18914 10628 19156 10656
rect 18914 10625 18926 10628
rect 18868 10619 18926 10625
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19444 10656 19472 10684
rect 20346 10665 20352 10668
rect 19444 10628 20033 10656
rect 13504 10560 13768 10588
rect 18064 10560 18736 10588
rect 20005 10588 20033 10628
rect 20340 10619 20352 10665
rect 20404 10656 20410 10668
rect 21928 10656 21956 10764
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 22094 10684 22100 10736
rect 22152 10724 22158 10736
rect 23017 10727 23075 10733
rect 22152 10696 22197 10724
rect 22152 10684 22158 10696
rect 23017 10693 23029 10727
rect 23063 10724 23075 10727
rect 23382 10724 23388 10736
rect 23063 10696 23388 10724
rect 23063 10693 23075 10696
rect 23017 10687 23075 10693
rect 23382 10684 23388 10696
rect 23440 10684 23446 10736
rect 22189 10659 22247 10665
rect 20404 10628 20440 10656
rect 21928 10628 22094 10656
rect 20346 10616 20352 10619
rect 20404 10616 20410 10628
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 20005 10560 20085 10588
rect 13504 10548 13510 10560
rect 18064 10529 18092 10560
rect 20073 10557 20085 10560
rect 20119 10557 20131 10591
rect 20073 10551 20131 10557
rect 21726 10548 21732 10600
rect 21784 10588 21790 10600
rect 21913 10591 21971 10597
rect 21913 10588 21925 10591
rect 21784 10560 21925 10588
rect 21784 10548 21790 10560
rect 21913 10557 21925 10560
rect 21959 10557 21971 10591
rect 22066 10588 22094 10628
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22278 10656 22284 10668
rect 22235 10628 22284 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 22649 10591 22707 10597
rect 22649 10588 22661 10591
rect 22066 10560 22661 10588
rect 21913 10551 21971 10557
rect 22649 10557 22661 10560
rect 22695 10557 22707 10591
rect 22649 10551 22707 10557
rect 10229 10523 10287 10529
rect 10229 10489 10241 10523
rect 10275 10520 10287 10523
rect 18049 10523 18107 10529
rect 10275 10492 10732 10520
rect 10275 10489 10287 10492
rect 10229 10483 10287 10489
rect 10502 10452 10508 10464
rect 8864 10424 10508 10452
rect 8297 10415 8355 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 10704 10452 10732 10492
rect 18049 10489 18061 10523
rect 18095 10489 18107 10523
rect 22848 10520 22876 10619
rect 18049 10483 18107 10489
rect 21468 10492 22876 10520
rect 21468 10464 21496 10492
rect 13170 10452 13176 10464
rect 10704 10424 13176 10452
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 13541 10455 13599 10461
rect 13541 10452 13553 10455
rect 13412 10424 13553 10452
rect 13412 10412 13418 10424
rect 13541 10421 13553 10424
rect 13587 10421 13599 10455
rect 13541 10415 13599 10421
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 19794 10452 19800 10464
rect 18555 10424 19800 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 19794 10412 19800 10424
rect 19852 10412 19858 10464
rect 19981 10455 20039 10461
rect 19981 10421 19993 10455
rect 20027 10452 20039 10455
rect 21266 10452 21272 10464
rect 20027 10424 21272 10452
rect 20027 10421 20039 10424
rect 19981 10415 20039 10421
rect 21266 10412 21272 10424
rect 21324 10412 21330 10464
rect 21450 10452 21456 10464
rect 21411 10424 21456 10452
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 22094 10452 22100 10464
rect 21600 10424 22100 10452
rect 21600 10412 21606 10424
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 1104 10362 23460 10384
rect 1104 10310 3749 10362
rect 3801 10310 3813 10362
rect 3865 10310 3877 10362
rect 3929 10310 3941 10362
rect 3993 10310 4005 10362
rect 4057 10310 9347 10362
rect 9399 10310 9411 10362
rect 9463 10310 9475 10362
rect 9527 10310 9539 10362
rect 9591 10310 9603 10362
rect 9655 10310 14945 10362
rect 14997 10310 15009 10362
rect 15061 10310 15073 10362
rect 15125 10310 15137 10362
rect 15189 10310 15201 10362
rect 15253 10310 20543 10362
rect 20595 10310 20607 10362
rect 20659 10310 20671 10362
rect 20723 10310 20735 10362
rect 20787 10310 20799 10362
rect 20851 10310 23460 10362
rect 1104 10288 23460 10310
rect 3602 10248 3608 10260
rect 3563 10220 3608 10248
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 4614 10248 4620 10260
rect 4571 10220 4620 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 7282 10248 7288 10260
rect 7195 10220 7288 10248
rect 7282 10208 7288 10220
rect 7340 10248 7346 10260
rect 10502 10248 10508 10260
rect 7340 10220 9168 10248
rect 10463 10220 10508 10248
rect 7340 10208 7346 10220
rect 3973 10115 4031 10121
rect 3973 10081 3985 10115
rect 4019 10112 4031 10115
rect 4154 10112 4160 10124
rect 4019 10084 4160 10112
rect 4019 10081 4031 10084
rect 3973 10075 4031 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 5350 10112 5356 10124
rect 5092 10084 5356 10112
rect 5092 10056 5120 10084
rect 5350 10072 5356 10084
rect 5408 10112 5414 10124
rect 5629 10115 5687 10121
rect 5629 10112 5641 10115
rect 5408 10084 5641 10112
rect 5408 10072 5414 10084
rect 5629 10081 5641 10084
rect 5675 10081 5687 10115
rect 5902 10112 5908 10124
rect 5863 10084 5908 10112
rect 5629 10075 5687 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 3418 10044 3424 10056
rect 3379 10016 3424 10044
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5074 10044 5080 10056
rect 4939 10016 5080 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5583 10016 7696 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 3786 9936 3792 9988
rect 3844 9976 3850 9988
rect 4157 9979 4215 9985
rect 4157 9976 4169 9979
rect 3844 9948 4169 9976
rect 3844 9936 3850 9948
rect 4157 9945 4169 9948
rect 4203 9945 4215 9979
rect 4157 9939 4215 9945
rect 4430 9936 4436 9988
rect 4488 9976 4494 9988
rect 6178 9985 6184 9988
rect 4709 9979 4767 9985
rect 4709 9976 4721 9979
rect 4488 9948 4721 9976
rect 4488 9936 4494 9948
rect 4709 9945 4721 9948
rect 4755 9945 4767 9979
rect 6172 9976 6184 9985
rect 6139 9948 6184 9976
rect 4709 9939 4767 9945
rect 6172 9939 6184 9948
rect 6178 9936 6184 9939
rect 6236 9936 6242 9988
rect 7668 9976 7696 10016
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 8260 10016 8769 10044
rect 8260 10004 8266 10016
rect 8757 10013 8769 10016
rect 8803 10013 8815 10047
rect 8757 10007 8815 10013
rect 8490 9979 8548 9985
rect 8490 9976 8502 9979
rect 7668 9948 8502 9976
rect 8490 9945 8502 9948
rect 8536 9976 8548 9979
rect 9140 9976 9168 10220
rect 10502 10208 10508 10220
rect 10560 10248 10566 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10560 10220 10609 10248
rect 10560 10208 10566 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10248 12955 10251
rect 20346 10248 20352 10260
rect 12943 10220 20352 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 10318 10140 10324 10192
rect 10376 10180 10382 10192
rect 10376 10152 12434 10180
rect 10376 10140 10382 10152
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 11664 10084 11713 10112
rect 11664 10072 11670 10084
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 12406 10112 12434 10152
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13814 10180 13820 10192
rect 13228 10152 13676 10180
rect 13775 10152 13820 10180
rect 13228 10140 13234 10152
rect 13354 10112 13360 10124
rect 12406 10084 13360 10112
rect 11701 10075 11759 10081
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 13538 10112 13544 10124
rect 13499 10084 13544 10112
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13648 10112 13676 10152
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 15378 10140 15384 10192
rect 15436 10180 15442 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15436 10152 15485 10180
rect 15436 10140 15442 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 15654 10180 15660 10192
rect 15615 10152 15660 10180
rect 15473 10143 15531 10149
rect 15654 10140 15660 10152
rect 15712 10180 15718 10192
rect 15749 10183 15807 10189
rect 15749 10180 15761 10183
rect 15712 10152 15761 10180
rect 15712 10140 15718 10152
rect 15749 10149 15761 10152
rect 15795 10149 15807 10183
rect 15749 10143 15807 10149
rect 15933 10183 15991 10189
rect 15933 10149 15945 10183
rect 15979 10180 15991 10183
rect 16114 10180 16120 10192
rect 15979 10152 16120 10180
rect 15979 10149 15991 10152
rect 15933 10143 15991 10149
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 18414 10140 18420 10192
rect 18472 10180 18478 10192
rect 18472 10152 18828 10180
rect 18472 10140 18478 10152
rect 16577 10115 16635 10121
rect 13648 10084 14228 10112
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 10502 10044 10508 10056
rect 10367 10016 10508 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 12986 10044 12992 10056
rect 12023 10016 12992 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13872 10016 14105 10044
rect 13872 10004 13878 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14200 10044 14228 10084
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 16850 10112 16856 10124
rect 16623 10084 16856 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 18800 10121 18828 10152
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10081 18843 10115
rect 18785 10075 18843 10081
rect 14349 10047 14407 10053
rect 14349 10044 14361 10047
rect 14200 10016 14361 10044
rect 14093 10007 14151 10013
rect 14349 10013 14361 10016
rect 14395 10013 14407 10047
rect 14349 10007 14407 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 17034 10044 17040 10056
rect 16807 10016 17040 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 17034 10004 17040 10016
rect 17092 10004 17098 10056
rect 19076 10053 19104 10220
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 20456 10220 22140 10248
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10044 19303 10047
rect 19334 10044 19340 10056
rect 19291 10016 19340 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 10054 9979 10112 9985
rect 10054 9976 10066 9979
rect 8536 9948 8984 9976
rect 9140 9948 10066 9976
rect 8536 9945 8548 9948
rect 8490 9939 8548 9945
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3568 9880 4077 9908
rect 3568 9868 3574 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 5074 9908 5080 9920
rect 5035 9880 5080 9908
rect 4065 9871 4123 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9908 5503 9911
rect 6454 9908 6460 9920
rect 5491 9880 6460 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 6454 9868 6460 9880
rect 6512 9908 6518 9920
rect 8956 9917 8984 9948
rect 10054 9945 10066 9948
rect 10100 9945 10112 9979
rect 10054 9939 10112 9945
rect 11885 9979 11943 9985
rect 11885 9945 11897 9979
rect 11931 9976 11943 9979
rect 12713 9979 12771 9985
rect 11931 9948 12664 9976
rect 11931 9945 11943 9948
rect 11885 9939 11943 9945
rect 7377 9911 7435 9917
rect 7377 9908 7389 9911
rect 6512 9880 7389 9908
rect 6512 9868 6518 9880
rect 7377 9877 7389 9880
rect 7423 9877 7435 9911
rect 7377 9871 7435 9877
rect 8941 9911 8999 9917
rect 8941 9877 8953 9911
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 12345 9911 12403 9917
rect 12345 9908 12357 9911
rect 12124 9880 12357 9908
rect 12124 9868 12130 9880
rect 12345 9877 12357 9880
rect 12391 9877 12403 9911
rect 12636 9908 12664 9948
rect 12713 9945 12725 9979
rect 12759 9976 12771 9979
rect 13262 9976 13268 9988
rect 12759 9948 13268 9976
rect 12759 9945 12771 9948
rect 12713 9939 12771 9945
rect 13262 9936 13268 9948
rect 13320 9976 13326 9988
rect 13832 9976 13860 10004
rect 13320 9948 13860 9976
rect 18172 9979 18230 9985
rect 13320 9936 13326 9948
rect 18172 9945 18184 9979
rect 18218 9976 18230 9979
rect 18322 9976 18328 9988
rect 18218 9948 18328 9976
rect 18218 9945 18230 9948
rect 18172 9939 18230 9945
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 18432 9976 18460 10007
rect 19260 9976 19288 10007
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 19518 10053 19524 10056
rect 19512 10007 19524 10053
rect 19576 10044 19582 10056
rect 19576 10016 19612 10044
rect 19518 10004 19524 10007
rect 19576 10004 19582 10016
rect 19794 10004 19800 10056
rect 19852 10044 19858 10056
rect 20456 10044 20484 10220
rect 20714 10180 20720 10192
rect 20675 10152 20720 10180
rect 20714 10140 20720 10152
rect 20772 10140 20778 10192
rect 22112 10180 22140 10220
rect 22112 10152 22324 10180
rect 22296 10112 22324 10152
rect 22741 10115 22799 10121
rect 22741 10112 22753 10115
rect 22296 10084 22753 10112
rect 22741 10081 22753 10084
rect 22787 10081 22799 10115
rect 22741 10075 22799 10081
rect 19852 10016 20484 10044
rect 19852 10004 19858 10016
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 21830 10047 21888 10053
rect 21830 10044 21842 10047
rect 21508 10016 21842 10044
rect 21508 10004 21514 10016
rect 21830 10013 21842 10016
rect 21876 10013 21888 10047
rect 22094 10044 22100 10056
rect 22055 10016 22100 10044
rect 21830 10007 21888 10013
rect 22094 10004 22100 10016
rect 22152 10044 22158 10056
rect 22646 10044 22652 10056
rect 22152 10016 22416 10044
rect 22607 10016 22652 10044
rect 22152 10004 22158 10016
rect 22278 9976 22284 9988
rect 18432 9948 19288 9976
rect 19352 9948 22284 9976
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12636 9880 13001 9908
rect 12345 9871 12403 9877
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 13354 9908 13360 9920
rect 13315 9880 13360 9908
rect 12989 9871 13047 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 13446 9868 13452 9920
rect 13504 9908 13510 9920
rect 16942 9908 16948 9920
rect 13504 9880 13549 9908
rect 16903 9880 16948 9908
rect 13504 9868 13510 9880
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 17037 9911 17095 9917
rect 17037 9877 17049 9911
rect 17083 9908 17095 9911
rect 17126 9908 17132 9920
rect 17083 9880 17132 9908
rect 17083 9877 17095 9880
rect 17037 9871 17095 9877
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 19352 9908 19380 9948
rect 22278 9936 22284 9948
rect 22336 9936 22342 9988
rect 22388 9976 22416 10016
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 23017 9979 23075 9985
rect 23017 9976 23029 9979
rect 22388 9948 23029 9976
rect 23017 9945 23029 9948
rect 23063 9945 23075 9979
rect 23017 9939 23075 9945
rect 17276 9880 19380 9908
rect 17276 9868 17282 9880
rect 20438 9868 20444 9920
rect 20496 9908 20502 9920
rect 20625 9911 20683 9917
rect 20625 9908 20637 9911
rect 20496 9880 20637 9908
rect 20496 9868 20502 9880
rect 20625 9877 20637 9880
rect 20671 9908 20683 9911
rect 22002 9908 22008 9920
rect 20671 9880 22008 9908
rect 20671 9877 20683 9880
rect 20625 9871 20683 9877
rect 22002 9868 22008 9880
rect 22060 9868 22066 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22189 9911 22247 9917
rect 22189 9908 22201 9911
rect 22152 9880 22201 9908
rect 22152 9868 22158 9880
rect 22189 9877 22201 9880
rect 22235 9877 22247 9911
rect 22189 9871 22247 9877
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 22557 9911 22615 9917
rect 22557 9908 22569 9911
rect 22428 9880 22569 9908
rect 22428 9868 22434 9880
rect 22557 9877 22569 9880
rect 22603 9908 22615 9911
rect 23474 9908 23480 9920
rect 22603 9880 23480 9908
rect 22603 9877 22615 9880
rect 22557 9871 22615 9877
rect 23474 9868 23480 9880
rect 23532 9868 23538 9920
rect 1104 9818 23460 9840
rect 1104 9766 6548 9818
rect 6600 9766 6612 9818
rect 6664 9766 6676 9818
rect 6728 9766 6740 9818
rect 6792 9766 6804 9818
rect 6856 9766 12146 9818
rect 12198 9766 12210 9818
rect 12262 9766 12274 9818
rect 12326 9766 12338 9818
rect 12390 9766 12402 9818
rect 12454 9766 17744 9818
rect 17796 9766 17808 9818
rect 17860 9766 17872 9818
rect 17924 9766 17936 9818
rect 17988 9766 18000 9818
rect 18052 9766 23460 9818
rect 1104 9744 23460 9766
rect 3510 9704 3516 9716
rect 3471 9676 3516 9704
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 3786 9704 3792 9716
rect 3747 9676 3792 9704
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 6825 9707 6883 9713
rect 6825 9673 6837 9707
rect 6871 9704 6883 9707
rect 6914 9704 6920 9716
rect 6871 9676 6920 9704
rect 6871 9673 6883 9676
rect 6825 9667 6883 9673
rect 6914 9664 6920 9676
rect 6972 9704 6978 9716
rect 7926 9704 7932 9716
rect 6972 9676 7932 9704
rect 6972 9664 6978 9676
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 9861 9707 9919 9713
rect 9861 9673 9873 9707
rect 9907 9704 9919 9707
rect 10502 9704 10508 9716
rect 9907 9676 10508 9704
rect 9907 9673 9919 9676
rect 9861 9667 9919 9673
rect 5077 9639 5135 9645
rect 5077 9605 5089 9639
rect 5123 9636 5135 9639
rect 7282 9636 7288 9648
rect 5123 9608 7288 9636
rect 5123 9605 5135 9608
rect 5077 9599 5135 9605
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 9410 9639 9468 9645
rect 9410 9636 9422 9639
rect 7432 9608 9422 9636
rect 7432 9596 7438 9608
rect 9410 9605 9422 9608
rect 9456 9605 9468 9639
rect 9410 9599 9468 9605
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9568 1458 9580
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1452 9540 1685 9568
rect 1452 9528 1458 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 3326 9568 3332 9580
rect 3287 9540 3332 9568
rect 1673 9531 1731 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3602 9568 3608 9580
rect 3563 9540 3608 9568
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4522 9568 4528 9580
rect 4387 9540 4528 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 4264 9432 4292 9531
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 6178 9568 6184 9580
rect 5215 9540 6184 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 6638 9528 6644 9580
rect 6696 9568 6702 9580
rect 7938 9571 7996 9577
rect 7938 9568 7950 9571
rect 6696 9540 7950 9568
rect 6696 9528 6702 9540
rect 7938 9537 7950 9540
rect 7984 9568 7996 9571
rect 9677 9571 9735 9577
rect 7984 9540 8340 9568
rect 7984 9537 7996 9540
rect 7938 9531 7996 9537
rect 4430 9500 4436 9512
rect 4391 9472 4436 9500
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 5350 9500 5356 9512
rect 5311 9472 5356 9500
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 6270 9432 6276 9444
rect 4264 9404 6276 9432
rect 6270 9392 6276 9404
rect 6328 9392 6334 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 3881 9367 3939 9373
rect 3881 9364 3893 9367
rect 3200 9336 3893 9364
rect 3200 9324 3206 9336
rect 3881 9333 3893 9336
rect 3927 9333 3939 9367
rect 3881 9327 3939 9333
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 4709 9367 4767 9373
rect 4709 9364 4721 9367
rect 4488 9336 4721 9364
rect 4488 9324 4494 9336
rect 4709 9333 4721 9336
rect 4755 9333 4767 9367
rect 4709 9327 4767 9333
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 6512 9336 6653 9364
rect 6512 9324 6518 9336
rect 6641 9333 6653 9336
rect 6687 9364 6699 9367
rect 8220 9364 8248 9463
rect 8312 9441 8340 9540
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 9876 9568 9904 9667
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 11701 9707 11759 9713
rect 11701 9673 11713 9707
rect 11747 9704 11759 9707
rect 11790 9704 11796 9716
rect 11747 9676 11796 9704
rect 11747 9673 11759 9676
rect 11701 9667 11759 9673
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 13262 9704 13268 9716
rect 13223 9676 13268 9704
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13412 9676 13461 9704
rect 13412 9664 13418 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 16393 9707 16451 9713
rect 16393 9704 16405 9707
rect 15712 9676 16405 9704
rect 15712 9664 15718 9676
rect 16393 9673 16405 9676
rect 16439 9704 16451 9707
rect 16669 9707 16727 9713
rect 16669 9704 16681 9707
rect 16439 9676 16681 9704
rect 16439 9673 16451 9676
rect 16393 9667 16451 9673
rect 16669 9673 16681 9676
rect 16715 9673 16727 9707
rect 16669 9667 16727 9673
rect 11609 9639 11667 9645
rect 11609 9605 11621 9639
rect 11655 9636 11667 9639
rect 13280 9636 13308 9664
rect 15672 9636 15700 9664
rect 11655 9608 13308 9636
rect 11655 9605 11667 9608
rect 11609 9599 11667 9605
rect 10594 9568 10600 9580
rect 9723 9540 9904 9568
rect 10555 9540 10600 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 12825 9571 12883 9577
rect 12825 9537 12837 9571
rect 12871 9568 12883 9571
rect 13081 9571 13139 9577
rect 12871 9540 13032 9568
rect 12871 9537 12883 9540
rect 12825 9531 12883 9537
rect 10686 9500 10692 9512
rect 10647 9472 10692 9500
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9500 10931 9503
rect 10919 9472 11192 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 8297 9435 8355 9441
rect 8297 9401 8309 9435
rect 8343 9401 8355 9435
rect 8297 9395 8355 9401
rect 6687 9336 8248 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 11164 9373 11192 9472
rect 11256 9432 11284 9531
rect 13004 9500 13032 9540
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13280 9568 13308 9608
rect 14936 9608 15700 9636
rect 16684 9636 16712 9667
rect 17034 9664 17040 9716
rect 17092 9704 17098 9716
rect 19334 9704 19340 9716
rect 17092 9676 19340 9704
rect 17092 9664 17098 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 21266 9704 21272 9716
rect 19536 9676 21272 9704
rect 16684 9608 18828 9636
rect 13127 9540 13308 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 14936 9577 14964 9608
rect 14562 9571 14620 9577
rect 14562 9568 14574 9571
rect 13504 9540 14574 9568
rect 13504 9528 13510 9540
rect 14562 9537 14574 9540
rect 14608 9537 14620 9571
rect 14562 9531 14620 9537
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14875 9540 14933 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 15188 9571 15246 9577
rect 15188 9537 15200 9571
rect 15234 9568 15246 9571
rect 15470 9568 15476 9580
rect 15234 9540 15476 9568
rect 15234 9537 15246 9540
rect 15188 9531 15246 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9568 16911 9571
rect 17034 9568 17040 9580
rect 16899 9540 17040 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9568 17187 9571
rect 17494 9568 17500 9580
rect 17175 9540 17500 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 17494 9528 17500 9540
rect 17552 9568 17558 9580
rect 17770 9568 17776 9580
rect 17552 9540 17776 9568
rect 17552 9528 17558 9540
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18800 9577 18828 9608
rect 18966 9596 18972 9648
rect 19024 9636 19030 9648
rect 19150 9636 19156 9648
rect 19024 9608 19156 9636
rect 19024 9596 19030 9608
rect 19150 9596 19156 9608
rect 19208 9636 19214 9648
rect 19536 9636 19564 9676
rect 21266 9664 21272 9676
rect 21324 9664 21330 9716
rect 19208 9608 19564 9636
rect 19208 9596 19214 9608
rect 19610 9596 19616 9648
rect 19668 9636 19674 9648
rect 22094 9636 22100 9648
rect 19668 9608 20208 9636
rect 19668 9596 19674 9608
rect 18529 9571 18587 9577
rect 18529 9537 18541 9571
rect 18575 9568 18587 9571
rect 18785 9571 18843 9577
rect 18575 9540 18736 9568
rect 18575 9537 18587 9540
rect 18529 9531 18587 9537
rect 13354 9500 13360 9512
rect 13004 9472 13360 9500
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 17218 9500 17224 9512
rect 16316 9472 17224 9500
rect 16316 9441 16344 9472
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 18708 9500 18736 9540
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 19628 9568 19656 9596
rect 19978 9568 19984 9580
rect 20036 9577 20042 9580
rect 18831 9540 19656 9568
rect 19948 9540 19984 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 19978 9528 19984 9540
rect 20036 9531 20048 9577
rect 20036 9528 20042 9531
rect 18966 9500 18972 9512
rect 18708 9472 18972 9500
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 20180 9500 20208 9608
rect 22066 9596 22100 9636
rect 22152 9596 22158 9648
rect 22830 9636 22836 9648
rect 22791 9608 22836 9636
rect 22830 9596 22836 9608
rect 22888 9596 22894 9648
rect 20346 9568 20352 9580
rect 20307 9540 20352 9568
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 22066 9568 22094 9596
rect 21499 9540 22094 9568
rect 22189 9571 22247 9577
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 20180 9472 20269 9500
rect 20257 9469 20269 9472
rect 20303 9500 20315 9503
rect 20717 9503 20775 9509
rect 20717 9500 20729 9503
rect 20303 9472 20729 9500
rect 20303 9469 20315 9472
rect 20257 9463 20315 9469
rect 20717 9469 20729 9472
rect 20763 9500 20775 9503
rect 21082 9500 21088 9512
rect 20763 9472 21088 9500
rect 20763 9469 20775 9472
rect 20717 9463 20775 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21910 9500 21916 9512
rect 21871 9472 21916 9500
rect 21910 9460 21916 9472
rect 21968 9460 21974 9512
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 16301 9435 16359 9441
rect 11256 9404 11836 9432
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 9088 9336 10241 9364
rect 9088 9324 9094 9336
rect 10229 9333 10241 9336
rect 10275 9333 10287 9367
rect 10229 9327 10287 9333
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11330 9364 11336 9376
rect 11195 9336 11336 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11808 9364 11836 9404
rect 16301 9401 16313 9435
rect 16347 9401 16359 9435
rect 16301 9395 16359 9401
rect 17037 9435 17095 9441
rect 17037 9401 17049 9435
rect 17083 9432 17095 9435
rect 21637 9435 21695 9441
rect 17083 9404 17908 9432
rect 17083 9401 17095 9404
rect 17037 9395 17095 9401
rect 13538 9364 13544 9376
rect 11808 9336 13544 9364
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17405 9367 17463 9373
rect 17405 9333 17417 9367
rect 17451 9364 17463 9367
rect 17770 9364 17776 9376
rect 17451 9336 17776 9364
rect 17451 9333 17463 9336
rect 17405 9327 17463 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 17880 9364 17908 9404
rect 18800 9404 19380 9432
rect 18800 9364 18828 9404
rect 19352 9376 19380 9404
rect 21637 9401 21649 9435
rect 21683 9432 21695 9435
rect 22112 9432 22140 9463
rect 21683 9404 22140 9432
rect 21683 9401 21695 9404
rect 21637 9395 21695 9401
rect 17880 9336 18828 9364
rect 18877 9367 18935 9373
rect 18877 9333 18889 9367
rect 18923 9364 18935 9367
rect 18966 9364 18972 9376
rect 18923 9336 18972 9364
rect 18923 9333 18935 9336
rect 18877 9327 18935 9333
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 19334 9324 19340 9376
rect 19392 9324 19398 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 22204 9364 22232 9531
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 22649 9503 22707 9509
rect 22649 9500 22661 9503
rect 22336 9472 22661 9500
rect 22336 9460 22342 9472
rect 22649 9469 22661 9472
rect 22695 9469 22707 9503
rect 22649 9463 22707 9469
rect 20312 9336 22232 9364
rect 22557 9367 22615 9373
rect 20312 9324 20318 9336
rect 22557 9333 22569 9367
rect 22603 9364 22615 9367
rect 22646 9364 22652 9376
rect 22603 9336 22652 9364
rect 22603 9333 22615 9336
rect 22557 9327 22615 9333
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23014 9364 23020 9376
rect 22975 9336 23020 9364
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 1104 9274 23460 9296
rect 1104 9222 3749 9274
rect 3801 9222 3813 9274
rect 3865 9222 3877 9274
rect 3929 9222 3941 9274
rect 3993 9222 4005 9274
rect 4057 9222 9347 9274
rect 9399 9222 9411 9274
rect 9463 9222 9475 9274
rect 9527 9222 9539 9274
rect 9591 9222 9603 9274
rect 9655 9222 14945 9274
rect 14997 9222 15009 9274
rect 15061 9222 15073 9274
rect 15125 9222 15137 9274
rect 15189 9222 15201 9274
rect 15253 9222 20543 9274
rect 20595 9222 20607 9274
rect 20659 9222 20671 9274
rect 20723 9222 20735 9274
rect 20787 9222 20799 9274
rect 20851 9222 23460 9274
rect 1104 9200 23460 9222
rect 3602 9160 3608 9172
rect 3563 9132 3608 9160
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 5350 9160 5356 9172
rect 4396 9132 5356 9160
rect 4396 9120 4402 9132
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 6270 9160 6276 9172
rect 6231 9132 6276 9160
rect 6270 9120 6276 9132
rect 6328 9120 6334 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 10928 9132 12909 9160
rect 10928 9120 10934 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 13814 9160 13820 9172
rect 13775 9132 13820 9160
rect 12897 9123 12955 9129
rect 13814 9120 13820 9132
rect 13872 9160 13878 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 13872 9132 14197 9160
rect 13872 9120 13878 9132
rect 14185 9129 14197 9132
rect 14231 9160 14243 9163
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 14231 9132 14381 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16206 9160 16212 9172
rect 15979 9132 16212 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 3973 9095 4031 9101
rect 3973 9092 3985 9095
rect 3384 9064 3985 9092
rect 3384 9052 3390 9064
rect 3973 9061 3985 9064
rect 4019 9061 4031 9095
rect 3973 9055 4031 9061
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 6638 9092 6644 9104
rect 4212 9064 4660 9092
rect 4212 9052 4218 9064
rect 4632 9036 4660 9064
rect 5276 9064 6644 9092
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 8993 3019 9027
rect 3142 9024 3148 9036
rect 3103 8996 3148 9024
rect 2961 8987 3019 8993
rect 2976 8956 3004 8987
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 4430 9024 4436 9036
rect 4391 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 5276 9033 5304 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 13832 9092 13860 9120
rect 12820 9064 13860 9092
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 8993 5319 9027
rect 5261 8987 5319 8993
rect 5350 8984 5356 9036
rect 5408 9024 5414 9036
rect 12820 9033 12848 9064
rect 12805 9027 12863 9033
rect 5408 8996 5453 9024
rect 5408 8984 5414 8996
rect 12805 8993 12817 9027
rect 12851 8993 12863 9027
rect 13538 9024 13544 9036
rect 13499 8996 13544 9024
rect 12805 8987 12863 8993
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 14384 9024 14412 9123
rect 16206 9120 16212 9132
rect 16264 9160 16270 9172
rect 16264 9132 18552 9160
rect 16264 9120 16270 9132
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 14384 8996 14565 9024
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 18524 9024 18552 9132
rect 18598 9120 18604 9172
rect 18656 9160 18662 9172
rect 20254 9160 20260 9172
rect 18656 9132 20260 9160
rect 18656 9120 18662 9132
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20622 9120 20628 9172
rect 20680 9160 20686 9172
rect 22094 9160 22100 9172
rect 20680 9132 22100 9160
rect 20680 9120 20686 9132
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 19058 9092 19064 9104
rect 19019 9064 19064 9092
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 22189 9095 22247 9101
rect 22189 9061 22201 9095
rect 22235 9092 22247 9095
rect 23198 9092 23204 9104
rect 22235 9064 23204 9092
rect 22235 9061 22247 9064
rect 22189 9055 22247 9061
rect 23198 9052 23204 9064
rect 23256 9052 23262 9104
rect 19426 9024 19432 9036
rect 18524 8996 19432 9024
rect 14553 8987 14611 8993
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 22646 9024 22652 9036
rect 22607 8996 22652 9024
rect 22646 8984 22652 8996
rect 22704 8984 22710 9036
rect 22738 8984 22744 9036
rect 22796 9024 22802 9036
rect 22796 8996 22841 9024
rect 22796 8984 22802 8996
rect 4154 8956 4160 8968
rect 2976 8928 4160 8956
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 5074 8956 5080 8968
rect 4387 8928 5080 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 6914 8956 6920 8968
rect 5215 8928 6920 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 7699 8928 7880 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 4522 8848 4528 8900
rect 4580 8888 4586 8900
rect 5718 8888 5724 8900
rect 4580 8860 5724 8888
rect 4580 8848 4586 8860
rect 5718 8848 5724 8860
rect 5776 8888 5782 8900
rect 7386 8891 7444 8897
rect 7386 8888 7398 8891
rect 5776 8860 7398 8888
rect 5776 8848 5782 8860
rect 7386 8857 7398 8860
rect 7432 8857 7444 8891
rect 7386 8851 7444 8857
rect 3234 8820 3240 8832
rect 3195 8792 3240 8820
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4488 8792 4813 8820
rect 4488 8780 4494 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 4801 8783 4859 8789
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 7282 8820 7288 8832
rect 4948 8792 7288 8820
rect 4948 8780 4954 8792
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7852 8829 7880 8928
rect 8266 8928 8401 8956
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8820 7895 8823
rect 8266 8820 8294 8928
rect 8389 8925 8401 8928
rect 8435 8956 8447 8959
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 8435 8928 8585 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8573 8925 8585 8928
rect 8619 8956 8631 8959
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 8619 8928 9965 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 9953 8925 9965 8928
rect 9999 8956 10011 8959
rect 10042 8956 10048 8968
rect 9999 8928 10048 8956
rect 9999 8925 10011 8928
rect 9953 8919 10011 8925
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 10220 8959 10278 8965
rect 10220 8925 10232 8959
rect 10266 8956 10278 8959
rect 10594 8956 10600 8968
rect 10266 8928 10600 8956
rect 10266 8925 10278 8928
rect 10220 8919 10278 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 14826 8965 14832 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 12728 8928 13369 8956
rect 12560 8891 12618 8897
rect 12560 8888 12572 8891
rect 11348 8860 12572 8888
rect 11348 8829 11376 8860
rect 12560 8857 12572 8860
rect 12606 8888 12618 8891
rect 12728 8888 12756 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 14820 8956 14832 8965
rect 14787 8928 14832 8956
rect 13357 8919 13415 8925
rect 14820 8919 14832 8928
rect 14826 8916 14832 8919
rect 14884 8916 14890 8968
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8956 17463 8959
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17451 8928 17509 8956
rect 17451 8925 17463 8928
rect 17405 8919 17463 8925
rect 17497 8925 17509 8928
rect 17543 8956 17555 8959
rect 18138 8956 18144 8968
rect 17543 8928 18144 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 20358 8959 20416 8965
rect 20358 8925 20370 8959
rect 20404 8925 20416 8959
rect 20358 8919 20416 8925
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8956 20683 8959
rect 21082 8956 21088 8968
rect 20671 8928 21088 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 12606 8860 12756 8888
rect 12820 8860 13277 8888
rect 12606 8857 12618 8860
rect 12560 8851 12618 8857
rect 7883 8792 8294 8820
rect 11333 8823 11391 8829
rect 7883 8789 7895 8792
rect 7837 8783 7895 8789
rect 11333 8789 11345 8823
rect 11379 8789 11391 8823
rect 11333 8783 11391 8789
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 12820 8820 12848 8860
rect 13265 8857 13277 8860
rect 13311 8857 13323 8891
rect 13265 8851 13323 8857
rect 17160 8891 17218 8897
rect 17160 8857 17172 8891
rect 17206 8888 17218 8891
rect 17764 8891 17822 8897
rect 17206 8860 17724 8888
rect 17206 8857 17218 8860
rect 17160 8851 17218 8857
rect 11480 8792 12848 8820
rect 16025 8823 16083 8829
rect 11480 8780 11486 8792
rect 16025 8789 16037 8823
rect 16071 8820 16083 8823
rect 16114 8820 16120 8832
rect 16071 8792 16120 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 17696 8820 17724 8860
rect 17764 8857 17776 8891
rect 17810 8888 17822 8891
rect 17954 8888 17960 8900
rect 17810 8860 17960 8888
rect 17810 8857 17822 8860
rect 17764 8851 17822 8857
rect 17954 8848 17960 8860
rect 18012 8888 18018 8900
rect 18322 8888 18328 8900
rect 18012 8860 18328 8888
rect 18012 8848 18018 8860
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 20254 8888 20260 8900
rect 18892 8860 20260 8888
rect 18230 8820 18236 8832
rect 17696 8792 18236 8820
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 18892 8829 18920 8860
rect 20254 8848 20260 8860
rect 20312 8848 20318 8900
rect 20364 8888 20392 8919
rect 21082 8916 21088 8928
rect 21140 8956 21146 8968
rect 22097 8959 22155 8965
rect 22097 8956 22109 8959
rect 21140 8928 22109 8956
rect 21140 8916 21146 8928
rect 22097 8925 22109 8928
rect 22143 8956 22155 8959
rect 23014 8956 23020 8968
rect 22143 8928 23020 8956
rect 22143 8925 22155 8928
rect 22097 8919 22155 8925
rect 23014 8916 23020 8928
rect 23072 8916 23078 8968
rect 20438 8888 20444 8900
rect 20364 8860 20444 8888
rect 20438 8848 20444 8860
rect 20496 8848 20502 8900
rect 20530 8848 20536 8900
rect 20588 8888 20594 8900
rect 20588 8860 20760 8888
rect 20588 8848 20594 8860
rect 18877 8823 18935 8829
rect 18877 8789 18889 8823
rect 18923 8789 18935 8823
rect 18877 8783 18935 8789
rect 19245 8823 19303 8829
rect 19245 8789 19257 8823
rect 19291 8820 19303 8823
rect 19794 8820 19800 8832
rect 19291 8792 19800 8820
rect 19291 8789 19303 8792
rect 19245 8783 19303 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 20622 8820 20628 8832
rect 19944 8792 20628 8820
rect 19944 8780 19950 8792
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20732 8829 20760 8860
rect 21818 8848 21824 8900
rect 21876 8897 21882 8900
rect 21876 8888 21888 8897
rect 22554 8888 22560 8900
rect 21876 8860 21921 8888
rect 22515 8860 22560 8888
rect 21876 8851 21888 8860
rect 21876 8848 21882 8851
rect 22554 8848 22560 8860
rect 22612 8848 22618 8900
rect 20717 8823 20775 8829
rect 20717 8789 20729 8823
rect 20763 8789 20775 8823
rect 23014 8820 23020 8832
rect 22975 8792 23020 8820
rect 20717 8783 20775 8789
rect 23014 8780 23020 8792
rect 23072 8780 23078 8832
rect 1104 8730 23460 8752
rect 1104 8678 6548 8730
rect 6600 8678 6612 8730
rect 6664 8678 6676 8730
rect 6728 8678 6740 8730
rect 6792 8678 6804 8730
rect 6856 8678 12146 8730
rect 12198 8678 12210 8730
rect 12262 8678 12274 8730
rect 12326 8678 12338 8730
rect 12390 8678 12402 8730
rect 12454 8678 17744 8730
rect 17796 8678 17808 8730
rect 17860 8678 17872 8730
rect 17924 8678 17936 8730
rect 17988 8678 18000 8730
rect 18052 8678 23460 8730
rect 1104 8656 23460 8678
rect 3513 8619 3571 8625
rect 3513 8585 3525 8619
rect 3559 8616 3571 8619
rect 3694 8616 3700 8628
rect 3559 8588 3700 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 4890 8616 4896 8628
rect 3896 8588 4896 8616
rect 3145 8551 3203 8557
rect 3145 8517 3157 8551
rect 3191 8548 3203 8551
rect 3896 8548 3924 8588
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 6178 8616 6184 8628
rect 6139 8588 6184 8616
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 6972 8588 8309 8616
rect 6972 8576 6978 8588
rect 8297 8585 8309 8588
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10594 8616 10600 8628
rect 9999 8588 10600 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16758 8616 16764 8628
rect 16347 8588 16764 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18414 8616 18420 8628
rect 18095 8588 18420 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18414 8576 18420 8588
rect 18472 8616 18478 8628
rect 19150 8616 19156 8628
rect 18472 8588 19156 8616
rect 18472 8576 18478 8588
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19518 8616 19524 8628
rect 19479 8588 19524 8616
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20404 8588 23152 8616
rect 20404 8576 20410 8588
rect 3191 8520 3924 8548
rect 3973 8551 4031 8557
rect 3191 8517 3203 8520
rect 3145 8511 3203 8517
rect 3973 8517 3985 8551
rect 4019 8548 4031 8551
rect 4430 8548 4436 8560
rect 4019 8520 4436 8548
rect 4019 8517 4031 8520
rect 3973 8511 4031 8517
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 6454 8548 6460 8560
rect 4816 8520 6460 8548
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 4816 8489 4844 8520
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 8478 8548 8484 8560
rect 7024 8520 8484 8548
rect 4801 8483 4859 8489
rect 3660 8452 4384 8480
rect 3660 8440 3666 8452
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 3878 8412 3884 8424
rect 3099 8384 3884 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 2976 8344 3004 8375
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8381 4123 8415
rect 4065 8375 4123 8381
rect 2976 8316 3372 8344
rect 3344 8276 3372 8316
rect 3418 8304 3424 8356
rect 3476 8344 3482 8356
rect 3605 8347 3663 8353
rect 3605 8344 3617 8347
rect 3476 8316 3617 8344
rect 3476 8304 3482 8316
rect 3605 8313 3617 8316
rect 3651 8313 3663 8347
rect 3605 8307 3663 8313
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4080 8344 4108 8375
rect 4154 8372 4160 8424
rect 4212 8412 4218 8424
rect 4356 8412 4384 8452
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 5057 8483 5115 8489
rect 5057 8480 5069 8483
rect 4801 8443 4859 8449
rect 4908 8452 5069 8480
rect 4908 8412 4936 8452
rect 5057 8449 5069 8452
rect 5103 8449 5115 8483
rect 7024 8480 7052 8520
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 9861 8551 9919 8557
rect 9861 8548 9873 8551
rect 9692 8520 9873 8548
rect 9692 8492 9720 8520
rect 9861 8517 9873 8520
rect 9907 8548 9919 8551
rect 10042 8548 10048 8560
rect 9907 8520 10048 8548
rect 9907 8517 9919 8520
rect 9861 8511 9919 8517
rect 10042 8508 10048 8520
rect 10100 8548 10106 8560
rect 16925 8551 16983 8557
rect 16925 8548 16937 8551
rect 10100 8520 11376 8548
rect 10100 8508 10106 8520
rect 7098 8489 7104 8492
rect 5057 8443 5115 8449
rect 6380 8452 7052 8480
rect 4212 8384 4257 8412
rect 4356 8384 4936 8412
rect 4212 8372 4218 8384
rect 3752 8316 4108 8344
rect 3752 8304 3758 8316
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 6380 8344 6408 8452
rect 7092 8443 7104 8489
rect 7156 8480 7162 8492
rect 9410 8483 9468 8489
rect 9410 8480 9422 8483
rect 7156 8452 7192 8480
rect 8220 8452 9422 8480
rect 7098 8440 7104 8443
rect 7156 8440 7162 8452
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 4304 8316 4844 8344
rect 4304 8304 4310 8316
rect 4338 8276 4344 8288
rect 3344 8248 4344 8276
rect 4338 8236 4344 8248
rect 4396 8236 4402 8288
rect 4816 8276 4844 8316
rect 5736 8316 6408 8344
rect 6472 8384 6837 8412
rect 5736 8276 5764 8316
rect 6472 8288 6500 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 8220 8353 8248 8452
rect 9410 8449 9422 8452
rect 9456 8449 9468 8483
rect 9674 8480 9680 8492
rect 9587 8452 9680 8480
rect 9410 8443 9468 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 11348 8489 11376 8520
rect 16868 8520 16937 8548
rect 11066 8483 11124 8489
rect 11066 8480 11078 8483
rect 10744 8452 11078 8480
rect 10744 8440 10750 8452
rect 11066 8449 11078 8452
rect 11112 8480 11124 8483
rect 11333 8483 11391 8489
rect 11112 8452 11284 8480
rect 11112 8449 11124 8452
rect 11066 8443 11124 8449
rect 11256 8412 11284 8452
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 12630 8483 12688 8489
rect 12630 8480 12642 8483
rect 11572 8452 12642 8480
rect 11572 8440 11578 8452
rect 12630 8449 12642 8452
rect 12676 8449 12688 8483
rect 12630 8443 12688 8449
rect 14820 8483 14878 8489
rect 14820 8449 14832 8483
rect 14866 8480 14878 8483
rect 16114 8480 16120 8492
rect 14866 8452 16120 8480
rect 14866 8449 14878 8452
rect 14820 8443 14878 8449
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16868 8480 16896 8520
rect 16925 8517 16937 8520
rect 16971 8517 16983 8551
rect 16925 8511 16983 8517
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 22833 8551 22891 8557
rect 22833 8548 22845 8551
rect 17092 8520 22845 8548
rect 17092 8508 17098 8520
rect 22833 8517 22845 8520
rect 22879 8517 22891 8551
rect 22833 8511 22891 8517
rect 23124 8492 23152 8588
rect 16816 8452 16896 8480
rect 18408 8483 18466 8489
rect 16816 8440 16822 8452
rect 18408 8449 18420 8483
rect 18454 8480 18466 8483
rect 19242 8480 19248 8492
rect 18454 8452 19248 8480
rect 18454 8449 18466 8452
rect 18408 8443 18466 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19869 8483 19927 8489
rect 19869 8480 19881 8483
rect 19352 8452 19881 8480
rect 12897 8415 12955 8421
rect 11256 8384 11560 8412
rect 11532 8353 11560 8384
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 14553 8415 14611 8421
rect 12943 8384 13124 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 8205 8347 8263 8353
rect 8205 8344 8217 8347
rect 8168 8316 8217 8344
rect 8168 8304 8174 8316
rect 8205 8313 8217 8316
rect 8251 8313 8263 8347
rect 8205 8307 8263 8313
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 6454 8276 6460 8288
rect 4816 8248 5764 8276
rect 6415 8248 6460 8276
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 13096 8285 13124 8384
rect 14553 8381 14565 8415
rect 14599 8381 14611 8415
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 14553 8375 14611 8381
rect 16408 8384 16681 8412
rect 13081 8279 13139 8285
rect 13081 8245 13093 8279
rect 13127 8276 13139 8279
rect 13357 8279 13415 8285
rect 13357 8276 13369 8279
rect 13127 8248 13369 8276
rect 13127 8245 13139 8248
rect 13081 8239 13139 8245
rect 13357 8245 13369 8248
rect 13403 8276 13415 8279
rect 13541 8279 13599 8285
rect 13541 8276 13553 8279
rect 13403 8248 13553 8276
rect 13403 8245 13415 8248
rect 13357 8239 13415 8245
rect 13541 8245 13553 8248
rect 13587 8276 13599 8279
rect 13725 8279 13783 8285
rect 13725 8276 13737 8279
rect 13587 8248 13737 8276
rect 13587 8245 13599 8248
rect 13541 8239 13599 8245
rect 13725 8245 13737 8248
rect 13771 8276 13783 8279
rect 13909 8279 13967 8285
rect 13909 8276 13921 8279
rect 13771 8248 13921 8276
rect 13771 8245 13783 8248
rect 13725 8239 13783 8245
rect 13909 8245 13921 8248
rect 13955 8276 13967 8279
rect 14093 8279 14151 8285
rect 14093 8276 14105 8279
rect 13955 8248 14105 8276
rect 13955 8245 13967 8248
rect 13909 8239 13967 8245
rect 14093 8245 14105 8248
rect 14139 8276 14151 8279
rect 14277 8279 14335 8285
rect 14277 8276 14289 8279
rect 14139 8248 14289 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 14277 8245 14289 8248
rect 14323 8276 14335 8279
rect 14461 8279 14519 8285
rect 14461 8276 14473 8279
rect 14323 8248 14473 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 14461 8245 14473 8248
rect 14507 8276 14519 8279
rect 14568 8276 14596 8375
rect 15930 8344 15936 8356
rect 15891 8316 15936 8344
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 16408 8353 16436 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 18138 8412 18144 8424
rect 18051 8384 18144 8412
rect 16669 8375 16727 8381
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 19352 8412 19380 8452
rect 19869 8449 19881 8452
rect 19915 8449 19927 8483
rect 21174 8480 21180 8492
rect 21135 8452 21180 8480
rect 19869 8443 19927 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 21542 8480 21548 8492
rect 21407 8452 21548 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 22060 8452 22201 8480
rect 22060 8440 22066 8452
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 23106 8480 23112 8492
rect 23067 8452 23112 8480
rect 22189 8443 22247 8449
rect 23106 8440 23112 8452
rect 23164 8440 23170 8492
rect 19610 8412 19616 8424
rect 19208 8384 19380 8412
rect 19571 8384 19616 8412
rect 19208 8372 19214 8384
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 22278 8412 22284 8424
rect 22239 8384 22284 8412
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 22373 8415 22431 8421
rect 22373 8381 22385 8415
rect 22419 8381 22431 8415
rect 23566 8412 23572 8424
rect 22373 8375 22431 8381
rect 22480 8384 23572 8412
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 16040 8316 16129 8344
rect 16040 8276 16068 8316
rect 16117 8313 16129 8316
rect 16163 8344 16175 8347
rect 16393 8347 16451 8353
rect 16393 8344 16405 8347
rect 16163 8316 16405 8344
rect 16163 8313 16175 8316
rect 16117 8307 16175 8313
rect 16393 8313 16405 8316
rect 16439 8344 16451 8347
rect 16439 8316 16712 8344
rect 16439 8313 16451 8316
rect 16393 8307 16451 8313
rect 14507 8248 16068 8276
rect 16684 8276 16712 8316
rect 18156 8276 18184 8372
rect 20548 8316 21220 8344
rect 19610 8276 19616 8288
rect 16684 8248 19616 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 20254 8236 20260 8288
rect 20312 8276 20318 8288
rect 20548 8276 20576 8316
rect 20312 8248 20576 8276
rect 20312 8236 20318 8248
rect 20622 8236 20628 8288
rect 20680 8276 20686 8288
rect 20993 8279 21051 8285
rect 20993 8276 21005 8279
rect 20680 8248 21005 8276
rect 20680 8236 20686 8248
rect 20993 8245 21005 8248
rect 21039 8245 21051 8279
rect 21192 8276 21220 8316
rect 21266 8304 21272 8356
rect 21324 8344 21330 8356
rect 21545 8347 21603 8353
rect 21545 8344 21557 8347
rect 21324 8316 21557 8344
rect 21324 8304 21330 8316
rect 21545 8313 21557 8316
rect 21591 8313 21603 8347
rect 21818 8344 21824 8356
rect 21779 8316 21824 8344
rect 21545 8307 21603 8313
rect 21818 8304 21824 8316
rect 21876 8304 21882 8356
rect 22388 8344 22416 8375
rect 21928 8316 22416 8344
rect 21928 8276 21956 8316
rect 21192 8248 21956 8276
rect 20993 8239 21051 8245
rect 22094 8236 22100 8288
rect 22152 8276 22158 8288
rect 22480 8276 22508 8384
rect 23566 8372 23572 8384
rect 23624 8372 23630 8424
rect 22152 8248 22508 8276
rect 22152 8236 22158 8248
rect 1104 8186 23460 8208
rect 1104 8134 3749 8186
rect 3801 8134 3813 8186
rect 3865 8134 3877 8186
rect 3929 8134 3941 8186
rect 3993 8134 4005 8186
rect 4057 8134 9347 8186
rect 9399 8134 9411 8186
rect 9463 8134 9475 8186
rect 9527 8134 9539 8186
rect 9591 8134 9603 8186
rect 9655 8134 14945 8186
rect 14997 8134 15009 8186
rect 15061 8134 15073 8186
rect 15125 8134 15137 8186
rect 15189 8134 15201 8186
rect 15253 8134 20543 8186
rect 20595 8134 20607 8186
rect 20659 8134 20671 8186
rect 20723 8134 20735 8186
rect 20787 8134 20799 8186
rect 20851 8134 23460 8186
rect 1104 8112 23460 8134
rect 7374 8072 7380 8084
rect 7335 8044 7380 8072
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 20990 8072 20996 8084
rect 19628 8044 20996 8072
rect 18785 8007 18843 8013
rect 18785 7973 18797 8007
rect 18831 8004 18843 8007
rect 19518 8004 19524 8016
rect 18831 7976 19524 8004
rect 18831 7973 18843 7976
rect 18785 7967 18843 7973
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 9769 7939 9827 7945
rect 9769 7936 9781 7939
rect 9732 7908 9781 7936
rect 9732 7896 9738 7908
rect 9769 7905 9781 7908
rect 9815 7905 9827 7939
rect 9769 7899 9827 7905
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 11388 7908 11805 7936
rect 11388 7896 11394 7908
rect 11793 7905 11805 7908
rect 11839 7905 11851 7939
rect 19628 7936 19656 8044
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 21082 7964 21088 8016
rect 21140 8004 21146 8016
rect 21140 7976 21312 8004
rect 21140 7964 21146 7976
rect 21174 7936 21180 7948
rect 11793 7899 11851 7905
rect 18340 7908 19656 7936
rect 20548 7908 21180 7936
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 5534 7868 5540 7880
rect 4479 7840 5540 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 7331 7840 8769 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 8757 7837 8769 7840
rect 8803 7868 8815 7871
rect 9692 7868 9720 7896
rect 8803 7840 8984 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 4700 7803 4758 7809
rect 4700 7769 4712 7803
rect 4746 7800 4758 7803
rect 5350 7800 5356 7812
rect 4746 7772 5356 7800
rect 4746 7769 4758 7772
rect 4700 7763 4758 7769
rect 5350 7760 5356 7772
rect 5408 7800 5414 7812
rect 6914 7800 6920 7812
rect 5408 7772 6920 7800
rect 5408 7760 5414 7772
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 7040 7803 7098 7809
rect 7040 7769 7052 7803
rect 7086 7800 7098 7803
rect 7086 7772 8432 7800
rect 7086 7769 7098 7772
rect 7040 7763 7098 7769
rect 5718 7692 5724 7744
rect 5776 7732 5782 7744
rect 5813 7735 5871 7741
rect 5813 7732 5825 7735
rect 5776 7704 5825 7732
rect 5776 7692 5782 7704
rect 5813 7701 5825 7704
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 8404 7732 8432 7772
rect 8478 7760 8484 7812
rect 8536 7809 8542 7812
rect 8536 7800 8548 7809
rect 8536 7772 8581 7800
rect 8536 7763 8548 7772
rect 8536 7760 8542 7763
rect 8956 7744 8984 7840
rect 9600 7840 9720 7868
rect 10036 7871 10094 7877
rect 8662 7732 8668 7744
rect 5960 7704 6005 7732
rect 8404 7704 8668 7732
rect 5960 7692 5966 7704
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 8938 7732 8944 7744
rect 8899 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7732 9002 7744
rect 9600 7741 9628 7840
rect 10036 7837 10048 7871
rect 10082 7868 10094 7871
rect 11422 7868 11428 7880
rect 10082 7840 11428 7868
rect 10082 7837 10094 7840
rect 10036 7831 10094 7837
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7868 12219 7871
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 12207 7840 12357 7868
rect 12207 7837 12219 7840
rect 12161 7831 12219 7837
rect 12345 7837 12357 7840
rect 12391 7868 12403 7871
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12391 7840 12541 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 12529 7837 12541 7840
rect 12575 7868 12587 7871
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 12575 7840 14105 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 14093 7837 14105 7840
rect 14139 7868 14151 7871
rect 14642 7868 14648 7880
rect 14139 7840 14648 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7868 15623 7871
rect 16206 7868 16212 7880
rect 15611 7840 16212 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 18161 7871 18219 7877
rect 18161 7837 18173 7871
rect 18207 7868 18219 7871
rect 18340 7868 18368 7908
rect 18207 7840 18368 7868
rect 18417 7871 18475 7877
rect 18207 7837 18219 7840
rect 18161 7831 18219 7837
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 18601 7871 18659 7877
rect 18601 7837 18613 7871
rect 18647 7868 18659 7871
rect 18874 7868 18880 7880
rect 18647 7840 18880 7868
rect 18647 7837 18659 7840
rect 18601 7831 18659 7837
rect 12802 7809 12808 7812
rect 11701 7803 11759 7809
rect 11701 7800 11713 7803
rect 11164 7772 11713 7800
rect 11164 7744 11192 7772
rect 11701 7769 11713 7772
rect 11747 7769 11759 7803
rect 12796 7800 12808 7809
rect 12763 7772 12808 7800
rect 11701 7763 11759 7769
rect 12796 7763 12808 7772
rect 12802 7760 12808 7763
rect 12860 7760 12866 7812
rect 12894 7760 12900 7812
rect 12952 7800 12958 7812
rect 14338 7803 14396 7809
rect 14338 7800 14350 7803
rect 12952 7772 14350 7800
rect 12952 7760 12958 7772
rect 14338 7769 14350 7772
rect 14384 7769 14396 7803
rect 14338 7763 14396 7769
rect 15832 7803 15890 7809
rect 15832 7769 15844 7803
rect 15878 7800 15890 7803
rect 18432 7800 18460 7831
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19061 7871 19119 7877
rect 19061 7837 19073 7871
rect 19107 7868 19119 7871
rect 20548 7868 20576 7908
rect 21174 7896 21180 7908
rect 21232 7896 21238 7948
rect 21284 7945 21312 7976
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7905 21327 7939
rect 21726 7936 21732 7948
rect 21690 7908 21732 7936
rect 21269 7899 21327 7905
rect 21726 7896 21732 7908
rect 21784 7896 21790 7948
rect 19107 7840 20576 7868
rect 20625 7871 20683 7877
rect 19107 7837 19119 7840
rect 19061 7831 19119 7837
rect 20625 7837 20637 7871
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 15878 7772 18092 7800
rect 18432 7772 19656 7800
rect 15878 7769 15890 7772
rect 15832 7763 15890 7769
rect 18064 7744 18092 7772
rect 19628 7744 19656 7772
rect 20254 7760 20260 7812
rect 20312 7800 20318 7812
rect 20358 7803 20416 7809
rect 20358 7800 20370 7803
rect 20312 7772 20370 7800
rect 20312 7760 20318 7772
rect 20358 7769 20370 7772
rect 20404 7769 20416 7803
rect 20358 7763 20416 7769
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 8996 7704 9137 7732
rect 8996 7692 9002 7704
rect 9125 7701 9137 7704
rect 9171 7732 9183 7735
rect 9585 7735 9643 7741
rect 9585 7732 9597 7735
rect 9171 7704 9597 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9585 7701 9597 7704
rect 9631 7701 9643 7735
rect 11146 7732 11152 7744
rect 11107 7704 11152 7732
rect 9585 7695 9643 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 11609 7735 11667 7741
rect 11296 7704 11341 7732
rect 11296 7692 11302 7704
rect 11609 7701 11621 7735
rect 11655 7732 11667 7735
rect 12066 7732 12072 7744
rect 11655 7704 12072 7732
rect 11655 7701 11667 7704
rect 11609 7695 11667 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 13906 7732 13912 7744
rect 13867 7704 13912 7732
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 15473 7735 15531 7741
rect 15473 7701 15485 7735
rect 15519 7732 15531 7735
rect 16758 7732 16764 7744
rect 15519 7704 16764 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 16942 7732 16948 7744
rect 16903 7704 16948 7732
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 17092 7704 17137 7732
rect 17092 7692 17098 7704
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 18322 7692 18328 7744
rect 18380 7732 18386 7744
rect 18690 7732 18696 7744
rect 18380 7704 18696 7732
rect 18380 7692 18386 7704
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 19242 7732 19248 7744
rect 19203 7704 19248 7732
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 20640 7732 20668 7831
rect 21358 7828 21364 7880
rect 21416 7868 21422 7880
rect 21592 7871 21650 7877
rect 21592 7868 21604 7871
rect 21416 7840 21604 7868
rect 21416 7828 21422 7840
rect 21592 7837 21604 7840
rect 21638 7837 21650 7871
rect 21592 7831 21650 7837
rect 22005 7871 22063 7877
rect 22005 7837 22017 7871
rect 22051 7868 22063 7871
rect 22370 7868 22376 7880
rect 22051 7840 22376 7868
rect 22051 7837 22063 7840
rect 22005 7831 22063 7837
rect 22370 7828 22376 7840
rect 22428 7828 22434 7880
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 20864 7772 20913 7800
rect 20864 7760 20870 7772
rect 20901 7769 20913 7772
rect 20947 7769 20959 7803
rect 20901 7763 20959 7769
rect 21085 7803 21143 7809
rect 21085 7769 21097 7803
rect 21131 7769 21143 7803
rect 21085 7763 21143 7769
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 19668 7704 20729 7732
rect 19668 7692 19674 7704
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 21100 7732 21128 7763
rect 22002 7732 22008 7744
rect 21100 7704 22008 7732
rect 20717 7695 20775 7701
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 23106 7732 23112 7744
rect 23067 7704 23112 7732
rect 23106 7692 23112 7704
rect 23164 7692 23170 7744
rect 1104 7642 23460 7664
rect 1104 7590 6548 7642
rect 6600 7590 6612 7642
rect 6664 7590 6676 7642
rect 6728 7590 6740 7642
rect 6792 7590 6804 7642
rect 6856 7590 12146 7642
rect 12198 7590 12210 7642
rect 12262 7590 12274 7642
rect 12326 7590 12338 7642
rect 12390 7590 12402 7642
rect 12454 7590 17744 7642
rect 17796 7590 17808 7642
rect 17860 7590 17872 7642
rect 17924 7590 17936 7642
rect 17988 7590 18000 7642
rect 18052 7590 23460 7642
rect 1104 7568 23460 7590
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3292 7500 3985 7528
rect 3292 7488 3298 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 3973 7491 4031 7497
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 6178 7528 6184 7540
rect 4387 7500 6184 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 9732 7500 11345 7528
rect 9732 7488 9738 7500
rect 11333 7497 11345 7500
rect 11379 7528 11391 7531
rect 11422 7528 11428 7540
rect 11379 7500 11428 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 13081 7531 13139 7537
rect 13081 7497 13093 7531
rect 13127 7528 13139 7531
rect 13446 7528 13452 7540
rect 13127 7500 13452 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 17954 7528 17960 7540
rect 14516 7500 17960 7528
rect 14516 7488 14522 7500
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 18049 7531 18107 7537
rect 18049 7497 18061 7531
rect 18095 7528 18107 7531
rect 18230 7528 18236 7540
rect 18095 7500 18236 7528
rect 18095 7497 18107 7500
rect 18049 7491 18107 7497
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 21450 7528 21456 7540
rect 21411 7500 21456 7528
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 21634 7488 21640 7540
rect 21692 7488 21698 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 22152 7500 22197 7528
rect 22152 7488 22158 7500
rect 22278 7488 22284 7540
rect 22336 7528 22342 7540
rect 22557 7531 22615 7537
rect 22557 7528 22569 7531
rect 22336 7500 22569 7528
rect 22336 7488 22342 7500
rect 22557 7497 22569 7500
rect 22603 7497 22615 7531
rect 22557 7491 22615 7497
rect 5534 7460 5540 7472
rect 4816 7432 5540 7460
rect 4816 7401 4844 7432
rect 5534 7420 5540 7432
rect 5592 7460 5598 7472
rect 6454 7460 6460 7472
rect 5592 7432 6460 7460
rect 5592 7420 5598 7432
rect 6454 7420 6460 7432
rect 6512 7460 6518 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 6512 7432 6653 7460
rect 6512 7420 6518 7432
rect 6641 7429 6653 7432
rect 6687 7460 6699 7463
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 6687 7432 6837 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 6825 7429 6837 7432
rect 6871 7460 6883 7463
rect 8938 7460 8944 7472
rect 6871 7432 8944 7460
rect 6871 7429 6883 7432
rect 6825 7423 6883 7429
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4801 7395 4859 7401
rect 4479 7364 4752 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 4525 7327 4583 7333
rect 4525 7324 4537 7327
rect 4396 7296 4537 7324
rect 4396 7284 4402 7296
rect 4525 7293 4537 7296
rect 4571 7293 4583 7327
rect 4724 7324 4752 7364
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 5068 7395 5126 7401
rect 5068 7392 5080 7395
rect 4801 7355 4859 7361
rect 4908 7364 5080 7392
rect 4908 7324 4936 7364
rect 5068 7361 5080 7364
rect 5114 7392 5126 7395
rect 5626 7392 5632 7404
rect 5114 7364 5632 7392
rect 5114 7361 5126 7364
rect 5068 7355 5126 7361
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 6932 7401 6960 7432
rect 8496 7401 8524 7432
rect 8938 7420 8944 7432
rect 8996 7460 9002 7472
rect 9858 7460 9864 7472
rect 8996 7432 9864 7460
rect 8996 7420 9002 7432
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 14286 7463 14344 7469
rect 14286 7460 14298 7463
rect 13964 7432 14298 7460
rect 13964 7420 13970 7432
rect 14286 7429 14298 7432
rect 14332 7460 14344 7463
rect 14550 7460 14556 7472
rect 14332 7432 14556 7460
rect 14332 7429 14344 7432
rect 14286 7423 14344 7429
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 17034 7420 17040 7472
rect 17092 7420 17098 7472
rect 18782 7420 18788 7472
rect 18840 7460 18846 7472
rect 19254 7463 19312 7469
rect 19254 7460 19266 7463
rect 18840 7432 19266 7460
rect 18840 7420 18846 7432
rect 19254 7429 19266 7432
rect 19300 7429 19312 7463
rect 19254 7423 19312 7429
rect 19426 7420 19432 7472
rect 19484 7460 19490 7472
rect 19858 7463 19916 7469
rect 19858 7460 19870 7463
rect 19484 7432 19870 7460
rect 19484 7420 19490 7432
rect 19858 7429 19870 7432
rect 19904 7429 19916 7463
rect 19858 7423 19916 7429
rect 21269 7463 21327 7469
rect 21269 7429 21281 7463
rect 21315 7460 21327 7463
rect 21652 7460 21680 7488
rect 22830 7460 22836 7472
rect 21315 7432 21680 7460
rect 22791 7432 22836 7460
rect 21315 7429 21327 7432
rect 21269 7423 21327 7429
rect 22830 7420 22836 7432
rect 22888 7420 22894 7472
rect 8754 7401 8760 7404
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 7173 7395 7231 7401
rect 7173 7392 7185 7395
rect 6917 7355 6975 7361
rect 7024 7364 7185 7392
rect 4724 7296 4936 7324
rect 4525 7287 4583 7293
rect 5810 7284 5816 7336
rect 5868 7324 5874 7336
rect 7024 7324 7052 7364
rect 7173 7361 7185 7364
rect 7219 7361 7231 7395
rect 7173 7355 7231 7361
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7361 8539 7395
rect 8748 7392 8760 7401
rect 8715 7364 8760 7392
rect 8481 7355 8539 7361
rect 8748 7355 8760 7364
rect 8754 7352 8760 7355
rect 8812 7352 8818 7404
rect 9876 7392 9904 7420
rect 10226 7401 10232 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9876 7364 9965 7392
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 10220 7392 10232 7401
rect 10187 7364 10232 7392
rect 9953 7355 10011 7361
rect 10220 7355 10232 7364
rect 10226 7352 10232 7355
rect 10284 7352 10290 7404
rect 11609 7395 11667 7401
rect 11609 7361 11621 7395
rect 11655 7392 11667 7395
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11655 7364 11713 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 11701 7361 11713 7364
rect 11747 7392 11759 7395
rect 11790 7392 11796 7404
rect 11747 7364 11796 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 11974 7401 11980 7404
rect 11968 7355 11980 7401
rect 12032 7392 12038 7404
rect 15769 7395 15827 7401
rect 12032 7364 12068 7392
rect 11974 7352 11980 7355
rect 12032 7352 12038 7364
rect 15769 7361 15781 7395
rect 15815 7392 15827 7395
rect 15930 7392 15936 7404
rect 15815 7364 15936 7392
rect 15815 7361 15827 7364
rect 15769 7355 15827 7361
rect 15930 7352 15936 7364
rect 15988 7352 15994 7404
rect 16936 7395 16994 7401
rect 16936 7361 16948 7395
rect 16982 7392 16994 7395
rect 17052 7392 17080 7420
rect 18874 7392 18880 7404
rect 16982 7364 18880 7392
rect 16982 7361 16994 7364
rect 16936 7355 16994 7361
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 21637 7395 21695 7401
rect 21637 7361 21649 7395
rect 21683 7361 21695 7395
rect 21637 7355 21695 7361
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22278 7392 22284 7404
rect 22235 7364 22284 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 5868 7296 7052 7324
rect 14553 7327 14611 7333
rect 5868 7284 5874 7296
rect 14553 7293 14565 7327
rect 14599 7324 14611 7327
rect 14642 7324 14648 7336
rect 14599 7296 14648 7324
rect 14599 7293 14611 7296
rect 14553 7287 14611 7293
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 16025 7327 16083 7333
rect 16025 7293 16037 7327
rect 16071 7324 16083 7327
rect 16669 7327 16727 7333
rect 16071 7296 16252 7324
rect 16071 7293 16083 7296
rect 16025 7287 16083 7293
rect 16224 7200 16252 7296
rect 16669 7293 16681 7327
rect 16715 7293 16727 7327
rect 16669 7287 16727 7293
rect 19521 7327 19579 7333
rect 19521 7293 19533 7327
rect 19567 7324 19579 7327
rect 19610 7324 19616 7336
rect 19567 7296 19616 7324
rect 19567 7293 19579 7296
rect 19521 7287 19579 7293
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8754 7188 8760 7200
rect 8343 7160 8760 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8754 7148 8760 7160
rect 8812 7148 8818 7200
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13228 7160 13273 7188
rect 13228 7148 13234 7160
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 14645 7191 14703 7197
rect 14645 7188 14657 7191
rect 14332 7160 14657 7188
rect 14332 7148 14338 7160
rect 14645 7157 14657 7160
rect 14691 7157 14703 7191
rect 16206 7188 16212 7200
rect 16119 7160 16212 7188
rect 14645 7151 14703 7157
rect 16206 7148 16212 7160
rect 16264 7188 16270 7200
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 16264 7160 16405 7188
rect 16264 7148 16270 7160
rect 16393 7157 16405 7160
rect 16439 7188 16451 7191
rect 16684 7188 16712 7287
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 18138 7256 18144 7268
rect 18099 7228 18144 7256
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 21652 7256 21680 7355
rect 22278 7352 22284 7364
rect 22336 7392 22342 7404
rect 22922 7392 22928 7404
rect 22336 7364 22928 7392
rect 22336 7352 22342 7364
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 21818 7284 21824 7336
rect 21876 7324 21882 7336
rect 21913 7327 21971 7333
rect 21913 7324 21925 7327
rect 21876 7296 21925 7324
rect 21876 7284 21882 7296
rect 21913 7293 21925 7296
rect 21959 7293 21971 7327
rect 21913 7287 21971 7293
rect 22094 7256 22100 7268
rect 20548 7228 21588 7256
rect 21652 7228 22100 7256
rect 17586 7188 17592 7200
rect 16439 7160 17592 7188
rect 16439 7157 16451 7160
rect 16393 7151 16451 7157
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 20548 7188 20576 7228
rect 19208 7160 20576 7188
rect 20993 7191 21051 7197
rect 19208 7148 19214 7160
rect 20993 7157 21005 7191
rect 21039 7188 21051 7191
rect 21450 7188 21456 7200
rect 21039 7160 21456 7188
rect 21039 7157 21051 7160
rect 20993 7151 21051 7157
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 21560 7188 21588 7228
rect 22094 7216 22100 7228
rect 22152 7216 22158 7268
rect 22646 7256 22652 7268
rect 22607 7228 22652 7256
rect 22646 7216 22652 7228
rect 22704 7216 22710 7268
rect 22370 7188 22376 7200
rect 21560 7160 22376 7188
rect 22370 7148 22376 7160
rect 22428 7188 22434 7200
rect 22830 7188 22836 7200
rect 22428 7160 22836 7188
rect 22428 7148 22434 7160
rect 22830 7148 22836 7160
rect 22888 7148 22894 7200
rect 23014 7188 23020 7200
rect 22975 7160 23020 7188
rect 23014 7148 23020 7160
rect 23072 7148 23078 7200
rect 1104 7098 23460 7120
rect 1104 7046 3749 7098
rect 3801 7046 3813 7098
rect 3865 7046 3877 7098
rect 3929 7046 3941 7098
rect 3993 7046 4005 7098
rect 4057 7046 9347 7098
rect 9399 7046 9411 7098
rect 9463 7046 9475 7098
rect 9527 7046 9539 7098
rect 9591 7046 9603 7098
rect 9655 7046 14945 7098
rect 14997 7046 15009 7098
rect 15061 7046 15073 7098
rect 15125 7046 15137 7098
rect 15189 7046 15201 7098
rect 15253 7046 20543 7098
rect 20595 7046 20607 7098
rect 20659 7046 20671 7098
rect 20723 7046 20735 7098
rect 20787 7046 20799 7098
rect 20851 7046 23460 7098
rect 1104 7024 23460 7046
rect 5626 6984 5632 6996
rect 5587 6956 5632 6984
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 8478 6984 8484 6996
rect 8439 6956 8484 6984
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 12124 6956 12173 6984
rect 12124 6944 12130 6956
rect 12161 6953 12173 6956
rect 12207 6953 12219 6987
rect 12618 6984 12624 6996
rect 12161 6947 12219 6953
rect 12268 6956 12624 6984
rect 11790 6876 11796 6928
rect 11848 6916 11854 6928
rect 12268 6916 12296 6956
rect 12618 6944 12624 6956
rect 12676 6984 12682 6996
rect 13817 6987 13875 6993
rect 13817 6984 13829 6987
rect 12676 6956 13829 6984
rect 12676 6944 12682 6956
rect 13817 6953 13829 6956
rect 13863 6984 13875 6987
rect 13906 6984 13912 6996
rect 13863 6956 13912 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 13906 6944 13912 6956
rect 13964 6984 13970 6996
rect 14185 6987 14243 6993
rect 14185 6984 14197 6987
rect 13964 6956 14197 6984
rect 13964 6944 13970 6956
rect 14185 6953 14197 6956
rect 14231 6984 14243 6987
rect 14369 6987 14427 6993
rect 14369 6984 14381 6987
rect 14231 6956 14381 6984
rect 14231 6953 14243 6956
rect 14185 6947 14243 6953
rect 14369 6953 14381 6956
rect 14415 6984 14427 6987
rect 14642 6984 14648 6996
rect 14415 6956 14648 6984
rect 14415 6953 14427 6956
rect 14369 6947 14427 6953
rect 14642 6944 14648 6956
rect 14700 6984 14706 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 14700 6956 14749 6984
rect 14700 6944 14706 6956
rect 14737 6953 14749 6956
rect 14783 6984 14795 6987
rect 16206 6984 16212 6996
rect 14783 6956 16212 6984
rect 14783 6953 14795 6956
rect 14737 6947 14795 6953
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 18748 6956 19104 6984
rect 18748 6944 18754 6956
rect 19076 6925 19104 6956
rect 19242 6944 19248 6996
rect 19300 6984 19306 6996
rect 22370 6984 22376 6996
rect 19300 6956 22376 6984
rect 19300 6944 19306 6956
rect 22370 6944 22376 6956
rect 22428 6944 22434 6996
rect 23106 6944 23112 6996
rect 23164 6944 23170 6996
rect 19061 6919 19119 6925
rect 11848 6888 12296 6916
rect 11848 6876 11854 6888
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1636 6752 1961 6780
rect 1636 6740 1642 6752
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 6178 6740 6184 6792
rect 6236 6780 6242 6792
rect 7009 6783 7067 6789
rect 6236 6752 6868 6780
rect 6236 6740 6242 6752
rect 6270 6672 6276 6724
rect 6328 6712 6334 6724
rect 6742 6715 6800 6721
rect 6742 6712 6754 6715
rect 6328 6684 6754 6712
rect 6328 6672 6334 6684
rect 6742 6681 6754 6684
rect 6788 6681 6800 6715
rect 6840 6712 6868 6752
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 7055 6752 7113 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7101 6749 7113 6752
rect 7147 6780 7159 6783
rect 8386 6780 8392 6792
rect 7147 6752 8392 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 8386 6740 8392 6752
rect 8444 6780 8450 6792
rect 8665 6783 8723 6789
rect 8665 6780 8677 6783
rect 8444 6752 8677 6780
rect 8444 6740 8450 6752
rect 8665 6749 8677 6752
rect 8711 6780 8723 6783
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8711 6752 9045 6780
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 9033 6749 9045 6752
rect 9079 6780 9091 6783
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9079 6752 9321 6780
rect 9079 6749 9091 6752
rect 9033 6743 9091 6749
rect 9309 6749 9321 6752
rect 9355 6780 9367 6783
rect 9950 6780 9956 6792
rect 9355 6752 9956 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 9950 6740 9956 6752
rect 10008 6780 10014 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10008 6752 10793 6780
rect 10008 6740 10014 6752
rect 10781 6749 10793 6752
rect 10827 6780 10839 6783
rect 11808 6780 11836 6876
rect 12268 6857 12296 6888
rect 17696 6888 18828 6916
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 10827 6752 11836 6780
rect 15942 6783 16000 6789
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 15942 6749 15954 6783
rect 15988 6780 16000 6783
rect 16206 6780 16212 6792
rect 15988 6752 16068 6780
rect 16167 6752 16212 6780
rect 15988 6749 16000 6752
rect 15942 6743 16000 6749
rect 16040 6724 16068 6752
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 17696 6789 17724 6888
rect 18322 6848 18328 6860
rect 17972 6820 18328 6848
rect 17972 6789 18000 6820
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 18506 6848 18512 6860
rect 18467 6820 18512 6848
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 17644 6752 17693 6780
rect 17644 6740 17650 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6749 18015 6783
rect 18800 6780 18828 6888
rect 19061 6885 19073 6919
rect 19107 6885 19119 6919
rect 19061 6879 19119 6885
rect 20530 6876 20536 6928
rect 20588 6916 20594 6928
rect 20625 6919 20683 6925
rect 20625 6916 20637 6919
rect 20588 6888 20637 6916
rect 20588 6876 20594 6888
rect 20625 6885 20637 6888
rect 20671 6885 20683 6919
rect 20625 6879 20683 6885
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 21082 6848 21088 6860
rect 20772 6820 21088 6848
rect 20772 6808 20778 6820
rect 21082 6808 21088 6820
rect 21140 6848 21146 6860
rect 21177 6851 21235 6857
rect 21177 6848 21189 6851
rect 21140 6820 21189 6848
rect 21140 6808 21146 6820
rect 21177 6817 21189 6820
rect 21223 6817 21235 6851
rect 21177 6811 21235 6817
rect 17957 6743 18015 6749
rect 18156 6752 18736 6780
rect 18800 6776 19104 6780
rect 19150 6776 19156 6792
rect 18800 6752 19156 6776
rect 7346 6715 7404 6721
rect 7346 6712 7358 6715
rect 6840 6684 7358 6712
rect 6742 6675 6800 6681
rect 7346 6681 7358 6684
rect 7392 6681 7404 6715
rect 7346 6675 7404 6681
rect 9576 6715 9634 6721
rect 9576 6681 9588 6715
rect 9622 6712 9634 6715
rect 9858 6712 9864 6724
rect 9622 6684 9864 6712
rect 9622 6681 9634 6684
rect 9576 6675 9634 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 11048 6715 11106 6721
rect 11048 6681 11060 6715
rect 11094 6712 11106 6715
rect 11146 6712 11152 6724
rect 11094 6684 11152 6712
rect 11094 6681 11106 6684
rect 11048 6675 11106 6681
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 12066 6672 12072 6724
rect 12124 6712 12130 6724
rect 12498 6715 12556 6721
rect 12498 6712 12510 6715
rect 12124 6684 12510 6712
rect 12124 6672 12130 6684
rect 12498 6681 12510 6684
rect 12544 6681 12556 6715
rect 15194 6712 15200 6724
rect 12498 6675 12556 6681
rect 13648 6684 15200 6712
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 3602 6644 3608 6656
rect 2179 6616 3608 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10226 6644 10232 6656
rect 9824 6616 10232 6644
rect 9824 6604 9830 6616
rect 10226 6604 10232 6616
rect 10284 6644 10290 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10284 6616 10701 6644
rect 10284 6604 10290 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 13262 6604 13268 6656
rect 13320 6644 13326 6656
rect 13648 6653 13676 6684
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 16022 6672 16028 6724
rect 16080 6672 16086 6724
rect 16942 6672 16948 6724
rect 17000 6712 17006 6724
rect 17414 6715 17472 6721
rect 17414 6712 17426 6715
rect 17000 6684 17426 6712
rect 17000 6672 17006 6684
rect 17414 6681 17426 6684
rect 17460 6681 17472 6715
rect 17414 6675 17472 6681
rect 13633 6647 13691 6653
rect 13633 6644 13645 6647
rect 13320 6616 13645 6644
rect 13320 6604 13326 6616
rect 13633 6613 13645 6616
rect 13679 6613 13691 6647
rect 13633 6607 13691 6613
rect 14182 6604 14188 6656
rect 14240 6644 14246 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 14240 6616 14473 6644
rect 14240 6604 14246 6616
rect 14461 6613 14473 6616
rect 14507 6644 14519 6647
rect 14734 6644 14740 6656
rect 14507 6616 14740 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 14829 6647 14887 6653
rect 14829 6613 14841 6647
rect 14875 6644 14887 6647
rect 15838 6644 15844 6656
rect 14875 6616 15844 6644
rect 14875 6613 14887 6616
rect 14829 6607 14887 6613
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 16298 6644 16304 6656
rect 16259 6616 16304 6644
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 17494 6604 17500 6656
rect 17552 6644 17558 6656
rect 18156 6653 18184 6752
rect 18598 6712 18604 6724
rect 18559 6684 18604 6712
rect 18598 6672 18604 6684
rect 18656 6672 18662 6724
rect 18708 6712 18736 6752
rect 19076 6748 19156 6752
rect 19150 6740 19156 6748
rect 19208 6780 19214 6792
rect 19242 6780 19248 6792
rect 19208 6752 19248 6780
rect 19208 6740 19214 6752
rect 19242 6740 19248 6752
rect 19300 6780 19306 6792
rect 19794 6780 19800 6792
rect 19300 6752 19800 6780
rect 19300 6740 19306 6752
rect 19794 6740 19800 6752
rect 19852 6780 19858 6792
rect 20898 6780 20904 6792
rect 19852 6752 20208 6780
rect 20859 6752 20904 6780
rect 19852 6740 19858 6752
rect 20180 6724 20208 6752
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 21192 6780 21220 6811
rect 21634 6808 21640 6860
rect 21692 6848 21698 6860
rect 21913 6851 21971 6857
rect 21692 6820 21737 6848
rect 21692 6808 21698 6820
rect 21913 6817 21925 6851
rect 21959 6848 21971 6851
rect 22278 6848 22284 6860
rect 21959 6820 22284 6848
rect 21959 6817 21971 6820
rect 21913 6811 21971 6817
rect 22278 6808 22284 6820
rect 22336 6848 22342 6860
rect 23124 6848 23152 6944
rect 23382 6848 23388 6860
rect 22336 6820 23388 6848
rect 22336 6808 22342 6820
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 22554 6780 22560 6792
rect 21192 6752 22560 6780
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 19334 6712 19340 6724
rect 18708 6684 19340 6712
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 19512 6715 19570 6721
rect 19512 6681 19524 6715
rect 19558 6712 19570 6715
rect 19610 6712 19616 6724
rect 19558 6684 19616 6712
rect 19558 6681 19570 6684
rect 19512 6675 19570 6681
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 20162 6672 20168 6724
rect 20220 6672 20226 6724
rect 20717 6715 20775 6721
rect 20717 6681 20729 6715
rect 20763 6712 20775 6715
rect 20806 6712 20812 6724
rect 20763 6684 20812 6712
rect 20763 6681 20775 6684
rect 20717 6675 20775 6681
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 17773 6647 17831 6653
rect 17773 6644 17785 6647
rect 17552 6616 17785 6644
rect 17552 6604 17558 6616
rect 17773 6613 17785 6616
rect 17819 6613 17831 6647
rect 17773 6607 17831 6613
rect 18141 6647 18199 6653
rect 18141 6613 18153 6647
rect 18187 6613 18199 6647
rect 18141 6607 18199 6613
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18693 6647 18751 6653
rect 18693 6644 18705 6647
rect 18380 6616 18705 6644
rect 18380 6604 18386 6616
rect 18693 6613 18705 6616
rect 18739 6613 18751 6647
rect 18693 6607 18751 6613
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 20622 6644 20628 6656
rect 19208 6616 20628 6644
rect 19208 6604 19214 6616
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 21082 6644 21088 6656
rect 21043 6616 21088 6644
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 21643 6647 21701 6653
rect 21643 6644 21655 6647
rect 21600 6616 21655 6644
rect 21600 6604 21606 6616
rect 21643 6613 21655 6616
rect 21689 6613 21701 6647
rect 21643 6607 21701 6613
rect 22646 6604 22652 6656
rect 22704 6644 22710 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22704 6616 23029 6644
rect 22704 6604 22710 6616
rect 23017 6613 23029 6616
rect 23063 6613 23075 6647
rect 23017 6607 23075 6613
rect 1104 6554 23460 6576
rect 1104 6502 6548 6554
rect 6600 6502 6612 6554
rect 6664 6502 6676 6554
rect 6728 6502 6740 6554
rect 6792 6502 6804 6554
rect 6856 6502 12146 6554
rect 12198 6502 12210 6554
rect 12262 6502 12274 6554
rect 12326 6502 12338 6554
rect 12390 6502 12402 6554
rect 12454 6502 17744 6554
rect 17796 6502 17808 6554
rect 17860 6502 17872 6554
rect 17924 6502 17936 6554
rect 17988 6502 18000 6554
rect 18052 6502 23460 6554
rect 1104 6480 23460 6502
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8849 6443 8907 6449
rect 8849 6409 8861 6443
rect 8895 6440 8907 6443
rect 9858 6440 9864 6452
rect 8895 6412 9864 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10505 6443 10563 6449
rect 10505 6409 10517 6443
rect 10551 6440 10563 6443
rect 11238 6440 11244 6452
rect 10551 6412 11244 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 13725 6443 13783 6449
rect 11532 6412 13492 6440
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 7662 6375 7720 6381
rect 7662 6372 7674 6375
rect 5960 6344 7674 6372
rect 5960 6332 5966 6344
rect 7662 6341 7674 6344
rect 7708 6341 7720 6375
rect 8404 6372 8432 6400
rect 7662 6335 7720 6341
rect 7944 6344 8432 6372
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 7944 6313 7972 6344
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 8941 6375 8999 6381
rect 8941 6372 8953 6375
rect 8812 6344 8953 6372
rect 8812 6332 8818 6344
rect 8941 6341 8953 6344
rect 8987 6341 8999 6375
rect 9766 6372 9772 6384
rect 9727 6344 9772 6372
rect 8941 6335 8999 6341
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 10597 6375 10655 6381
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 10870 6372 10876 6384
rect 10643 6344 10876 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 7929 6307 7987 6313
rect 2188 6276 7880 6304
rect 2188 6264 2194 6276
rect 7852 6236 7880 6276
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8251 6276 9536 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8938 6236 8944 6248
rect 7852 6208 8944 6236
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9122 6236 9128 6248
rect 9035 6208 9128 6236
rect 9122 6196 9128 6208
rect 9180 6236 9186 6248
rect 9180 6208 9444 6236
rect 9180 6196 9186 6208
rect 6546 6100 6552 6112
rect 6507 6072 6552 6100
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 8018 6100 8024 6112
rect 7979 6072 8024 6100
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8478 6100 8484 6112
rect 8439 6072 8484 6100
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9309 6103 9367 6109
rect 9309 6100 9321 6103
rect 9272 6072 9321 6100
rect 9272 6060 9278 6072
rect 9309 6069 9321 6072
rect 9355 6069 9367 6103
rect 9416 6100 9444 6208
rect 9508 6168 9536 6276
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 11149 6307 11207 6313
rect 11149 6304 11161 6307
rect 9732 6276 9777 6304
rect 9968 6276 11161 6304
rect 9732 6264 9738 6276
rect 9968 6245 9996 6276
rect 11149 6273 11161 6276
rect 11195 6304 11207 6307
rect 11330 6304 11336 6316
rect 11195 6276 11336 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11532 6313 11560 6412
rect 13170 6332 13176 6384
rect 13228 6332 13234 6384
rect 13262 6332 13268 6384
rect 13320 6381 13326 6384
rect 13320 6372 13332 6381
rect 13320 6344 13365 6372
rect 13320 6335 13332 6344
rect 13320 6332 13326 6335
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 13188 6304 13216 6332
rect 12023 6276 13216 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6205 10011 6239
rect 10778 6236 10784 6248
rect 10739 6208 10784 6236
rect 9953 6199 10011 6205
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 12526 6236 12532 6248
rect 11532 6208 12532 6236
rect 11532 6180 11560 6208
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 13464 6236 13492 6412
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 13906 6440 13912 6452
rect 13771 6412 13912 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 13740 6304 13768 6403
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6440 14519 6443
rect 16574 6440 16580 6452
rect 14507 6412 16580 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 18138 6400 18144 6452
rect 18196 6440 18202 6452
rect 18690 6440 18696 6452
rect 18196 6412 18696 6440
rect 18196 6400 18202 6412
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 20714 6440 20720 6452
rect 19076 6412 20720 6440
rect 14274 6332 14280 6384
rect 14332 6372 14338 6384
rect 15565 6375 15623 6381
rect 14332 6344 14780 6372
rect 14332 6332 14338 6344
rect 13587 6276 13768 6304
rect 14369 6307 14427 6313
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 14369 6273 14381 6307
rect 14415 6304 14427 6307
rect 14642 6304 14648 6316
rect 14415 6276 14648 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 14274 6236 14280 6248
rect 13464 6208 14280 6236
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 14752 6236 14780 6344
rect 15565 6341 15577 6375
rect 15611 6372 15623 6375
rect 16666 6372 16672 6384
rect 15611 6344 16672 6372
rect 15611 6341 15623 6344
rect 15565 6335 15623 6341
rect 16666 6332 16672 6344
rect 16724 6332 16730 6384
rect 17126 6332 17132 6384
rect 17184 6372 17190 6384
rect 19076 6372 19104 6412
rect 20714 6400 20720 6412
rect 20772 6400 20778 6452
rect 20898 6440 20904 6452
rect 20859 6412 20904 6440
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 21232 6412 21281 6440
rect 21232 6400 21238 6412
rect 21269 6409 21281 6412
rect 21315 6409 21327 6443
rect 21269 6403 21327 6409
rect 22741 6443 22799 6449
rect 22741 6409 22753 6443
rect 22787 6440 22799 6443
rect 23014 6440 23020 6452
rect 22787 6412 23020 6440
rect 22787 6409 22799 6412
rect 22741 6403 22799 6409
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 20104 6375 20162 6381
rect 20104 6372 20116 6375
rect 17184 6344 19104 6372
rect 19168 6344 20116 6372
rect 17184 6332 17190 6344
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14884 6276 15025 6304
rect 14884 6264 14890 6276
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15519 6276 15945 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16761 6307 16819 6313
rect 16761 6273 16773 6307
rect 16807 6304 16819 6307
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 16807 6276 17509 6304
rect 16807 6273 16819 6276
rect 16761 6267 16819 6273
rect 17497 6273 17509 6276
rect 17543 6304 17555 6307
rect 17586 6304 17592 6316
rect 17543 6276 17592 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 14608 6208 14653 6236
rect 14752 6208 15669 6236
rect 14608 6196 14614 6208
rect 15657 6205 15669 6208
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 10137 6171 10195 6177
rect 10137 6168 10149 6171
rect 9508 6140 10149 6168
rect 10137 6137 10149 6140
rect 10183 6137 10195 6171
rect 10137 6131 10195 6137
rect 11514 6128 11520 6180
rect 11572 6128 11578 6180
rect 11701 6171 11759 6177
rect 11701 6137 11713 6171
rect 11747 6168 11759 6171
rect 11974 6168 11980 6180
rect 11747 6140 11980 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 15105 6171 15163 6177
rect 15105 6137 15117 6171
rect 15151 6168 15163 6171
rect 15378 6168 15384 6180
rect 15151 6140 15384 6168
rect 15151 6137 15163 6140
rect 15105 6131 15163 6137
rect 15378 6128 15384 6140
rect 15436 6128 15442 6180
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 9416 6072 11069 6100
rect 9309 6063 9367 6069
rect 11057 6069 11069 6072
rect 11103 6069 11115 6103
rect 11057 6063 11115 6069
rect 11793 6103 11851 6109
rect 11793 6069 11805 6103
rect 11839 6100 11851 6103
rect 11882 6100 11888 6112
rect 11839 6072 11888 6100
rect 11839 6069 11851 6072
rect 11793 6063 11851 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12161 6103 12219 6109
rect 12161 6069 12173 6103
rect 12207 6100 12219 6103
rect 12894 6100 12900 6112
rect 12207 6072 12900 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13538 6060 13544 6112
rect 13596 6100 13602 6112
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13596 6072 14013 6100
rect 13596 6060 13602 6072
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 14090 6060 14096 6112
rect 14148 6100 14154 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14148 6072 14841 6100
rect 14148 6060 14154 6072
rect 14829 6069 14841 6072
rect 14875 6100 14887 6103
rect 15470 6100 15476 6112
rect 14875 6072 15476 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 15470 6060 15476 6072
rect 15528 6100 15534 6112
rect 16224 6100 16252 6267
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 17764 6307 17822 6313
rect 17764 6273 17776 6307
rect 17810 6304 17822 6307
rect 18690 6304 18696 6316
rect 17810 6276 18696 6304
rect 17810 6273 17822 6276
rect 17764 6267 17822 6273
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 19168 6304 19196 6344
rect 20104 6341 20116 6344
rect 20150 6372 20162 6375
rect 20530 6372 20536 6384
rect 20150 6344 20536 6372
rect 20150 6341 20162 6344
rect 20104 6335 20162 6341
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 22186 6372 22192 6384
rect 20640 6344 22094 6372
rect 22147 6344 22192 6372
rect 18800 6276 19196 6304
rect 17129 6239 17187 6245
rect 17129 6205 17141 6239
rect 17175 6205 17187 6239
rect 17402 6236 17408 6248
rect 17363 6208 17408 6236
rect 17129 6199 17187 6205
rect 17144 6168 17172 6199
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18800 6236 18828 6276
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 20640 6313 20668 6344
rect 20625 6307 20683 6313
rect 19300 6276 20484 6304
rect 19300 6264 19306 6276
rect 20349 6239 20407 6245
rect 18564 6208 18828 6236
rect 18984 6208 19334 6236
rect 18564 6196 18570 6208
rect 18984 6168 19012 6208
rect 17144 6140 17540 6168
rect 15528 6072 16252 6100
rect 16393 6103 16451 6109
rect 15528 6060 15534 6072
rect 16393 6069 16405 6103
rect 16439 6100 16451 6103
rect 17126 6100 17132 6112
rect 16439 6072 17132 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 17126 6060 17132 6072
rect 17184 6060 17190 6112
rect 17512 6100 17540 6140
rect 18423 6140 19012 6168
rect 19306 6168 19334 6208
rect 20349 6205 20361 6239
rect 20395 6205 20407 6239
rect 20456 6236 20484 6276
rect 20625 6273 20637 6307
rect 20671 6273 20683 6307
rect 22066 6304 22094 6344
rect 22186 6332 22192 6344
rect 22244 6332 22250 6384
rect 22278 6332 22284 6384
rect 22336 6372 22342 6384
rect 23474 6372 23480 6384
rect 22336 6344 22381 6372
rect 22756 6344 23480 6372
rect 22336 6332 22342 6344
rect 22756 6304 22784 6344
rect 23474 6332 23480 6344
rect 23532 6332 23538 6384
rect 20625 6267 20683 6273
rect 20732 6276 21496 6304
rect 22066 6276 22784 6304
rect 22833 6307 22891 6313
rect 20732 6236 20760 6276
rect 21358 6236 21364 6248
rect 20456 6208 20760 6236
rect 21319 6208 21364 6236
rect 20349 6199 20407 6205
rect 19306 6140 19472 6168
rect 18423 6100 18451 6140
rect 17512 6072 18451 6100
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 18877 6103 18935 6109
rect 18877 6100 18889 6103
rect 18840 6072 18889 6100
rect 18840 6060 18846 6072
rect 18877 6069 18889 6072
rect 18923 6069 18935 6103
rect 18877 6063 18935 6069
rect 18966 6060 18972 6112
rect 19024 6100 19030 6112
rect 19444 6100 19472 6140
rect 19978 6100 19984 6112
rect 19024 6072 19069 6100
rect 19444 6072 19984 6100
rect 19024 6060 19030 6072
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 20162 6060 20168 6112
rect 20220 6100 20226 6112
rect 20364 6100 20392 6199
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 21468 6245 21496 6276
rect 22833 6273 22845 6307
rect 22879 6304 22891 6307
rect 23290 6304 23296 6316
rect 22879 6276 23296 6304
rect 22879 6273 22891 6276
rect 22833 6267 22891 6273
rect 23290 6264 23296 6276
rect 23348 6264 23354 6316
rect 21453 6239 21511 6245
rect 21453 6205 21465 6239
rect 21499 6205 21511 6239
rect 21453 6199 21511 6205
rect 21818 6196 21824 6248
rect 21876 6236 21882 6248
rect 21876 6208 22094 6236
rect 21876 6196 21882 6208
rect 20809 6171 20867 6177
rect 20809 6137 20821 6171
rect 20855 6168 20867 6171
rect 21726 6168 21732 6180
rect 20855 6140 21732 6168
rect 20855 6137 20867 6140
rect 20809 6131 20867 6137
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 22066 6168 22094 6208
rect 22370 6196 22376 6248
rect 22428 6236 22434 6248
rect 22428 6208 22473 6236
rect 22428 6196 22434 6208
rect 22830 6168 22836 6180
rect 22066 6140 22836 6168
rect 22830 6128 22836 6140
rect 22888 6128 22894 6180
rect 23017 6171 23075 6177
rect 23017 6137 23029 6171
rect 23063 6168 23075 6171
rect 23106 6168 23112 6180
rect 23063 6140 23112 6168
rect 23063 6137 23075 6140
rect 23017 6131 23075 6137
rect 23106 6128 23112 6140
rect 23164 6128 23170 6180
rect 20441 6103 20499 6109
rect 20441 6100 20453 6103
rect 20220 6072 20453 6100
rect 20220 6060 20226 6072
rect 20441 6069 20453 6072
rect 20487 6069 20499 6103
rect 21818 6100 21824 6112
rect 21779 6072 21824 6100
rect 20441 6063 20499 6069
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 1104 6010 23460 6032
rect 1104 5958 3749 6010
rect 3801 5958 3813 6010
rect 3865 5958 3877 6010
rect 3929 5958 3941 6010
rect 3993 5958 4005 6010
rect 4057 5958 9347 6010
rect 9399 5958 9411 6010
rect 9463 5958 9475 6010
rect 9527 5958 9539 6010
rect 9591 5958 9603 6010
rect 9655 5958 14945 6010
rect 14997 5958 15009 6010
rect 15061 5958 15073 6010
rect 15125 5958 15137 6010
rect 15189 5958 15201 6010
rect 15253 5958 20543 6010
rect 20595 5958 20607 6010
rect 20659 5958 20671 6010
rect 20723 5958 20735 6010
rect 20787 5958 20799 6010
rect 20851 5958 23460 6010
rect 1104 5936 23460 5958
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 5920 5868 7481 5896
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5350 5760 5356 5772
rect 5311 5732 5356 5760
rect 5169 5723 5227 5729
rect 5184 5624 5212 5723
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 5920 5769 5948 5868
rect 7469 5865 7481 5868
rect 7515 5896 7527 5899
rect 8386 5896 8392 5908
rect 7515 5868 8392 5896
rect 7515 5865 7527 5868
rect 7469 5859 7527 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 11609 5899 11667 5905
rect 11609 5896 11621 5899
rect 8720 5868 11621 5896
rect 8720 5856 8726 5868
rect 11609 5865 11621 5868
rect 11655 5865 11667 5899
rect 11609 5859 11667 5865
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11756 5868 11897 5896
rect 11756 5856 11762 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 12345 5899 12403 5905
rect 12345 5865 12357 5899
rect 12391 5896 12403 5899
rect 12618 5896 12624 5908
rect 12391 5868 12624 5896
rect 12391 5865 12403 5868
rect 12345 5859 12403 5865
rect 7006 5788 7012 5840
rect 7064 5828 7070 5840
rect 9033 5831 9091 5837
rect 9033 5828 9045 5831
rect 7064 5800 9045 5828
rect 7064 5788 7070 5800
rect 9033 5797 9045 5800
rect 9079 5797 9091 5831
rect 9953 5831 10011 5837
rect 9953 5828 9965 5831
rect 9033 5791 9091 5797
rect 9692 5800 9965 5828
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5729 5963 5763
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 5905 5723 5963 5729
rect 6932 5732 8401 5760
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5692 5503 5695
rect 5718 5692 5724 5704
rect 5491 5664 5724 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 6172 5695 6230 5701
rect 6172 5692 6184 5695
rect 5868 5664 6184 5692
rect 5868 5652 5874 5664
rect 6172 5661 6184 5664
rect 6218 5692 6230 5695
rect 6546 5692 6552 5704
rect 6218 5664 6552 5692
rect 6218 5661 6230 5664
rect 6172 5655 6230 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 5626 5624 5632 5636
rect 5184 5596 5632 5624
rect 5626 5584 5632 5596
rect 5684 5624 5690 5636
rect 6932 5624 6960 5732
rect 8389 5729 8401 5732
rect 8435 5760 8447 5763
rect 9122 5760 9128 5772
rect 8435 5732 9128 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9214 5720 9220 5772
rect 9272 5760 9278 5772
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 9272 5732 9505 5760
rect 9272 5720 9278 5732
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9692 5769 9720 5800
rect 9953 5797 9965 5800
rect 9999 5828 10011 5831
rect 10778 5828 10784 5840
rect 9999 5800 10784 5828
rect 9999 5797 10011 5800
rect 9953 5791 10011 5797
rect 10778 5788 10784 5800
rect 10836 5828 10842 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 10836 5800 10977 5828
rect 10836 5788 10842 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 11422 5828 11428 5840
rect 11383 5800 11428 5828
rect 10965 5791 11023 5797
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9640 5732 9689 5760
rect 9640 5720 9646 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 10873 5763 10931 5769
rect 10873 5729 10885 5763
rect 10919 5760 10931 5763
rect 12360 5760 12388 5859
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 14550 5896 14556 5908
rect 13924 5868 14556 5896
rect 13924 5837 13952 5868
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17000 5868 19840 5896
rect 17000 5856 17006 5868
rect 13909 5831 13967 5837
rect 13909 5797 13921 5831
rect 13955 5797 13967 5831
rect 17218 5828 17224 5840
rect 13909 5791 13967 5797
rect 15948 5800 17224 5828
rect 10919 5732 12388 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 13228 5732 13277 5760
rect 13228 5720 13234 5732
rect 13265 5729 13277 5732
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 13449 5763 13507 5769
rect 13449 5729 13461 5763
rect 13495 5760 13507 5763
rect 13538 5760 13544 5772
rect 13495 5732 13544 5760
rect 13495 5729 13507 5732
rect 13449 5723 13507 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 14090 5720 14096 5772
rect 14148 5760 14154 5772
rect 14148 5732 14193 5760
rect 14148 5720 14154 5732
rect 14550 5720 14556 5772
rect 14608 5758 14614 5772
rect 14608 5730 14651 5758
rect 14608 5720 14614 5730
rect 14734 5720 14740 5772
rect 14792 5760 14798 5772
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 14792 5732 14841 5760
rect 14792 5720 14798 5732
rect 14829 5729 14841 5732
rect 14875 5760 14887 5763
rect 15948 5760 15976 5800
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 19058 5828 19064 5840
rect 19019 5800 19064 5828
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 16114 5760 16120 5772
rect 14875 5732 15976 5760
rect 16075 5732 16120 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 17494 5720 17500 5772
rect 17552 5760 17558 5772
rect 19812 5769 19840 5868
rect 19978 5856 19984 5908
rect 20036 5896 20042 5908
rect 20898 5896 20904 5908
rect 20036 5868 20904 5896
rect 20036 5856 20042 5868
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 21726 5856 21732 5908
rect 21784 5896 21790 5908
rect 22094 5896 22100 5908
rect 21784 5868 22100 5896
rect 21784 5856 21790 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 23014 5896 23020 5908
rect 22975 5868 23020 5896
rect 23014 5856 23020 5868
rect 23072 5856 23078 5908
rect 20438 5788 20444 5840
rect 20496 5828 20502 5840
rect 20625 5831 20683 5837
rect 20625 5828 20637 5831
rect 20496 5800 20637 5828
rect 20496 5788 20502 5800
rect 20625 5797 20637 5800
rect 20671 5797 20683 5831
rect 20625 5791 20683 5797
rect 17684 5763 17742 5769
rect 17684 5760 17696 5763
rect 17552 5732 17696 5760
rect 17552 5720 17558 5732
rect 17684 5729 17696 5732
rect 17730 5729 17742 5763
rect 19797 5763 19855 5769
rect 17684 5723 17742 5729
rect 19306 5732 19656 5760
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 9088 5664 9413 5692
rect 9088 5652 9094 5664
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 11238 5692 11244 5704
rect 11199 5664 11244 5692
rect 9401 5655 9459 5661
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11698 5652 11704 5704
rect 11756 5692 11762 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11756 5664 11805 5692
rect 11756 5652 11762 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16574 5692 16580 5704
rect 16439 5664 16580 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 17126 5652 17132 5704
rect 17184 5692 17190 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 17184 5664 17233 5692
rect 17184 5652 17190 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 17644 5664 17969 5692
rect 17644 5652 17650 5664
rect 17957 5661 17969 5664
rect 18003 5692 18015 5695
rect 18598 5692 18604 5704
rect 18003 5664 18604 5692
rect 18003 5661 18015 5664
rect 17957 5655 18015 5661
rect 18598 5652 18604 5664
rect 18656 5692 18662 5704
rect 19306 5692 19334 5732
rect 19628 5701 19656 5732
rect 19797 5729 19809 5763
rect 19843 5729 19855 5763
rect 19797 5723 19855 5729
rect 19904 5732 21128 5760
rect 18656 5664 19334 5692
rect 19613 5695 19671 5701
rect 18656 5652 18662 5664
rect 19613 5661 19625 5695
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 8205 5627 8263 5633
rect 8205 5624 8217 5627
rect 5684 5596 6960 5624
rect 7300 5596 8217 5624
rect 5684 5584 5690 5596
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6914 5556 6920 5568
rect 5859 5528 6920 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7300 5565 7328 5596
rect 8205 5593 8217 5596
rect 8251 5593 8263 5627
rect 8205 5587 8263 5593
rect 16206 5584 16212 5636
rect 16264 5624 16270 5636
rect 16945 5627 17003 5633
rect 16945 5624 16957 5627
rect 16264 5596 16957 5624
rect 16264 5584 16270 5596
rect 16945 5593 16957 5596
rect 16991 5593 17003 5627
rect 19904 5624 19932 5732
rect 20070 5692 20076 5704
rect 20031 5664 20076 5692
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 16945 5587 17003 5593
rect 19076 5596 19932 5624
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 7156 5528 7297 5556
rect 7156 5516 7162 5528
rect 7285 5525 7297 5528
rect 7331 5525 7343 5559
rect 7742 5556 7748 5568
rect 7703 5528 7748 5556
rect 7285 5519 7343 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 13596 5528 13641 5556
rect 13596 5516 13602 5528
rect 14366 5516 14372 5568
rect 14424 5556 14430 5568
rect 14559 5559 14617 5565
rect 14559 5556 14571 5559
rect 14424 5528 14571 5556
rect 14424 5516 14430 5528
rect 14559 5525 14571 5528
rect 14605 5525 14617 5559
rect 14559 5519 14617 5525
rect 15933 5559 15991 5565
rect 15933 5525 15945 5559
rect 15979 5556 15991 5559
rect 16298 5556 16304 5568
rect 15979 5528 16304 5556
rect 15979 5525 15991 5528
rect 15933 5519 15991 5525
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 16761 5559 16819 5565
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 16850 5556 16856 5568
rect 16807 5528 16856 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17037 5559 17095 5565
rect 17037 5525 17049 5559
rect 17083 5556 17095 5559
rect 17687 5559 17745 5565
rect 17687 5556 17699 5559
rect 17083 5528 17699 5556
rect 17083 5525 17095 5528
rect 17037 5519 17095 5525
rect 17687 5525 17699 5528
rect 17733 5556 17745 5559
rect 19076 5556 19104 5596
rect 20162 5584 20168 5636
rect 20220 5624 20226 5636
rect 20349 5627 20407 5633
rect 20349 5624 20361 5627
rect 20220 5596 20361 5624
rect 20220 5584 20226 5596
rect 20349 5593 20361 5596
rect 20395 5593 20407 5627
rect 20349 5587 20407 5593
rect 17733 5528 19104 5556
rect 17733 5525 17745 5528
rect 17687 5519 17745 5525
rect 19150 5516 19156 5568
rect 19208 5556 19214 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 19208 5528 19257 5556
rect 19208 5516 19214 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19245 5519 19303 5525
rect 19705 5559 19763 5565
rect 19705 5525 19717 5559
rect 19751 5556 19763 5559
rect 20070 5556 20076 5568
rect 19751 5528 20076 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 21100 5556 21128 5732
rect 21910 5720 21916 5772
rect 21968 5760 21974 5772
rect 22002 5763 22060 5769
rect 22002 5760 22014 5763
rect 21968 5732 22014 5760
rect 21968 5720 21974 5732
rect 22002 5729 22014 5732
rect 22048 5729 22060 5763
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 22002 5723 22060 5729
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 23658 5760 23664 5772
rect 22756 5732 23664 5760
rect 21174 5668 21180 5720
rect 21232 5692 21238 5720
rect 22756 5701 22784 5732
rect 23658 5720 23664 5732
rect 23716 5720 23722 5772
rect 21729 5695 21787 5701
rect 21729 5692 21741 5695
rect 21232 5668 21741 5692
rect 21192 5664 21741 5668
rect 21729 5661 21741 5664
rect 21775 5661 21787 5695
rect 21729 5655 21787 5661
rect 22741 5695 22799 5701
rect 22741 5661 22753 5695
rect 22787 5661 22799 5695
rect 22741 5655 22799 5661
rect 22830 5652 22836 5704
rect 22888 5692 22894 5704
rect 22888 5664 22933 5692
rect 22888 5652 22894 5664
rect 21450 5556 21456 5568
rect 21100 5528 21456 5556
rect 21450 5516 21456 5528
rect 21508 5556 21514 5568
rect 21998 5559 22056 5565
rect 21998 5556 22010 5559
rect 21508 5528 22010 5556
rect 21508 5516 21514 5528
rect 21998 5525 22010 5528
rect 22044 5525 22056 5559
rect 22554 5556 22560 5568
rect 22515 5528 22560 5556
rect 21998 5519 22056 5525
rect 22554 5516 22560 5528
rect 22612 5516 22618 5568
rect 1104 5466 23460 5488
rect 1104 5414 6548 5466
rect 6600 5414 6612 5466
rect 6664 5414 6676 5466
rect 6728 5414 6740 5466
rect 6792 5414 6804 5466
rect 6856 5414 12146 5466
rect 12198 5414 12210 5466
rect 12262 5414 12274 5466
rect 12326 5414 12338 5466
rect 12390 5414 12402 5466
rect 12454 5414 17744 5466
rect 17796 5414 17808 5466
rect 17860 5414 17872 5466
rect 17924 5414 17936 5466
rect 17988 5414 18000 5466
rect 18052 5414 23460 5466
rect 1104 5392 23460 5414
rect 5810 5352 5816 5364
rect 5771 5324 5816 5352
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5352 6791 5355
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 6779 5324 7113 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 7101 5321 7113 5324
rect 7147 5321 7159 5355
rect 7101 5315 7159 5321
rect 7193 5355 7251 5361
rect 7193 5321 7205 5355
rect 7239 5352 7251 5355
rect 8018 5352 8024 5364
rect 7239 5324 8024 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 9582 5352 9588 5364
rect 8619 5324 9588 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 5721 5287 5779 5293
rect 5721 5253 5733 5287
rect 5767 5284 5779 5287
rect 5902 5284 5908 5296
rect 5767 5256 5908 5284
rect 5767 5253 5779 5256
rect 5721 5247 5779 5253
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 8113 5287 8171 5293
rect 8113 5284 8125 5287
rect 6972 5256 8125 5284
rect 6972 5244 6978 5256
rect 8113 5253 8125 5256
rect 8159 5253 8171 5287
rect 8113 5247 8171 5253
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 7006 5216 7012 5228
rect 6595 5188 7012 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 8478 5216 8484 5228
rect 8067 5188 8484 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 5626 5148 5632 5160
rect 5587 5120 5632 5148
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 6914 5148 6920 5160
rect 6827 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5148 6978 5160
rect 7834 5148 7840 5160
rect 6972 5120 7840 5148
rect 6972 5108 6978 5120
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5148 8355 5151
rect 8386 5148 8392 5160
rect 8343 5120 8392 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 8386 5108 8392 5120
rect 8444 5148 8450 5160
rect 8588 5148 8616 5315
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 9977 5324 10977 5352
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9977 5225 10005 5324
rect 10965 5321 10977 5324
rect 11011 5352 11023 5355
rect 11054 5352 11060 5364
rect 11011 5324 11060 5352
rect 11011 5321 11023 5324
rect 10965 5315 11023 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 13538 5352 13544 5364
rect 13499 5324 13544 5352
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 15019 5355 15077 5361
rect 15019 5352 15031 5355
rect 14047 5324 15031 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 15019 5321 15031 5324
rect 15065 5352 15077 5355
rect 16206 5352 16212 5364
rect 15065 5324 16212 5352
rect 15065 5321 15077 5324
rect 15019 5315 15077 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 17494 5352 17500 5364
rect 17455 5324 17500 5352
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 17957 5355 18015 5361
rect 17957 5321 17969 5355
rect 18003 5352 18015 5355
rect 19150 5352 19156 5364
rect 18003 5324 19156 5352
rect 18003 5321 18015 5324
rect 17957 5315 18015 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 20070 5352 20076 5364
rect 19260 5324 20076 5352
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 13909 5287 13967 5293
rect 13909 5284 13921 5287
rect 10928 5256 13921 5284
rect 10928 5244 10934 5256
rect 13909 5253 13921 5256
rect 13955 5284 13967 5287
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13955 5256 14197 5284
rect 13955 5253 13967 5256
rect 13909 5247 13967 5253
rect 14185 5253 14197 5256
rect 14231 5284 14243 5287
rect 14366 5284 14372 5296
rect 14231 5256 14372 5284
rect 14231 5253 14243 5256
rect 14185 5247 14243 5253
rect 14366 5244 14372 5256
rect 14424 5244 14430 5296
rect 16390 5244 16396 5296
rect 16448 5284 16454 5296
rect 16448 5256 17448 5284
rect 16448 5244 16454 5256
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 8996 5188 9965 5216
rect 8996 5176 9002 5188
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 10689 5219 10747 5225
rect 10689 5216 10701 5219
rect 9953 5179 10011 5185
rect 10060 5188 10701 5216
rect 8444 5120 8616 5148
rect 8444 5108 8450 5120
rect 10060 5092 10088 5188
rect 10689 5185 10701 5188
rect 10735 5185 10747 5219
rect 15286 5216 15292 5228
rect 15247 5188 15292 5216
rect 10689 5179 10747 5185
rect 15286 5176 15292 5188
rect 15344 5216 15350 5228
rect 16022 5216 16028 5228
rect 15344 5188 16028 5216
rect 15344 5176 15350 5188
rect 16022 5176 16028 5188
rect 16080 5216 16086 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16080 5188 17049 5216
rect 16080 5176 16086 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17310 5216 17316 5228
rect 17175 5188 17316 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 10192 5120 10241 5148
rect 10192 5108 10198 5120
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 10778 5148 10784 5160
rect 10275 5120 10784 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5148 14611 5151
rect 14826 5148 14832 5160
rect 14599 5120 14832 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 15059 5151 15117 5157
rect 15059 5117 15071 5151
rect 15105 5148 15117 5151
rect 15378 5148 15384 5160
rect 15105 5120 15384 5148
rect 15105 5117 15117 5120
rect 15059 5111 15117 5117
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 15930 5108 15936 5160
rect 15988 5148 15994 5160
rect 17221 5151 17279 5157
rect 17221 5148 17233 5151
rect 15988 5120 17233 5148
rect 15988 5108 15994 5120
rect 17221 5117 17233 5120
rect 17267 5117 17279 5151
rect 17420 5148 17448 5256
rect 18782 5244 18788 5296
rect 18840 5284 18846 5296
rect 19260 5284 19288 5324
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 20254 5312 20260 5364
rect 20312 5352 20318 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 20312 5324 20637 5352
rect 20312 5312 20318 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20990 5352 20996 5364
rect 20951 5324 20996 5352
rect 20625 5315 20683 5321
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 21358 5312 21364 5364
rect 21416 5352 21422 5364
rect 21913 5355 21971 5361
rect 21913 5352 21925 5355
rect 21416 5324 21925 5352
rect 21416 5312 21422 5324
rect 21913 5321 21925 5324
rect 21959 5321 21971 5355
rect 22278 5352 22284 5364
rect 22239 5324 22284 5352
rect 21913 5315 21971 5321
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 22373 5355 22431 5361
rect 22373 5321 22385 5355
rect 22419 5352 22431 5355
rect 22646 5352 22652 5364
rect 22419 5324 22652 5352
rect 22419 5321 22431 5324
rect 22373 5315 22431 5321
rect 22646 5312 22652 5324
rect 22704 5312 22710 5364
rect 22922 5352 22928 5364
rect 22883 5324 22928 5352
rect 22922 5312 22928 5324
rect 22980 5312 22986 5364
rect 20530 5284 20536 5296
rect 18840 5256 19288 5284
rect 20491 5256 20536 5284
rect 18840 5244 18846 5256
rect 20530 5244 20536 5256
rect 20588 5244 20594 5296
rect 22186 5244 22192 5296
rect 22244 5284 22250 5296
rect 22244 5256 22508 5284
rect 22244 5244 22250 5256
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 17911 5188 18337 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 19817 5219 19875 5225
rect 19817 5185 19829 5219
rect 19863 5216 19875 5219
rect 19978 5216 19984 5228
rect 19863 5188 19984 5216
rect 19863 5185 19875 5188
rect 19817 5179 19875 5185
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 21542 5216 21548 5228
rect 21503 5188 21548 5216
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17420 5120 18061 5148
rect 17221 5111 17279 5117
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5148 20131 5151
rect 20162 5148 20168 5160
rect 20119 5120 20168 5148
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 20162 5108 20168 5120
rect 20220 5108 20226 5160
rect 22480 5157 22508 5256
rect 22554 5176 22560 5228
rect 22612 5216 22618 5228
rect 22741 5219 22799 5225
rect 22741 5216 22753 5219
rect 22612 5188 22753 5216
rect 22612 5176 22618 5188
rect 22741 5185 22753 5188
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 20717 5151 20775 5157
rect 20717 5148 20729 5151
rect 20272 5120 20729 5148
rect 7561 5083 7619 5089
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 10042 5080 10048 5092
rect 7607 5052 10048 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 10042 5040 10048 5052
rect 10100 5040 10106 5092
rect 10873 5083 10931 5089
rect 10873 5049 10885 5083
rect 10919 5080 10931 5083
rect 14366 5080 14372 5092
rect 10919 5052 14372 5080
rect 10919 5049 10931 5052
rect 10873 5043 10931 5049
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 20272 5080 20300 5120
rect 20717 5117 20729 5120
rect 20763 5117 20775 5151
rect 20717 5111 20775 5117
rect 22465 5151 22523 5157
rect 22465 5117 22477 5151
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 20088 5052 20300 5080
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 7466 5012 7472 5024
rect 6227 4984 7472 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 7708 4984 7753 5012
rect 7708 4972 7714 4984
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8757 5015 8815 5021
rect 8757 5012 8769 5015
rect 7892 4984 8769 5012
rect 7892 4972 7898 4984
rect 8757 4981 8769 4984
rect 8803 5012 8815 5015
rect 10686 5012 10692 5024
rect 8803 4984 10692 5012
rect 8803 4981 8815 4984
rect 8757 4975 8815 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16393 5015 16451 5021
rect 16393 5012 16405 5015
rect 16172 4984 16405 5012
rect 16172 4972 16178 4984
rect 16393 4981 16405 4984
rect 16439 4981 16451 5015
rect 18690 5012 18696 5024
rect 18651 4984 18696 5012
rect 16393 4975 16451 4981
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 19702 4972 19708 5024
rect 19760 5012 19766 5024
rect 20088 5012 20116 5052
rect 19760 4984 20116 5012
rect 20165 5015 20223 5021
rect 19760 4972 19766 4984
rect 20165 4981 20177 5015
rect 20211 5012 20223 5015
rect 20438 5012 20444 5024
rect 20211 4984 20444 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 1104 4922 23460 4944
rect 1104 4870 3749 4922
rect 3801 4870 3813 4922
rect 3865 4870 3877 4922
rect 3929 4870 3941 4922
rect 3993 4870 4005 4922
rect 4057 4870 9347 4922
rect 9399 4870 9411 4922
rect 9463 4870 9475 4922
rect 9527 4870 9539 4922
rect 9591 4870 9603 4922
rect 9655 4870 14945 4922
rect 14997 4870 15009 4922
rect 15061 4870 15073 4922
rect 15125 4870 15137 4922
rect 15189 4870 15201 4922
rect 15253 4870 20543 4922
rect 20595 4870 20607 4922
rect 20659 4870 20671 4922
rect 20723 4870 20735 4922
rect 20787 4870 20799 4922
rect 20851 4870 23460 4922
rect 1104 4848 23460 4870
rect 6914 4808 6920 4820
rect 6564 4780 6920 4808
rect 6564 4681 6592 4780
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7101 4811 7159 4817
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 17405 4811 17463 4817
rect 7147 4780 9904 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 7193 4743 7251 4749
rect 7193 4740 7205 4743
rect 6656 4712 7205 4740
rect 6656 4681 6684 4712
rect 7193 4709 7205 4712
rect 7239 4709 7251 4743
rect 7193 4703 7251 4709
rect 7466 4700 7472 4752
rect 7524 4740 7530 4752
rect 8386 4740 8392 4752
rect 7524 4712 8064 4740
rect 7524 4700 7530 4712
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 6641 4675 6699 4681
rect 6641 4641 6653 4675
rect 6687 4641 6699 4675
rect 7650 4672 7656 4684
rect 6641 4635 6699 4641
rect 6840 4644 7656 4672
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6840 4604 6868 4644
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 8036 4681 8064 4712
rect 8220 4712 8392 4740
rect 8220 4681 8248 4712
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4641 8263 4675
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 8205 4635 8263 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 9876 4672 9904 4780
rect 17405 4777 17417 4811
rect 17451 4808 17463 4811
rect 17586 4808 17592 4820
rect 17451 4780 17592 4808
rect 17451 4777 17463 4780
rect 17405 4771 17463 4777
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 19245 4811 19303 4817
rect 19245 4777 19257 4811
rect 19291 4808 19303 4811
rect 19978 4808 19984 4820
rect 19291 4780 19984 4808
rect 19291 4777 19303 4780
rect 19245 4771 19303 4777
rect 19978 4768 19984 4780
rect 20036 4808 20042 4820
rect 21269 4811 21327 4817
rect 20036 4780 20668 4808
rect 20036 4768 20042 4780
rect 20640 4740 20668 4780
rect 21269 4777 21281 4811
rect 21315 4808 21327 4811
rect 21634 4808 21640 4820
rect 21315 4780 21640 4808
rect 21315 4777 21327 4780
rect 21269 4771 21327 4777
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 23290 4740 23296 4752
rect 20640 4712 21312 4740
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9876 4644 9965 4672
rect 9953 4641 9965 4644
rect 9999 4672 10011 4675
rect 10410 4672 10416 4684
rect 9999 4644 10416 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 15470 4632 15476 4684
rect 15528 4672 15534 4684
rect 15565 4675 15623 4681
rect 15565 4672 15577 4675
rect 15528 4644 15577 4672
rect 15528 4632 15534 4644
rect 15565 4641 15577 4644
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 16044 4675 16102 4681
rect 16044 4641 16056 4675
rect 16090 4672 16102 4675
rect 16298 4672 16304 4684
rect 16090 4644 16160 4672
rect 16259 4644 16304 4672
rect 16090 4641 16102 4644
rect 16044 4635 16102 4641
rect 6135 4576 6868 4604
rect 7377 4607 7435 4613
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7423 4576 7604 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 6733 4539 6791 4545
rect 6733 4536 6745 4539
rect 6288 4508 6745 4536
rect 6288 4477 6316 4508
rect 6733 4505 6745 4508
rect 6779 4505 6791 4539
rect 6733 4499 6791 4505
rect 7576 4477 7604 4576
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7800 4576 7941 4604
rect 7800 4564 7806 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 10042 4604 10048 4616
rect 10003 4576 10048 4604
rect 7929 4567 7987 4573
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 16132 4604 16160 4644
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4672 18199 4675
rect 18230 4672 18236 4684
rect 18187 4644 18236 4672
rect 18187 4641 18199 4644
rect 18141 4635 18199 4641
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 18874 4672 18880 4684
rect 18835 4644 18880 4672
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 16132 4576 16979 4604
rect 16951 4536 16979 4576
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 17865 4607 17923 4613
rect 17865 4604 17877 4607
rect 17460 4576 17877 4604
rect 17460 4564 17466 4576
rect 17865 4573 17877 4576
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 20070 4604 20076 4616
rect 18748 4576 20076 4604
rect 18748 4564 18754 4576
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 20180 4576 20637 4604
rect 20180 4548 20208 4576
rect 20625 4573 20637 4576
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 20806 4564 20812 4616
rect 20864 4604 20870 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20864 4576 20913 4604
rect 20864 4564 20870 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 21174 4604 21180 4616
rect 21135 4576 21180 4604
rect 20901 4567 20959 4573
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 21284 4604 21312 4712
rect 21928 4712 23296 4740
rect 21729 4675 21787 4681
rect 21729 4641 21741 4675
rect 21775 4672 21787 4675
rect 21818 4672 21824 4684
rect 21775 4644 21824 4672
rect 21775 4641 21787 4644
rect 21729 4635 21787 4641
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 21928 4681 21956 4712
rect 23290 4700 23296 4712
rect 23348 4700 23354 4752
rect 21913 4675 21971 4681
rect 21913 4641 21925 4675
rect 21959 4641 21971 4675
rect 21913 4635 21971 4641
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 22646 4672 22652 4684
rect 22152 4644 22508 4672
rect 22607 4644 22652 4672
rect 22152 4632 22158 4644
rect 22278 4604 22284 4616
rect 21284 4576 22284 4604
rect 22278 4564 22284 4576
rect 22336 4564 22342 4616
rect 22480 4613 22508 4644
rect 22646 4632 22652 4644
rect 22704 4632 22710 4684
rect 22465 4607 22523 4613
rect 22465 4573 22477 4607
rect 22511 4573 22523 4607
rect 22465 4567 22523 4573
rect 22557 4607 22615 4613
rect 22557 4573 22569 4607
rect 22603 4604 22615 4607
rect 23382 4604 23388 4616
rect 22603 4576 23388 4604
rect 22603 4573 22615 4576
rect 22557 4567 22615 4573
rect 23382 4564 23388 4576
rect 23440 4564 23446 4616
rect 18230 4536 18236 4548
rect 16951 4508 18236 4536
rect 18230 4496 18236 4508
rect 18288 4496 18294 4548
rect 18785 4539 18843 4545
rect 18785 4505 18797 4539
rect 18831 4536 18843 4539
rect 19334 4536 19340 4548
rect 18831 4508 19340 4536
rect 18831 4505 18843 4508
rect 18785 4499 18843 4505
rect 19334 4496 19340 4508
rect 19392 4496 19398 4548
rect 20162 4496 20168 4548
rect 20220 4496 20226 4548
rect 20254 4496 20260 4548
rect 20312 4536 20318 4548
rect 20358 4539 20416 4545
rect 20358 4536 20370 4539
rect 20312 4508 20370 4536
rect 20312 4496 20318 4508
rect 20358 4505 20370 4508
rect 20404 4505 20416 4539
rect 20358 4499 20416 4505
rect 20530 4496 20536 4548
rect 20588 4536 20594 4548
rect 21637 4539 21695 4545
rect 20588 4508 21036 4536
rect 20588 4496 20594 4508
rect 6273 4471 6331 4477
rect 6273 4437 6285 4471
rect 6319 4437 6331 4471
rect 6273 4431 6331 4437
rect 7561 4471 7619 4477
rect 7561 4437 7573 4471
rect 7607 4437 7619 4471
rect 7561 4431 7619 4437
rect 10413 4471 10471 4477
rect 10413 4437 10425 4471
rect 10459 4468 10471 4471
rect 10870 4468 10876 4480
rect 10459 4440 10876 4468
rect 10459 4437 10471 4440
rect 10413 4431 10471 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 16031 4471 16089 4477
rect 16031 4437 16043 4471
rect 16077 4468 16089 4471
rect 16206 4468 16212 4480
rect 16077 4440 16212 4468
rect 16077 4437 16089 4440
rect 16031 4431 16089 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 16632 4440 17509 4468
rect 16632 4428 16638 4440
rect 17497 4437 17509 4440
rect 17543 4437 17555 4471
rect 17497 4431 17555 4437
rect 17957 4471 18015 4477
rect 17957 4437 17969 4471
rect 18003 4468 18015 4471
rect 18325 4471 18383 4477
rect 18325 4468 18337 4471
rect 18003 4440 18337 4468
rect 18003 4437 18015 4440
rect 17957 4431 18015 4437
rect 18325 4437 18337 4440
rect 18371 4437 18383 4471
rect 18690 4468 18696 4480
rect 18651 4440 18696 4468
rect 18325 4431 18383 4437
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 18966 4428 18972 4480
rect 19024 4468 19030 4480
rect 19702 4468 19708 4480
rect 19024 4440 19708 4468
rect 19024 4428 19030 4440
rect 19702 4428 19708 4440
rect 19760 4428 19766 4480
rect 19794 4428 19800 4480
rect 19852 4468 19858 4480
rect 21008 4477 21036 4508
rect 21637 4505 21649 4539
rect 21683 4536 21695 4539
rect 22925 4539 22983 4545
rect 22925 4536 22937 4539
rect 21683 4508 22937 4536
rect 21683 4505 21695 4508
rect 21637 4499 21695 4505
rect 22925 4505 22937 4508
rect 22971 4505 22983 4539
rect 22925 4499 22983 4505
rect 20717 4471 20775 4477
rect 20717 4468 20729 4471
rect 19852 4440 20729 4468
rect 19852 4428 19858 4440
rect 20717 4437 20729 4440
rect 20763 4437 20775 4471
rect 20717 4431 20775 4437
rect 20993 4471 21051 4477
rect 20993 4437 21005 4471
rect 21039 4437 21051 4471
rect 20993 4431 21051 4437
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22152 4440 22197 4468
rect 22152 4428 22158 4440
rect 1104 4378 23460 4400
rect 1104 4326 6548 4378
rect 6600 4326 6612 4378
rect 6664 4326 6676 4378
rect 6728 4326 6740 4378
rect 6792 4326 6804 4378
rect 6856 4326 12146 4378
rect 12198 4326 12210 4378
rect 12262 4326 12274 4378
rect 12326 4326 12338 4378
rect 12390 4326 12402 4378
rect 12454 4326 17744 4378
rect 17796 4326 17808 4378
rect 17860 4326 17872 4378
rect 17924 4326 17936 4378
rect 17988 4326 18000 4378
rect 18052 4326 23460 4378
rect 1104 4304 23460 4326
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7193 4267 7251 4273
rect 7193 4264 7205 4267
rect 6972 4236 7205 4264
rect 6972 4224 6978 4236
rect 7193 4233 7205 4236
rect 7239 4233 7251 4267
rect 7193 4227 7251 4233
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 17865 4267 17923 4273
rect 17865 4264 17877 4267
rect 15988 4236 17877 4264
rect 15988 4224 15994 4236
rect 17865 4233 17877 4236
rect 17911 4233 17923 4267
rect 17865 4227 17923 4233
rect 18690 4224 18696 4276
rect 18748 4264 18754 4276
rect 19153 4267 19211 4273
rect 19153 4264 19165 4267
rect 18748 4236 19165 4264
rect 18748 4224 18754 4236
rect 19153 4233 19165 4236
rect 19199 4233 19211 4267
rect 19794 4264 19800 4276
rect 19755 4236 19800 4264
rect 19153 4227 19211 4233
rect 19794 4224 19800 4236
rect 19852 4224 19858 4276
rect 20438 4224 20444 4276
rect 20496 4264 20502 4276
rect 20717 4267 20775 4273
rect 20717 4264 20729 4267
rect 20496 4236 20729 4264
rect 20496 4224 20502 4236
rect 20717 4233 20729 4236
rect 20763 4233 20775 4267
rect 20717 4227 20775 4233
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 22152 4236 22197 4264
rect 22152 4224 22158 4236
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 14884 4168 15976 4196
rect 14884 4156 14890 4168
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 10870 4128 10876 4140
rect 10831 4100 10876 4128
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 15948 4137 15976 4168
rect 16022 4156 16028 4208
rect 16080 4196 16086 4208
rect 16117 4199 16175 4205
rect 16117 4196 16129 4199
rect 16080 4168 16129 4196
rect 16080 4156 16086 4168
rect 16117 4165 16129 4168
rect 16163 4165 16175 4199
rect 16117 4159 16175 4165
rect 16485 4199 16543 4205
rect 16485 4165 16497 4199
rect 16531 4196 16543 4199
rect 17037 4199 17095 4205
rect 17037 4196 17049 4199
rect 16531 4168 17049 4196
rect 16531 4165 16543 4168
rect 16485 4159 16543 4165
rect 17037 4165 17049 4168
rect 17083 4165 17095 4199
rect 17037 4159 17095 4165
rect 17310 4156 17316 4208
rect 17368 4196 17374 4208
rect 20456 4196 20484 4224
rect 22189 4199 22247 4205
rect 22189 4196 22201 4199
rect 17368 4168 18736 4196
rect 17368 4156 17374 4168
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16356 4100 16896 4128
rect 16356 4088 16362 4100
rect 15654 4020 15660 4072
rect 15712 4060 15718 4072
rect 16390 4060 16396 4072
rect 15712 4032 16396 4060
rect 15712 4020 15718 4032
rect 16390 4020 16396 4032
rect 16448 4060 16454 4072
rect 16448 4032 16620 4060
rect 16448 4020 16454 4032
rect 16114 3952 16120 4004
rect 16172 3992 16178 4004
rect 16298 3992 16304 4004
rect 16172 3964 16304 3992
rect 16172 3952 16178 3964
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11057 3927 11115 3933
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 12526 3924 12532 3936
rect 11103 3896 12532 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 16482 3924 16488 3936
rect 15896 3896 16488 3924
rect 15896 3884 15902 3896
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 16592 3924 16620 4032
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16724 4032 16773 4060
rect 16724 4020 16730 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 16868 3992 16896 4100
rect 16942 4088 16948 4140
rect 17000 4128 17006 4140
rect 17000 4100 17045 4128
rect 17000 4088 17006 4100
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 18708 4137 18736 4168
rect 19352 4168 20484 4196
rect 22112 4168 22201 4196
rect 19352 4137 19380 4168
rect 22112 4140 22140 4168
rect 22189 4165 22201 4168
rect 22235 4165 22247 4199
rect 22189 4159 22247 4165
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17276 4100 17785 4128
rect 17276 4088 17282 4100
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 19337 4131 19395 4137
rect 19337 4097 19349 4131
rect 19383 4097 19395 4131
rect 19337 4091 19395 4097
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 20530 4128 20536 4140
rect 19751 4100 20536 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20625 4131 20683 4137
rect 20625 4097 20637 4131
rect 20671 4097 20683 4131
rect 21266 4128 21272 4140
rect 21227 4100 21272 4128
rect 20625 4091 20683 4097
rect 17034 4020 17040 4072
rect 17092 4060 17098 4072
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 17092 4032 17601 4060
rect 17092 4020 17098 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 18414 4060 18420 4072
rect 18375 4032 18420 4060
rect 17589 4023 17647 4029
rect 18414 4020 18420 4032
rect 18472 4020 18478 4072
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4029 18659 4063
rect 19518 4060 19524 4072
rect 19479 4032 19524 4060
rect 18601 4023 18659 4029
rect 18616 3992 18644 4023
rect 19518 4020 19524 4032
rect 19576 4020 19582 4072
rect 20438 4060 20444 4072
rect 20180 4032 20444 4060
rect 20180 4001 20208 4032
rect 20438 4020 20444 4032
rect 20496 4060 20502 4072
rect 20640 4060 20668 4091
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 21358 4088 21364 4140
rect 21416 4128 21422 4140
rect 21416 4100 21461 4128
rect 21416 4088 21422 4100
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 22833 4131 22891 4137
rect 22833 4097 22845 4131
rect 22879 4128 22891 4131
rect 23566 4128 23572 4140
rect 22879 4100 23572 4128
rect 22879 4097 22891 4100
rect 22833 4091 22891 4097
rect 23566 4088 23572 4100
rect 23624 4088 23630 4140
rect 20496 4032 20668 4060
rect 20901 4063 20959 4069
rect 20496 4020 20502 4032
rect 20901 4029 20913 4063
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22738 4060 22744 4072
rect 22051 4032 22744 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 16868 3964 18644 3992
rect 20165 3995 20223 4001
rect 20165 3961 20177 3995
rect 20211 3961 20223 3995
rect 20916 3992 20944 4023
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 23750 4060 23756 4072
rect 22848 4032 23756 4060
rect 21085 3995 21143 4001
rect 21085 3992 21097 3995
rect 20916 3964 21097 3992
rect 20165 3955 20223 3961
rect 21085 3961 21097 3964
rect 21131 3961 21143 3995
rect 21085 3955 21143 3961
rect 21358 3952 21364 4004
rect 21416 3992 21422 4004
rect 22848 3992 22876 4032
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 21416 3964 22876 3992
rect 23017 3995 23075 4001
rect 21416 3952 21422 3964
rect 23017 3961 23029 3995
rect 23063 3992 23075 3995
rect 23198 3992 23204 4004
rect 23063 3964 23204 3992
rect 23063 3961 23075 3964
rect 23017 3955 23075 3961
rect 23198 3952 23204 3964
rect 23256 3952 23262 4004
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 16592 3896 17417 3924
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17405 3887 17463 3893
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 18104 3896 18245 3924
rect 18104 3884 18110 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3924 19119 3927
rect 19978 3924 19984 3936
rect 19107 3896 19984 3924
rect 19107 3893 19119 3896
rect 19061 3887 19119 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 21542 3924 21548 3936
rect 20312 3896 20357 3924
rect 21503 3896 21548 3924
rect 20312 3884 20318 3896
rect 21542 3884 21548 3896
rect 21600 3884 21606 3936
rect 22462 3884 22468 3936
rect 22520 3924 22526 3936
rect 22557 3927 22615 3933
rect 22557 3924 22569 3927
rect 22520 3896 22569 3924
rect 22520 3884 22526 3896
rect 22557 3893 22569 3896
rect 22603 3893 22615 3927
rect 22557 3887 22615 3893
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 22704 3896 22749 3924
rect 22704 3884 22710 3896
rect 1104 3834 23460 3856
rect 1104 3782 3749 3834
rect 3801 3782 3813 3834
rect 3865 3782 3877 3834
rect 3929 3782 3941 3834
rect 3993 3782 4005 3834
rect 4057 3782 9347 3834
rect 9399 3782 9411 3834
rect 9463 3782 9475 3834
rect 9527 3782 9539 3834
rect 9591 3782 9603 3834
rect 9655 3782 14945 3834
rect 14997 3782 15009 3834
rect 15061 3782 15073 3834
rect 15125 3782 15137 3834
rect 15189 3782 15201 3834
rect 15253 3782 20543 3834
rect 20595 3782 20607 3834
rect 20659 3782 20671 3834
rect 20723 3782 20735 3834
rect 20787 3782 20799 3834
rect 20851 3782 23460 3834
rect 1104 3760 23460 3782
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 17218 3720 17224 3732
rect 9824 3692 16804 3720
rect 17179 3692 17224 3720
rect 9824 3680 9830 3692
rect 12894 3652 12900 3664
rect 12360 3624 12900 3652
rect 12360 3593 12388 3624
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 16776 3652 16804 3692
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 19334 3720 19340 3732
rect 19295 3692 19340 3720
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 19613 3723 19671 3729
rect 19613 3720 19625 3723
rect 19444 3692 19625 3720
rect 19444 3652 19472 3692
rect 19613 3689 19625 3692
rect 19659 3689 19671 3723
rect 19613 3683 19671 3689
rect 20070 3680 20076 3732
rect 20128 3720 20134 3732
rect 20625 3723 20683 3729
rect 20128 3692 20392 3720
rect 20128 3680 20134 3692
rect 20254 3652 20260 3664
rect 16776 3624 19472 3652
rect 19536 3624 20260 3652
rect 12345 3587 12403 3593
rect 12345 3553 12357 3587
rect 12391 3553 12403 3587
rect 12526 3584 12532 3596
rect 12487 3556 12532 3584
rect 12345 3547 12403 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 15844 3587 15902 3593
rect 15844 3584 15856 3587
rect 14424 3556 15856 3584
rect 14424 3544 14430 3556
rect 15844 3553 15856 3556
rect 15890 3584 15902 3587
rect 15930 3584 15936 3596
rect 15890 3556 15936 3584
rect 15890 3553 15902 3556
rect 15844 3547 15902 3553
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 16540 3556 17877 3584
rect 16540 3544 16546 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 18046 3584 18052 3596
rect 18007 3556 18052 3584
rect 17865 3547 17923 3553
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 18138 3544 18144 3596
rect 18196 3584 18202 3596
rect 19150 3584 19156 3596
rect 18196 3556 19156 3584
rect 18196 3544 18202 3556
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 5074 3516 5080 3528
rect 1627 3488 5080 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 10652 3488 12633 3516
rect 10652 3476 10658 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 15470 3516 15476 3528
rect 15427 3488 15476 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 16080 3488 17601 3516
rect 16080 3476 16086 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18969 3519 19027 3525
rect 18380 3488 18828 3516
rect 18380 3476 18386 3488
rect 18141 3451 18199 3457
rect 18141 3417 18153 3451
rect 18187 3448 18199 3451
rect 18601 3451 18659 3457
rect 18601 3448 18613 3451
rect 18187 3420 18613 3448
rect 18187 3417 18199 3420
rect 18141 3411 18199 3417
rect 18601 3417 18613 3420
rect 18647 3417 18659 3451
rect 18800 3448 18828 3488
rect 18969 3485 18981 3519
rect 19015 3516 19027 3519
rect 19334 3516 19340 3528
rect 19015 3488 19340 3516
rect 19015 3485 19027 3488
rect 18969 3479 19027 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19536 3525 19564 3624
rect 20254 3612 20260 3624
rect 20312 3612 20318 3664
rect 20364 3652 20392 3692
rect 20625 3689 20637 3723
rect 20671 3720 20683 3723
rect 21358 3720 21364 3732
rect 20671 3692 21364 3720
rect 20671 3689 20683 3692
rect 20625 3683 20683 3689
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 22370 3680 22376 3732
rect 22428 3720 22434 3732
rect 22557 3723 22615 3729
rect 22557 3720 22569 3723
rect 22428 3692 22569 3720
rect 22428 3680 22434 3692
rect 22557 3689 22569 3692
rect 22603 3689 22615 3723
rect 23014 3720 23020 3732
rect 22975 3692 23020 3720
rect 22557 3683 22615 3689
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 22830 3652 22836 3664
rect 20364 3624 21496 3652
rect 19702 3544 19708 3596
rect 19760 3584 19766 3596
rect 19981 3587 20039 3593
rect 19981 3584 19993 3587
rect 19760 3556 19993 3584
rect 19760 3544 19766 3556
rect 19981 3553 19993 3556
rect 20027 3553 20039 3587
rect 21082 3584 21088 3596
rect 19981 3547 20039 3553
rect 20088 3556 21088 3584
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3516 19855 3519
rect 20088 3516 20116 3556
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 21468 3593 21496 3624
rect 22572 3624 22836 3652
rect 21453 3587 21511 3593
rect 21453 3553 21465 3587
rect 21499 3553 21511 3587
rect 22278 3584 22284 3596
rect 22239 3556 22284 3584
rect 21453 3547 21511 3553
rect 22278 3544 22284 3556
rect 22336 3544 22342 3596
rect 19843 3488 20116 3516
rect 19843 3485 19855 3488
rect 19797 3479 19855 3485
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 20220 3488 20729 3516
rect 20220 3476 20226 3488
rect 20717 3485 20729 3488
rect 20763 3485 20775 3519
rect 20717 3479 20775 3485
rect 20898 3476 20904 3528
rect 20956 3516 20962 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20956 3488 21281 3516
rect 20956 3476 20962 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 22189 3519 22247 3525
rect 22189 3485 22201 3519
rect 22235 3516 22247 3519
rect 22572 3516 22600 3624
rect 22830 3612 22836 3624
rect 22888 3612 22894 3664
rect 22738 3516 22744 3528
rect 22235 3488 22600 3516
rect 22699 3488 22744 3516
rect 22235 3485 22247 3488
rect 22189 3479 22247 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 21082 3448 21088 3460
rect 18800 3420 21088 3448
rect 18601 3411 18659 3417
rect 21082 3408 21088 3420
rect 21140 3408 21146 3460
rect 22278 3408 22284 3460
rect 22336 3448 22342 3460
rect 22462 3448 22468 3460
rect 22336 3420 22468 3448
rect 22336 3408 22342 3420
rect 22462 3408 22468 3420
rect 22520 3448 22526 3460
rect 22848 3448 22876 3479
rect 22520 3420 22876 3448
rect 22520 3408 22526 3420
rect 1394 3380 1400 3392
rect 1355 3352 1400 3380
rect 1394 3340 1400 3352
rect 1452 3340 1458 3392
rect 12986 3380 12992 3392
rect 12947 3352 12992 3380
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 15847 3383 15905 3389
rect 15847 3349 15859 3383
rect 15893 3380 15905 3383
rect 16206 3380 16212 3392
rect 15893 3352 16212 3380
rect 15893 3349 15905 3352
rect 15847 3343 15905 3349
rect 16206 3340 16212 3352
rect 16264 3340 16270 3392
rect 17310 3340 17316 3392
rect 17368 3380 17374 3392
rect 18506 3380 18512 3392
rect 17368 3352 17413 3380
rect 18467 3352 18512 3380
rect 17368 3340 17374 3352
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 19150 3340 19156 3392
rect 19208 3380 19214 3392
rect 20165 3383 20223 3389
rect 20165 3380 20177 3383
rect 19208 3352 20177 3380
rect 19208 3340 19214 3352
rect 20165 3349 20177 3352
rect 20211 3349 20223 3383
rect 20165 3343 20223 3349
rect 20257 3383 20315 3389
rect 20257 3349 20269 3383
rect 20303 3380 20315 3383
rect 20438 3380 20444 3392
rect 20303 3352 20444 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 20901 3383 20959 3389
rect 20901 3349 20913 3383
rect 20947 3380 20959 3383
rect 21266 3380 21272 3392
rect 20947 3352 21272 3380
rect 20947 3349 20959 3352
rect 20901 3343 20959 3349
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 21361 3383 21419 3389
rect 21361 3349 21373 3383
rect 21407 3380 21419 3383
rect 21729 3383 21787 3389
rect 21729 3380 21741 3383
rect 21407 3352 21741 3380
rect 21407 3349 21419 3352
rect 21361 3343 21419 3349
rect 21729 3349 21741 3352
rect 21775 3349 21787 3383
rect 21729 3343 21787 3349
rect 22097 3383 22155 3389
rect 22097 3349 22109 3383
rect 22143 3380 22155 3383
rect 22554 3380 22560 3392
rect 22143 3352 22560 3380
rect 22143 3349 22155 3352
rect 22097 3343 22155 3349
rect 22554 3340 22560 3352
rect 22612 3340 22618 3392
rect 1104 3290 23460 3312
rect 1104 3238 6548 3290
rect 6600 3238 6612 3290
rect 6664 3238 6676 3290
rect 6728 3238 6740 3290
rect 6792 3238 6804 3290
rect 6856 3238 12146 3290
rect 12198 3238 12210 3290
rect 12262 3238 12274 3290
rect 12326 3238 12338 3290
rect 12390 3238 12402 3290
rect 12454 3238 17744 3290
rect 17796 3238 17808 3290
rect 17860 3238 17872 3290
rect 17924 3238 17936 3290
rect 17988 3238 18000 3290
rect 18052 3238 23460 3290
rect 1104 3216 23460 3238
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 16945 3179 17003 3185
rect 16945 3176 16957 3179
rect 13044 3148 16957 3176
rect 13044 3136 13050 3148
rect 16945 3145 16957 3148
rect 16991 3145 17003 3179
rect 16945 3139 17003 3145
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 17310 3176 17316 3188
rect 17083 3148 17316 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 17310 3136 17316 3148
rect 17368 3136 17374 3188
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 18325 3179 18383 3185
rect 17460 3148 17505 3176
rect 17460 3136 17466 3148
rect 18325 3145 18337 3179
rect 18371 3176 18383 3179
rect 18785 3179 18843 3185
rect 18785 3176 18797 3179
rect 18371 3148 18797 3176
rect 18371 3145 18383 3148
rect 18325 3139 18383 3145
rect 18785 3145 18797 3148
rect 18831 3176 18843 3179
rect 20346 3176 20352 3188
rect 18831 3148 20352 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 5074 3068 5080 3120
rect 5132 3108 5138 3120
rect 17865 3111 17923 3117
rect 17865 3108 17877 3111
rect 5132 3080 17877 3108
rect 5132 3068 5138 3080
rect 17865 3077 17877 3080
rect 17911 3077 17923 3111
rect 17865 3071 17923 3077
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6595 3012 6776 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 4522 2796 4528 2848
rect 4580 2836 4586 2848
rect 6748 2845 6776 3012
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 18141 3043 18199 3049
rect 11112 3012 18092 3040
rect 11112 3000 11118 3012
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 18064 2972 18092 3012
rect 18141 3009 18153 3043
rect 18187 3040 18199 3043
rect 18340 3040 18368 3139
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 21361 3179 21419 3185
rect 21361 3176 21373 3179
rect 20496 3148 21373 3176
rect 20496 3136 20502 3148
rect 21361 3145 21373 3148
rect 21407 3145 21419 3179
rect 21361 3139 21419 3145
rect 23017 3179 23075 3185
rect 23017 3145 23029 3179
rect 23063 3176 23075 3179
rect 23106 3176 23112 3188
rect 23063 3148 23112 3176
rect 23063 3145 23075 3148
rect 23017 3139 23075 3145
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19794 3108 19800 3120
rect 19484 3080 19800 3108
rect 19484 3068 19490 3080
rect 19794 3068 19800 3080
rect 19852 3068 19858 3120
rect 20533 3111 20591 3117
rect 20533 3077 20545 3111
rect 20579 3108 20591 3111
rect 21821 3111 21879 3117
rect 21821 3108 21833 3111
rect 20579 3080 21833 3108
rect 20579 3077 20591 3080
rect 20533 3071 20591 3077
rect 21821 3077 21833 3080
rect 21867 3077 21879 3111
rect 21821 3071 21879 3077
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18187 3012 18368 3040
rect 18708 3012 19257 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 18708 2972 18736 3012
rect 19245 3009 19257 3012
rect 19291 3040 19303 3043
rect 19518 3040 19524 3052
rect 19291 3012 19524 3040
rect 19291 3009 19303 3012
rect 19245 3003 19303 3009
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20625 3043 20683 3049
rect 20625 3040 20637 3043
rect 20036 3012 20637 3040
rect 20036 3000 20042 3012
rect 20625 3009 20637 3012
rect 20671 3009 20683 3043
rect 20625 3003 20683 3009
rect 20898 3000 20904 3052
rect 20956 3040 20962 3052
rect 21174 3040 21180 3052
rect 20956 3012 21180 3040
rect 20956 3000 20962 3012
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3009 21327 3043
rect 22646 3040 22652 3052
rect 22607 3012 22652 3040
rect 21269 3003 21327 3009
rect 18064 2944 18736 2972
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2972 19119 2975
rect 19334 2972 19340 2984
rect 19107 2944 19340 2972
rect 19107 2941 19119 2944
rect 19061 2935 19119 2941
rect 19334 2932 19340 2944
rect 19392 2972 19398 2984
rect 19705 2975 19763 2981
rect 19705 2972 19717 2975
rect 19392 2944 19717 2972
rect 19392 2932 19398 2944
rect 19705 2941 19717 2944
rect 19751 2972 19763 2975
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19751 2944 20085 2972
rect 19751 2941 19763 2944
rect 19705 2935 19763 2941
rect 20073 2941 20085 2944
rect 20119 2972 20131 2975
rect 20162 2972 20168 2984
rect 20119 2944 20168 2972
rect 20119 2941 20131 2944
rect 20073 2935 20131 2941
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 20717 2975 20775 2981
rect 20717 2972 20729 2975
rect 20272 2944 20729 2972
rect 16390 2864 16396 2916
rect 16448 2904 16454 2916
rect 19426 2904 19432 2916
rect 16448 2876 19432 2904
rect 16448 2864 16454 2876
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 19518 2864 19524 2916
rect 19576 2904 19582 2916
rect 19576 2876 19621 2904
rect 19576 2864 19582 2876
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 20272 2904 20300 2944
rect 20717 2941 20729 2944
rect 20763 2941 20775 2975
rect 20717 2935 20775 2941
rect 19944 2876 20300 2904
rect 19944 2864 19950 2876
rect 20530 2864 20536 2916
rect 20588 2904 20594 2916
rect 21284 2904 21312 3003
rect 22646 3000 22652 3012
rect 22704 3000 22710 3052
rect 22738 3000 22744 3052
rect 22796 3040 22802 3052
rect 22833 3043 22891 3049
rect 22833 3040 22845 3043
rect 22796 3012 22845 3040
rect 22796 3000 22802 3012
rect 22833 3009 22845 3012
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 22186 2932 22192 2984
rect 22244 2972 22250 2984
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 22244 2944 22385 2972
rect 22244 2932 22250 2944
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 20588 2876 21312 2904
rect 20588 2864 20594 2876
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 4580 2808 6377 2836
rect 4580 2796 4586 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 6733 2839 6791 2845
rect 6733 2805 6745 2839
rect 6779 2836 6791 2839
rect 10594 2836 10600 2848
rect 6779 2808 10600 2836
rect 6779 2805 6791 2808
rect 6733 2799 6791 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 19334 2836 19340 2848
rect 14240 2808 19340 2836
rect 14240 2796 14246 2808
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20165 2839 20223 2845
rect 20165 2836 20177 2839
rect 20036 2808 20177 2836
rect 20036 2796 20042 2808
rect 20165 2805 20177 2808
rect 20211 2836 20223 2839
rect 20346 2836 20352 2848
rect 20211 2808 20352 2836
rect 20211 2805 20223 2808
rect 20165 2799 20223 2805
rect 20346 2796 20352 2808
rect 20404 2796 20410 2848
rect 21082 2836 21088 2848
rect 21043 2808 21088 2836
rect 21082 2796 21088 2808
rect 21140 2796 21146 2848
rect 1104 2746 23460 2768
rect 1104 2694 3749 2746
rect 3801 2694 3813 2746
rect 3865 2694 3877 2746
rect 3929 2694 3941 2746
rect 3993 2694 4005 2746
rect 4057 2694 9347 2746
rect 9399 2694 9411 2746
rect 9463 2694 9475 2746
rect 9527 2694 9539 2746
rect 9591 2694 9603 2746
rect 9655 2694 14945 2746
rect 14997 2694 15009 2746
rect 15061 2694 15073 2746
rect 15125 2694 15137 2746
rect 15189 2694 15201 2746
rect 15253 2694 20543 2746
rect 20595 2694 20607 2746
rect 20659 2694 20671 2746
rect 20723 2694 20735 2746
rect 20787 2694 20799 2746
rect 20851 2694 23460 2746
rect 1104 2672 23460 2694
rect 19334 2632 19340 2644
rect 19295 2604 19340 2632
rect 19334 2592 19340 2604
rect 19392 2632 19398 2644
rect 19978 2632 19984 2644
rect 19392 2604 19984 2632
rect 19392 2592 19398 2604
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20162 2632 20168 2644
rect 20123 2604 20168 2632
rect 20162 2592 20168 2604
rect 20220 2632 20226 2644
rect 20349 2635 20407 2641
rect 20349 2632 20361 2635
rect 20220 2604 20361 2632
rect 20220 2592 20226 2604
rect 20349 2601 20361 2604
rect 20395 2601 20407 2635
rect 20349 2595 20407 2601
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 19797 2567 19855 2573
rect 19797 2564 19809 2567
rect 19300 2536 19809 2564
rect 19300 2524 19306 2536
rect 19797 2533 19809 2536
rect 19843 2533 19855 2567
rect 20364 2564 20392 2595
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 20533 2635 20591 2641
rect 20533 2632 20545 2635
rect 20496 2604 20545 2632
rect 20496 2592 20502 2604
rect 20533 2601 20545 2604
rect 20579 2632 20591 2635
rect 22646 2632 22652 2644
rect 20579 2604 22652 2632
rect 20579 2601 20591 2604
rect 20533 2595 20591 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 23014 2632 23020 2644
rect 22975 2604 23020 2632
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 20717 2567 20775 2573
rect 20717 2564 20729 2567
rect 20364 2536 20729 2564
rect 19797 2527 19855 2533
rect 20717 2533 20729 2536
rect 20763 2564 20775 2567
rect 20901 2567 20959 2573
rect 20901 2564 20913 2567
rect 20763 2536 20913 2564
rect 20763 2533 20775 2536
rect 20717 2527 20775 2533
rect 20901 2533 20913 2536
rect 20947 2564 20959 2567
rect 21085 2567 21143 2573
rect 21085 2564 21097 2567
rect 20947 2536 21097 2564
rect 20947 2533 20959 2536
rect 20901 2527 20959 2533
rect 21085 2533 21097 2536
rect 21131 2564 21143 2567
rect 21545 2567 21603 2573
rect 21545 2564 21557 2567
rect 21131 2536 21557 2564
rect 21131 2533 21143 2536
rect 21085 2527 21143 2533
rect 21545 2533 21557 2536
rect 21591 2533 21603 2567
rect 21545 2527 21603 2533
rect 21652 2536 22416 2564
rect 19518 2496 19524 2508
rect 19431 2468 19524 2496
rect 19518 2456 19524 2468
rect 19576 2496 19582 2508
rect 21652 2496 21680 2536
rect 19576 2468 21680 2496
rect 19576 2456 19582 2468
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22388 2496 22416 2536
rect 22462 2524 22468 2576
rect 22520 2564 22526 2576
rect 23842 2564 23848 2576
rect 22520 2536 23848 2564
rect 22520 2524 22526 2536
rect 23842 2524 23848 2536
rect 23900 2524 23906 2576
rect 22738 2496 22744 2508
rect 22152 2468 22197 2496
rect 22388 2468 22744 2496
rect 22152 2456 22158 2468
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 4522 2428 4528 2440
rect 2547 2400 4528 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 6178 2388 6184 2440
rect 6236 2428 6242 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6236 2400 6377 2428
rect 6236 2388 6242 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 10594 2428 10600 2440
rect 10507 2400 10600 2428
rect 6365 2391 6423 2397
rect 10594 2388 10600 2400
rect 10652 2428 10658 2440
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 10652 2400 10793 2428
rect 10652 2388 10658 2400
rect 10781 2397 10793 2400
rect 10827 2428 10839 2431
rect 19794 2428 19800 2440
rect 10827 2400 19800 2428
rect 10827 2397 10839 2400
rect 10781 2391 10839 2397
rect 19794 2388 19800 2400
rect 19852 2388 19858 2440
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 20898 2428 20904 2440
rect 20119 2400 20904 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20898 2388 20904 2400
rect 20956 2388 20962 2440
rect 21361 2431 21419 2437
rect 21361 2397 21373 2431
rect 21407 2428 21419 2431
rect 22002 2428 22008 2440
rect 21407 2400 22008 2428
rect 21407 2397 21419 2400
rect 21361 2391 21419 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22186 2428 22192 2440
rect 22147 2400 22192 2428
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 22462 2428 22468 2440
rect 22423 2400 22468 2428
rect 22462 2388 22468 2400
rect 22520 2388 22526 2440
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 19628 2332 20300 2360
rect 2130 2252 2136 2304
rect 2188 2292 2194 2304
rect 2317 2295 2375 2301
rect 2317 2292 2329 2295
rect 2188 2264 2329 2292
rect 2188 2252 2194 2264
rect 2317 2261 2329 2264
rect 2363 2261 2375 2295
rect 2317 2255 2375 2261
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 10284 2264 10425 2292
rect 10284 2252 10290 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 19628 2301 19656 2332
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 15528 2264 19625 2292
rect 15528 2252 15534 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 20272 2292 20300 2332
rect 20346 2320 20352 2372
rect 20404 2360 20410 2372
rect 22848 2360 22876 2391
rect 20404 2332 22876 2360
rect 20404 2320 20410 2332
rect 22186 2292 22192 2304
rect 20272 2264 22192 2292
rect 19613 2255 19671 2261
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 22370 2292 22376 2304
rect 22331 2264 22376 2292
rect 22370 2252 22376 2264
rect 22428 2252 22434 2304
rect 22646 2292 22652 2304
rect 22607 2264 22652 2292
rect 22646 2252 22652 2264
rect 22704 2252 22710 2304
rect 1104 2202 23460 2224
rect 1104 2150 6548 2202
rect 6600 2150 6612 2202
rect 6664 2150 6676 2202
rect 6728 2150 6740 2202
rect 6792 2150 6804 2202
rect 6856 2150 12146 2202
rect 12198 2150 12210 2202
rect 12262 2150 12274 2202
rect 12326 2150 12338 2202
rect 12390 2150 12402 2202
rect 12454 2150 17744 2202
rect 17796 2150 17808 2202
rect 17860 2150 17872 2202
rect 17924 2150 17936 2202
rect 17988 2150 18000 2202
rect 18052 2150 23460 2202
rect 1104 2128 23460 2150
<< via1 >>
rect 4068 22720 4120 22772
rect 5448 22720 5500 22772
rect 6184 22720 6236 22772
rect 9312 22720 9364 22772
rect 11428 22720 11480 22772
rect 11888 22720 11940 22772
rect 3608 22652 3660 22704
rect 12164 22652 12216 22704
rect 4988 22584 5040 22636
rect 14372 22584 14424 22636
rect 19616 22584 19668 22636
rect 22008 22584 22060 22636
rect 4620 22516 4672 22568
rect 6736 22516 6788 22568
rect 7196 22516 7248 22568
rect 5540 22448 5592 22500
rect 8668 22448 8720 22500
rect 10876 22448 10928 22500
rect 11520 22448 11572 22500
rect 12532 22448 12584 22500
rect 12716 22448 12768 22500
rect 18328 22448 18380 22500
rect 21456 22448 21508 22500
rect 5448 22380 5500 22432
rect 8024 22380 8076 22432
rect 12164 22380 12216 22432
rect 14004 22380 14056 22432
rect 14096 22380 14148 22432
rect 18144 22380 18196 22432
rect 3749 22278 3801 22330
rect 3813 22278 3865 22330
rect 3877 22278 3929 22330
rect 3941 22278 3993 22330
rect 4005 22278 4057 22330
rect 9347 22278 9399 22330
rect 9411 22278 9463 22330
rect 9475 22278 9527 22330
rect 9539 22278 9591 22330
rect 9603 22278 9655 22330
rect 14945 22278 14997 22330
rect 15009 22278 15061 22330
rect 15073 22278 15125 22330
rect 15137 22278 15189 22330
rect 15201 22278 15253 22330
rect 20543 22278 20595 22330
rect 20607 22278 20659 22330
rect 20671 22278 20723 22330
rect 20735 22278 20787 22330
rect 20799 22278 20851 22330
rect 5356 22219 5408 22228
rect 5356 22185 5365 22219
rect 5365 22185 5399 22219
rect 5399 22185 5408 22219
rect 5356 22176 5408 22185
rect 2320 22040 2372 22092
rect 5172 22108 5224 22160
rect 5264 22108 5316 22160
rect 3148 22040 3200 22092
rect 9036 22108 9088 22160
rect 2596 22015 2648 22024
rect 2596 21981 2605 22015
rect 2605 21981 2639 22015
rect 2639 21981 2648 22015
rect 2596 21972 2648 21981
rect 3056 21972 3108 22024
rect 3240 22015 3292 22024
rect 3240 21981 3249 22015
rect 3249 21981 3283 22015
rect 3283 21981 3292 22015
rect 3240 21972 3292 21981
rect 3608 22015 3660 22024
rect 3608 21981 3617 22015
rect 3617 21981 3651 22015
rect 3651 21981 3660 22015
rect 3608 21972 3660 21981
rect 4068 22015 4120 22024
rect 4068 21981 4070 22015
rect 4070 21981 4104 22015
rect 4104 21981 4120 22015
rect 4068 21972 4120 21981
rect 4344 21972 4396 22024
rect 4620 22015 4672 22024
rect 4620 21981 4629 22015
rect 4629 21981 4663 22015
rect 4663 21981 4672 22015
rect 4620 21972 4672 21981
rect 4804 21972 4856 22024
rect 5172 21972 5224 22024
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 5448 21972 5500 21981
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 8760 22040 8812 22092
rect 6184 22015 6236 22024
rect 6184 21981 6185 22015
rect 6185 21981 6219 22015
rect 6219 21981 6236 22015
rect 6184 21972 6236 21981
rect 6368 21972 6420 22024
rect 6736 22015 6788 22024
rect 6736 21981 6745 22015
rect 6745 21981 6779 22015
rect 6779 21981 6788 22015
rect 6736 21972 6788 21981
rect 2688 21904 2740 21956
rect 1584 21836 1636 21888
rect 2228 21836 2280 21888
rect 2872 21836 2924 21888
rect 3424 21879 3476 21888
rect 3424 21845 3433 21879
rect 3433 21845 3467 21879
rect 3467 21845 3476 21879
rect 3424 21836 3476 21845
rect 3608 21836 3660 21888
rect 4160 21836 4212 21888
rect 4712 21836 4764 21888
rect 4896 21836 4948 21888
rect 5632 21879 5684 21888
rect 5632 21845 5641 21879
rect 5641 21845 5675 21879
rect 5675 21845 5684 21879
rect 5632 21836 5684 21845
rect 7380 21904 7432 21956
rect 9128 21972 9180 22024
rect 10968 22176 11020 22228
rect 14372 22176 14424 22228
rect 21640 22176 21692 22228
rect 22008 22219 22060 22228
rect 22008 22185 22017 22219
rect 22017 22185 22051 22219
rect 22051 22185 22060 22219
rect 22008 22176 22060 22185
rect 10232 22083 10284 22092
rect 10232 22049 10241 22083
rect 10241 22049 10275 22083
rect 10275 22049 10284 22083
rect 10232 22040 10284 22049
rect 12072 22083 12124 22092
rect 12072 22049 12081 22083
rect 12081 22049 12115 22083
rect 12115 22049 12124 22083
rect 12072 22040 12124 22049
rect 12164 22083 12216 22092
rect 12164 22049 12173 22083
rect 12173 22049 12207 22083
rect 12207 22049 12216 22083
rect 12164 22040 12216 22049
rect 10876 22015 10928 22024
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 6184 21836 6236 21888
rect 6460 21836 6512 21888
rect 6644 21836 6696 21888
rect 7564 21879 7616 21888
rect 7564 21845 7573 21879
rect 7573 21845 7607 21879
rect 7607 21845 7616 21879
rect 7564 21836 7616 21845
rect 7932 21879 7984 21888
rect 7932 21845 7941 21879
rect 7941 21845 7975 21879
rect 7975 21845 7984 21879
rect 7932 21836 7984 21845
rect 8668 21904 8720 21956
rect 10140 21904 10192 21956
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 13084 21972 13136 22024
rect 14096 22108 14148 22160
rect 14280 22108 14332 22160
rect 13268 21972 13320 22024
rect 13360 21972 13412 22024
rect 15568 22040 15620 22092
rect 16120 22108 16172 22160
rect 18420 22108 18472 22160
rect 20812 22151 20864 22160
rect 20812 22117 20821 22151
rect 20821 22117 20855 22151
rect 20855 22117 20864 22151
rect 20812 22108 20864 22117
rect 17592 22083 17644 22092
rect 17592 22049 17601 22083
rect 17601 22049 17635 22083
rect 17635 22049 17644 22083
rect 17592 22040 17644 22049
rect 18788 22040 18840 22092
rect 19156 22040 19208 22092
rect 20168 22083 20220 22092
rect 20168 22049 20177 22083
rect 20177 22049 20211 22083
rect 20211 22049 20220 22083
rect 20168 22040 20220 22049
rect 21732 22108 21784 22160
rect 22284 22040 22336 22092
rect 8116 21836 8168 21888
rect 8576 21836 8628 21888
rect 9312 21836 9364 21888
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 10416 21879 10468 21888
rect 10416 21845 10425 21879
rect 10425 21845 10459 21879
rect 10459 21845 10468 21879
rect 10416 21836 10468 21845
rect 12624 21947 12676 21956
rect 12624 21913 12633 21947
rect 12633 21913 12667 21947
rect 12667 21913 12676 21947
rect 12624 21904 12676 21913
rect 14464 21972 14516 22024
rect 14648 21972 14700 22024
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15476 21972 15528 21981
rect 16672 21972 16724 22024
rect 18052 21972 18104 22024
rect 21824 22015 21876 22024
rect 15936 21904 15988 21956
rect 17132 21904 17184 21956
rect 17316 21904 17368 21956
rect 18144 21904 18196 21956
rect 19340 21904 19392 21956
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 22100 21972 22152 22024
rect 22560 22015 22612 22024
rect 22560 21981 22569 22015
rect 22569 21981 22603 22015
rect 22603 21981 22612 22015
rect 22560 21972 22612 21981
rect 20628 21904 20680 21956
rect 20904 21904 20956 21956
rect 11336 21879 11388 21888
rect 11336 21845 11345 21879
rect 11345 21845 11379 21879
rect 11379 21845 11388 21879
rect 11336 21836 11388 21845
rect 11704 21836 11756 21888
rect 11980 21879 12032 21888
rect 11980 21845 11989 21879
rect 11989 21845 12023 21879
rect 12023 21845 12032 21879
rect 11980 21836 12032 21845
rect 13084 21879 13136 21888
rect 13084 21845 13093 21879
rect 13093 21845 13127 21879
rect 13127 21845 13136 21879
rect 13084 21836 13136 21845
rect 14740 21836 14792 21888
rect 15108 21836 15160 21888
rect 15660 21879 15712 21888
rect 15660 21845 15669 21879
rect 15669 21845 15703 21879
rect 15703 21845 15712 21879
rect 15660 21836 15712 21845
rect 15844 21836 15896 21888
rect 16304 21836 16356 21888
rect 17224 21836 17276 21888
rect 17408 21879 17460 21888
rect 17408 21845 17417 21879
rect 17417 21845 17451 21879
rect 17451 21845 17460 21879
rect 17408 21836 17460 21845
rect 17500 21836 17552 21888
rect 18236 21879 18288 21888
rect 18236 21845 18245 21879
rect 18245 21845 18279 21879
rect 18279 21845 18288 21879
rect 18236 21836 18288 21845
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 19064 21879 19116 21888
rect 18696 21836 18748 21845
rect 19064 21845 19073 21879
rect 19073 21845 19107 21879
rect 19107 21845 19116 21879
rect 19064 21836 19116 21845
rect 19616 21879 19668 21888
rect 19616 21845 19625 21879
rect 19625 21845 19659 21879
rect 19659 21845 19668 21879
rect 19616 21836 19668 21845
rect 19708 21879 19760 21888
rect 19708 21845 19717 21879
rect 19717 21845 19751 21879
rect 19751 21845 19760 21879
rect 20352 21879 20404 21888
rect 19708 21836 19760 21845
rect 20352 21845 20361 21879
rect 20361 21845 20395 21879
rect 20395 21845 20404 21879
rect 20352 21836 20404 21845
rect 20444 21879 20496 21888
rect 20444 21845 20453 21879
rect 20453 21845 20487 21879
rect 20487 21845 20496 21879
rect 21272 21879 21324 21888
rect 20444 21836 20496 21845
rect 21272 21845 21281 21879
rect 21281 21845 21315 21879
rect 21315 21845 21324 21879
rect 21272 21836 21324 21845
rect 21364 21879 21416 21888
rect 21364 21845 21373 21879
rect 21373 21845 21407 21879
rect 21407 21845 21416 21879
rect 21364 21836 21416 21845
rect 23204 21972 23256 22024
rect 23388 21836 23440 21888
rect 6548 21734 6600 21786
rect 6612 21734 6664 21786
rect 6676 21734 6728 21786
rect 6740 21734 6792 21786
rect 6804 21734 6856 21786
rect 12146 21734 12198 21786
rect 12210 21734 12262 21786
rect 12274 21734 12326 21786
rect 12338 21734 12390 21786
rect 12402 21734 12454 21786
rect 17744 21734 17796 21786
rect 17808 21734 17860 21786
rect 17872 21734 17924 21786
rect 17936 21734 17988 21786
rect 18000 21734 18052 21786
rect 296 21632 348 21684
rect 2688 21632 2740 21684
rect 3240 21632 3292 21684
rect 4068 21632 4120 21684
rect 3148 21564 3200 21616
rect 5448 21632 5500 21684
rect 7564 21632 7616 21684
rect 9312 21632 9364 21684
rect 9404 21675 9456 21684
rect 9404 21641 9413 21675
rect 9413 21641 9447 21675
rect 9447 21641 9456 21675
rect 9404 21632 9456 21641
rect 4712 21564 4764 21616
rect 2320 21539 2372 21548
rect 2320 21505 2329 21539
rect 2329 21505 2363 21539
rect 2363 21505 2372 21539
rect 2320 21496 2372 21505
rect 2688 21496 2740 21548
rect 3056 21539 3108 21548
rect 3056 21505 3065 21539
rect 3065 21505 3099 21539
rect 3099 21505 3108 21539
rect 3056 21496 3108 21505
rect 3240 21496 3292 21548
rect 2872 21428 2924 21480
rect 3516 21496 3568 21548
rect 3792 21539 3844 21548
rect 3792 21505 3801 21539
rect 3801 21505 3835 21539
rect 3835 21505 3844 21539
rect 3792 21496 3844 21505
rect 3976 21496 4028 21548
rect 4528 21539 4580 21548
rect 4528 21505 4537 21539
rect 4537 21505 4571 21539
rect 4571 21505 4580 21539
rect 4528 21496 4580 21505
rect 940 21360 992 21412
rect 2596 21360 2648 21412
rect 4160 21428 4212 21480
rect 4988 21496 5040 21548
rect 4896 21428 4948 21480
rect 5448 21496 5500 21548
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 10232 21632 10284 21684
rect 10508 21632 10560 21684
rect 12072 21632 12124 21684
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 6092 21428 6144 21480
rect 4436 21360 4488 21412
rect 4804 21403 4856 21412
rect 4804 21369 4813 21403
rect 4813 21369 4847 21403
rect 4847 21369 4856 21403
rect 4804 21360 4856 21369
rect 5172 21403 5224 21412
rect 5172 21369 5181 21403
rect 5181 21369 5215 21403
rect 5215 21369 5224 21403
rect 5172 21360 5224 21369
rect 5356 21360 5408 21412
rect 6000 21360 6052 21412
rect 6460 21360 6512 21412
rect 6644 21403 6696 21412
rect 6644 21369 6653 21403
rect 6653 21369 6687 21403
rect 6687 21369 6696 21403
rect 6644 21360 6696 21369
rect 2504 21292 2556 21344
rect 3884 21292 3936 21344
rect 4068 21292 4120 21344
rect 4252 21335 4304 21344
rect 4252 21301 4261 21335
rect 4261 21301 4295 21335
rect 4295 21301 4304 21335
rect 4252 21292 4304 21301
rect 4344 21292 4396 21344
rect 4988 21292 5040 21344
rect 5264 21292 5316 21344
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 5540 21292 5592 21344
rect 7288 21428 7340 21480
rect 7564 21471 7616 21480
rect 7564 21437 7573 21471
rect 7573 21437 7607 21471
rect 7607 21437 7616 21471
rect 8024 21496 8076 21548
rect 8208 21539 8260 21548
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 11152 21564 11204 21616
rect 13912 21632 13964 21684
rect 12532 21564 12584 21616
rect 12716 21564 12768 21616
rect 15660 21632 15712 21684
rect 16304 21632 16356 21684
rect 17500 21632 17552 21684
rect 18328 21632 18380 21684
rect 19064 21632 19116 21684
rect 7564 21428 7616 21437
rect 8116 21471 8168 21480
rect 8116 21437 8125 21471
rect 8125 21437 8159 21471
rect 8159 21437 8168 21471
rect 8116 21428 8168 21437
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 10692 21496 10744 21548
rect 11612 21496 11664 21548
rect 9496 21471 9548 21480
rect 9496 21437 9505 21471
rect 9505 21437 9539 21471
rect 9539 21437 9548 21471
rect 9496 21428 9548 21437
rect 9864 21428 9916 21480
rect 10324 21428 10376 21480
rect 10416 21428 10468 21480
rect 11796 21428 11848 21480
rect 12900 21428 12952 21480
rect 14464 21496 14516 21548
rect 13268 21428 13320 21480
rect 13452 21471 13504 21480
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 14372 21428 14424 21480
rect 14740 21471 14792 21480
rect 14740 21437 14749 21471
rect 14749 21437 14783 21471
rect 14783 21437 14792 21471
rect 14740 21428 14792 21437
rect 7012 21335 7064 21344
rect 7012 21301 7021 21335
rect 7021 21301 7055 21335
rect 7055 21301 7064 21335
rect 7012 21292 7064 21301
rect 8116 21292 8168 21344
rect 9680 21292 9732 21344
rect 11060 21292 11112 21344
rect 12072 21292 12124 21344
rect 12716 21292 12768 21344
rect 16120 21496 16172 21548
rect 16856 21564 16908 21616
rect 19800 21632 19852 21684
rect 20444 21632 20496 21684
rect 20812 21632 20864 21684
rect 21364 21632 21416 21684
rect 21548 21632 21600 21684
rect 21916 21564 21968 21616
rect 22836 21632 22888 21684
rect 15844 21471 15896 21480
rect 15844 21437 15853 21471
rect 15853 21437 15887 21471
rect 15887 21437 15896 21471
rect 15844 21428 15896 21437
rect 16580 21428 16632 21480
rect 17040 21496 17092 21548
rect 18144 21539 18196 21548
rect 18144 21505 18153 21539
rect 18153 21505 18187 21539
rect 18187 21505 18196 21539
rect 18144 21496 18196 21505
rect 18052 21428 18104 21480
rect 18512 21496 18564 21548
rect 19248 21496 19300 21548
rect 19340 21496 19392 21548
rect 21364 21539 21416 21548
rect 21364 21505 21373 21539
rect 21373 21505 21407 21539
rect 21407 21505 21416 21539
rect 21364 21496 21416 21505
rect 21456 21496 21508 21548
rect 18420 21428 18472 21480
rect 19892 21428 19944 21480
rect 19984 21428 20036 21480
rect 15568 21335 15620 21344
rect 15568 21301 15577 21335
rect 15577 21301 15611 21335
rect 15611 21301 15620 21335
rect 15568 21292 15620 21301
rect 16304 21292 16356 21344
rect 16488 21292 16540 21344
rect 18236 21292 18288 21344
rect 18420 21292 18472 21344
rect 21088 21428 21140 21480
rect 22192 21496 22244 21548
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 22744 21496 22796 21548
rect 20720 21360 20772 21412
rect 20812 21292 20864 21344
rect 23020 21335 23072 21344
rect 23020 21301 23029 21335
rect 23029 21301 23063 21335
rect 23063 21301 23072 21335
rect 23020 21292 23072 21301
rect 3749 21190 3801 21242
rect 3813 21190 3865 21242
rect 3877 21190 3929 21242
rect 3941 21190 3993 21242
rect 4005 21190 4057 21242
rect 9347 21190 9399 21242
rect 9411 21190 9463 21242
rect 9475 21190 9527 21242
rect 9539 21190 9591 21242
rect 9603 21190 9655 21242
rect 14945 21190 14997 21242
rect 15009 21190 15061 21242
rect 15073 21190 15125 21242
rect 15137 21190 15189 21242
rect 15201 21190 15253 21242
rect 20543 21190 20595 21242
rect 20607 21190 20659 21242
rect 20671 21190 20723 21242
rect 20735 21190 20787 21242
rect 20799 21190 20851 21242
rect 2504 21131 2556 21140
rect 2504 21097 2513 21131
rect 2513 21097 2547 21131
rect 2547 21097 2556 21131
rect 2504 21088 2556 21097
rect 2780 21131 2832 21140
rect 2780 21097 2789 21131
rect 2789 21097 2823 21131
rect 2823 21097 2832 21131
rect 2780 21088 2832 21097
rect 3240 21088 3292 21140
rect 5724 21088 5776 21140
rect 7380 21088 7432 21140
rect 7932 21088 7984 21140
rect 3792 21020 3844 21072
rect 6828 21020 6880 21072
rect 3148 20952 3200 21004
rect 5540 20952 5592 21004
rect 2044 20927 2096 20936
rect 2044 20893 2053 20927
rect 2053 20893 2087 20927
rect 2087 20893 2096 20927
rect 2044 20884 2096 20893
rect 3056 20884 3108 20936
rect 3424 20884 3476 20936
rect 3608 20927 3660 20936
rect 3608 20893 3617 20927
rect 3617 20893 3651 20927
rect 3651 20893 3660 20927
rect 3608 20884 3660 20893
rect 3700 20884 3752 20936
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4988 20884 5040 20936
rect 5356 20884 5408 20936
rect 5724 20952 5776 21004
rect 6184 20995 6236 21004
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 7012 20952 7064 21004
rect 8116 20952 8168 21004
rect 8208 20952 8260 21004
rect 8852 21088 8904 21140
rect 9220 21088 9272 21140
rect 9496 21088 9548 21140
rect 11336 21088 11388 21140
rect 10692 21020 10744 21072
rect 13728 21063 13780 21072
rect 13728 21029 13737 21063
rect 13737 21029 13771 21063
rect 13771 21029 13780 21063
rect 13728 21020 13780 21029
rect 13820 21020 13872 21072
rect 14556 21020 14608 21072
rect 15292 21020 15344 21072
rect 9680 20995 9732 21004
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9680 20952 9732 20961
rect 11704 20952 11756 21004
rect 12992 20952 13044 21004
rect 6460 20927 6512 20936
rect 6460 20893 6469 20927
rect 6469 20893 6503 20927
rect 6503 20893 6512 20927
rect 6460 20884 6512 20893
rect 6552 20884 6604 20936
rect 6828 20884 6880 20936
rect 2964 20816 3016 20868
rect 2780 20748 2832 20800
rect 3424 20791 3476 20800
rect 3424 20757 3433 20791
rect 3433 20757 3467 20791
rect 3467 20757 3476 20791
rect 3424 20748 3476 20757
rect 7288 20816 7340 20868
rect 8852 20884 8904 20936
rect 9496 20884 9548 20936
rect 9772 20884 9824 20936
rect 10508 20884 10560 20936
rect 11888 20884 11940 20936
rect 12900 20927 12952 20936
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 13268 20884 13320 20936
rect 14372 20995 14424 21004
rect 14372 20961 14381 20995
rect 14381 20961 14415 20995
rect 14415 20961 14424 20995
rect 14372 20952 14424 20961
rect 14464 20884 14516 20936
rect 15384 20927 15436 20936
rect 15384 20893 15393 20927
rect 15393 20893 15427 20927
rect 15427 20893 15436 20927
rect 15384 20884 15436 20893
rect 14556 20816 14608 20868
rect 14832 20816 14884 20868
rect 16304 21088 16356 21140
rect 16304 20859 16356 20868
rect 4252 20791 4304 20800
rect 4252 20757 4261 20791
rect 4261 20757 4295 20791
rect 4295 20757 4304 20791
rect 4252 20748 4304 20757
rect 4712 20791 4764 20800
rect 4712 20757 4721 20791
rect 4721 20757 4755 20791
rect 4755 20757 4764 20791
rect 4712 20748 4764 20757
rect 4896 20748 4948 20800
rect 5908 20748 5960 20800
rect 6276 20748 6328 20800
rect 6552 20748 6604 20800
rect 6920 20748 6972 20800
rect 7196 20748 7248 20800
rect 7656 20748 7708 20800
rect 8116 20748 8168 20800
rect 10416 20748 10468 20800
rect 10692 20748 10744 20800
rect 10876 20791 10928 20800
rect 10876 20757 10885 20791
rect 10885 20757 10919 20791
rect 10919 20757 10928 20791
rect 10876 20748 10928 20757
rect 12532 20748 12584 20800
rect 12808 20748 12860 20800
rect 13268 20791 13320 20800
rect 13268 20757 13277 20791
rect 13277 20757 13311 20791
rect 13311 20757 13320 20791
rect 13268 20748 13320 20757
rect 13360 20791 13412 20800
rect 13360 20757 13369 20791
rect 13369 20757 13403 20791
rect 13403 20757 13412 20791
rect 13360 20748 13412 20757
rect 14188 20748 14240 20800
rect 14740 20748 14792 20800
rect 14924 20791 14976 20800
rect 14924 20757 14933 20791
rect 14933 20757 14967 20791
rect 14967 20757 14976 20791
rect 14924 20748 14976 20757
rect 16304 20825 16313 20859
rect 16313 20825 16347 20859
rect 16347 20825 16356 20859
rect 16672 20952 16724 21004
rect 17408 20884 17460 20936
rect 18420 20952 18472 21004
rect 19156 20952 19208 21004
rect 18512 20884 18564 20936
rect 19708 21088 19760 21140
rect 20996 21088 21048 21140
rect 21456 21088 21508 21140
rect 22652 21131 22704 21140
rect 22652 21097 22661 21131
rect 22661 21097 22695 21131
rect 22695 21097 22704 21131
rect 22652 21088 22704 21097
rect 20904 20952 20956 21004
rect 21824 21020 21876 21072
rect 16672 20859 16724 20868
rect 16304 20816 16356 20825
rect 16672 20825 16681 20859
rect 16681 20825 16715 20859
rect 16715 20825 16724 20859
rect 16672 20816 16724 20825
rect 16948 20816 17000 20868
rect 15936 20748 15988 20800
rect 17132 20791 17184 20800
rect 17132 20757 17141 20791
rect 17141 20757 17175 20791
rect 17175 20757 17184 20791
rect 17132 20748 17184 20757
rect 20260 20816 20312 20868
rect 20536 20884 20588 20936
rect 20996 20884 21048 20936
rect 22284 20884 22336 20936
rect 23664 20884 23716 20936
rect 22192 20816 22244 20868
rect 18328 20748 18380 20800
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 19892 20748 19944 20800
rect 21180 20748 21232 20800
rect 22008 20791 22060 20800
rect 22008 20757 22017 20791
rect 22017 20757 22051 20791
rect 22051 20757 22060 20791
rect 23020 20791 23072 20800
rect 22008 20748 22060 20757
rect 23020 20757 23029 20791
rect 23029 20757 23063 20791
rect 23063 20757 23072 20791
rect 23020 20748 23072 20757
rect 6548 20646 6600 20698
rect 6612 20646 6664 20698
rect 6676 20646 6728 20698
rect 6740 20646 6792 20698
rect 6804 20646 6856 20698
rect 12146 20646 12198 20698
rect 12210 20646 12262 20698
rect 12274 20646 12326 20698
rect 12338 20646 12390 20698
rect 12402 20646 12454 20698
rect 17744 20646 17796 20698
rect 17808 20646 17860 20698
rect 17872 20646 17924 20698
rect 17936 20646 17988 20698
rect 18000 20646 18052 20698
rect 2320 20544 2372 20596
rect 2872 20587 2924 20596
rect 2872 20553 2881 20587
rect 2881 20553 2915 20587
rect 2915 20553 2924 20587
rect 2872 20544 2924 20553
rect 3516 20544 3568 20596
rect 4344 20544 4396 20596
rect 4620 20476 4672 20528
rect 5632 20544 5684 20596
rect 6736 20544 6788 20596
rect 5724 20476 5776 20528
rect 5816 20476 5868 20528
rect 8668 20544 8720 20596
rect 9496 20587 9548 20596
rect 9496 20553 9505 20587
rect 9505 20553 9539 20587
rect 9539 20553 9548 20587
rect 9496 20544 9548 20553
rect 10600 20544 10652 20596
rect 13360 20544 13412 20596
rect 3332 20408 3384 20460
rect 4160 20408 4212 20460
rect 3792 20340 3844 20392
rect 4436 20383 4488 20392
rect 4436 20349 4445 20383
rect 4445 20349 4479 20383
rect 4479 20349 4488 20383
rect 4620 20383 4672 20392
rect 4436 20340 4488 20349
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 3424 20204 3476 20256
rect 3608 20204 3660 20256
rect 4804 20272 4856 20324
rect 6000 20408 6052 20460
rect 8576 20451 8628 20460
rect 8576 20417 8585 20451
rect 8585 20417 8619 20451
rect 8619 20417 8628 20451
rect 8576 20408 8628 20417
rect 9772 20476 9824 20528
rect 11152 20476 11204 20528
rect 10324 20408 10376 20460
rect 10784 20408 10836 20460
rect 18144 20544 18196 20596
rect 18512 20544 18564 20596
rect 18880 20544 18932 20596
rect 19156 20544 19208 20596
rect 21548 20544 21600 20596
rect 22376 20544 22428 20596
rect 6736 20340 6788 20392
rect 8300 20383 8352 20392
rect 8300 20349 8309 20383
rect 8309 20349 8343 20383
rect 8343 20349 8352 20383
rect 8300 20340 8352 20349
rect 8668 20340 8720 20392
rect 4436 20204 4488 20256
rect 5816 20204 5868 20256
rect 6092 20204 6144 20256
rect 8944 20272 8996 20324
rect 9220 20272 9272 20324
rect 9680 20340 9732 20392
rect 11060 20340 11112 20392
rect 11152 20340 11204 20392
rect 12256 20383 12308 20392
rect 12256 20349 12265 20383
rect 12265 20349 12299 20383
rect 12299 20349 12308 20383
rect 14096 20408 14148 20460
rect 12256 20340 12308 20349
rect 14740 20383 14792 20392
rect 13452 20272 13504 20324
rect 14740 20349 14749 20383
rect 14749 20349 14783 20383
rect 14783 20349 14792 20383
rect 14740 20340 14792 20349
rect 16028 20408 16080 20460
rect 15292 20383 15344 20392
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 15476 20383 15528 20392
rect 15476 20349 15485 20383
rect 15485 20349 15519 20383
rect 15519 20349 15528 20383
rect 15476 20340 15528 20349
rect 16396 20451 16448 20460
rect 16396 20417 16405 20451
rect 16405 20417 16439 20451
rect 16439 20417 16448 20451
rect 16396 20408 16448 20417
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 16672 20340 16724 20392
rect 16948 20340 17000 20392
rect 17500 20476 17552 20528
rect 17868 20519 17920 20528
rect 17868 20485 17877 20519
rect 17877 20485 17911 20519
rect 17911 20485 17920 20519
rect 17868 20476 17920 20485
rect 19248 20476 19300 20528
rect 19064 20408 19116 20460
rect 14832 20272 14884 20324
rect 15660 20272 15712 20324
rect 13268 20204 13320 20256
rect 13544 20204 13596 20256
rect 14924 20204 14976 20256
rect 15568 20204 15620 20256
rect 17408 20340 17460 20392
rect 17960 20383 18012 20392
rect 17960 20349 17969 20383
rect 17969 20349 18003 20383
rect 18003 20349 18012 20383
rect 17960 20340 18012 20349
rect 18144 20383 18196 20392
rect 18144 20349 18153 20383
rect 18153 20349 18187 20383
rect 18187 20349 18196 20383
rect 18144 20340 18196 20349
rect 19892 20383 19944 20392
rect 17408 20204 17460 20256
rect 19892 20349 19901 20383
rect 19901 20349 19935 20383
rect 19935 20349 19944 20383
rect 19892 20340 19944 20349
rect 21364 20408 21416 20460
rect 22192 20408 22244 20460
rect 20628 20272 20680 20324
rect 20904 20340 20956 20392
rect 22928 20408 22980 20460
rect 23572 20340 23624 20392
rect 19340 20204 19392 20256
rect 23112 20272 23164 20324
rect 21088 20204 21140 20256
rect 21364 20247 21416 20256
rect 21364 20213 21373 20247
rect 21373 20213 21407 20247
rect 21407 20213 21416 20247
rect 21364 20204 21416 20213
rect 23296 20204 23348 20256
rect 3749 20102 3801 20154
rect 3813 20102 3865 20154
rect 3877 20102 3929 20154
rect 3941 20102 3993 20154
rect 4005 20102 4057 20154
rect 9347 20102 9399 20154
rect 9411 20102 9463 20154
rect 9475 20102 9527 20154
rect 9539 20102 9591 20154
rect 9603 20102 9655 20154
rect 14945 20102 14997 20154
rect 15009 20102 15061 20154
rect 15073 20102 15125 20154
rect 15137 20102 15189 20154
rect 15201 20102 15253 20154
rect 20543 20102 20595 20154
rect 20607 20102 20659 20154
rect 20671 20102 20723 20154
rect 20735 20102 20787 20154
rect 20799 20102 20851 20154
rect 4160 20043 4212 20052
rect 4160 20009 4169 20043
rect 4169 20009 4203 20043
rect 4203 20009 4212 20043
rect 4160 20000 4212 20009
rect 4344 20043 4396 20052
rect 4344 20009 4353 20043
rect 4353 20009 4387 20043
rect 4387 20009 4396 20043
rect 4344 20000 4396 20009
rect 5080 20000 5132 20052
rect 6000 20000 6052 20052
rect 6184 20000 6236 20052
rect 8392 20000 8444 20052
rect 10232 20000 10284 20052
rect 12808 20000 12860 20052
rect 13084 20000 13136 20052
rect 13360 20000 13412 20052
rect 14740 20000 14792 20052
rect 15200 20000 15252 20052
rect 5356 19932 5408 19984
rect 12072 19932 12124 19984
rect 14188 19932 14240 19984
rect 3608 19839 3660 19848
rect 3608 19805 3617 19839
rect 3617 19805 3651 19839
rect 3651 19805 3660 19839
rect 3608 19796 3660 19805
rect 4344 19796 4396 19848
rect 6092 19864 6144 19916
rect 12164 19864 12216 19916
rect 12808 19864 12860 19916
rect 13544 19864 13596 19916
rect 14096 19907 14148 19916
rect 14096 19873 14105 19907
rect 14105 19873 14139 19907
rect 14139 19873 14148 19907
rect 14096 19864 14148 19873
rect 17684 20000 17736 20052
rect 19064 20000 19116 20052
rect 20812 20000 20864 20052
rect 21272 20000 21324 20052
rect 23480 20000 23532 20052
rect 17500 19932 17552 19984
rect 16304 19864 16356 19916
rect 16764 19864 16816 19916
rect 17316 19907 17368 19916
rect 17316 19873 17325 19907
rect 17325 19873 17359 19907
rect 17359 19873 17368 19907
rect 17316 19864 17368 19873
rect 21088 19932 21140 19984
rect 22744 19932 22796 19984
rect 22100 19907 22152 19916
rect 22100 19873 22109 19907
rect 22109 19873 22143 19907
rect 22143 19873 22152 19907
rect 22100 19864 22152 19873
rect 5816 19796 5868 19848
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 10876 19796 10928 19848
rect 12716 19796 12768 19848
rect 13176 19796 13228 19848
rect 13360 19796 13412 19848
rect 3056 19660 3108 19712
rect 3516 19660 3568 19712
rect 5356 19771 5408 19780
rect 5356 19737 5365 19771
rect 5365 19737 5399 19771
rect 5399 19737 5408 19771
rect 5356 19728 5408 19737
rect 6092 19728 6144 19780
rect 7288 19728 7340 19780
rect 7564 19728 7616 19780
rect 8760 19728 8812 19780
rect 9220 19771 9272 19780
rect 9220 19737 9232 19771
rect 9232 19737 9272 19771
rect 9220 19728 9272 19737
rect 5264 19703 5316 19712
rect 5264 19669 5273 19703
rect 5273 19669 5307 19703
rect 5307 19669 5316 19703
rect 5264 19660 5316 19669
rect 5724 19703 5776 19712
rect 5724 19669 5733 19703
rect 5733 19669 5767 19703
rect 5767 19669 5776 19703
rect 5724 19660 5776 19669
rect 8852 19660 8904 19712
rect 11152 19728 11204 19780
rect 11980 19728 12032 19780
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10692 19703 10744 19712
rect 10416 19660 10468 19669
rect 10692 19669 10701 19703
rect 10701 19669 10735 19703
rect 10735 19669 10744 19703
rect 10692 19660 10744 19669
rect 13084 19703 13136 19712
rect 13084 19669 13093 19703
rect 13093 19669 13127 19703
rect 13127 19669 13136 19703
rect 13084 19660 13136 19669
rect 13176 19660 13228 19712
rect 15568 19796 15620 19848
rect 15660 19796 15712 19848
rect 15936 19796 15988 19848
rect 15292 19728 15344 19780
rect 16488 19728 16540 19780
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 19340 19796 19392 19848
rect 20444 19796 20496 19848
rect 20720 19796 20772 19848
rect 21456 19796 21508 19848
rect 22836 19839 22888 19848
rect 22836 19805 22845 19839
rect 22845 19805 22879 19839
rect 22879 19805 22888 19839
rect 22836 19796 22888 19805
rect 17960 19771 18012 19780
rect 15936 19660 15988 19712
rect 16028 19660 16080 19712
rect 16304 19660 16356 19712
rect 16580 19703 16632 19712
rect 16580 19669 16589 19703
rect 16589 19669 16623 19703
rect 16623 19669 16632 19703
rect 16580 19660 16632 19669
rect 16856 19660 16908 19712
rect 17224 19660 17276 19712
rect 17960 19737 17994 19771
rect 17994 19737 18012 19771
rect 17960 19728 18012 19737
rect 19616 19728 19668 19780
rect 17408 19660 17460 19712
rect 18604 19660 18656 19712
rect 20260 19728 20312 19780
rect 20352 19660 20404 19712
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 22284 19703 22336 19712
rect 22284 19669 22293 19703
rect 22293 19669 22327 19703
rect 22327 19669 22336 19703
rect 22284 19660 22336 19669
rect 22376 19703 22428 19712
rect 22376 19669 22385 19703
rect 22385 19669 22419 19703
rect 22419 19669 22428 19703
rect 22376 19660 22428 19669
rect 22560 19660 22612 19712
rect 23020 19703 23072 19712
rect 23020 19669 23029 19703
rect 23029 19669 23063 19703
rect 23063 19669 23072 19703
rect 23020 19660 23072 19669
rect 6548 19558 6600 19610
rect 6612 19558 6664 19610
rect 6676 19558 6728 19610
rect 6740 19558 6792 19610
rect 6804 19558 6856 19610
rect 12146 19558 12198 19610
rect 12210 19558 12262 19610
rect 12274 19558 12326 19610
rect 12338 19558 12390 19610
rect 12402 19558 12454 19610
rect 17744 19558 17796 19610
rect 17808 19558 17860 19610
rect 17872 19558 17924 19610
rect 17936 19558 17988 19610
rect 18000 19558 18052 19610
rect 3056 19499 3108 19508
rect 3056 19465 3065 19499
rect 3065 19465 3099 19499
rect 3099 19465 3108 19499
rect 3056 19456 3108 19465
rect 3240 19456 3292 19508
rect 4344 19499 4396 19508
rect 4344 19465 4353 19499
rect 4353 19465 4387 19499
rect 4387 19465 4396 19499
rect 4344 19456 4396 19465
rect 4620 19499 4672 19508
rect 4620 19465 4629 19499
rect 4629 19465 4663 19499
rect 4663 19465 4672 19499
rect 4620 19456 4672 19465
rect 5356 19456 5408 19508
rect 9680 19456 9732 19508
rect 9864 19456 9916 19508
rect 10968 19499 11020 19508
rect 10968 19465 10977 19499
rect 10977 19465 11011 19499
rect 11011 19465 11020 19499
rect 10968 19456 11020 19465
rect 11152 19499 11204 19508
rect 11152 19465 11161 19499
rect 11161 19465 11195 19499
rect 11195 19465 11204 19499
rect 11152 19456 11204 19465
rect 12072 19456 12124 19508
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 13636 19456 13688 19508
rect 15384 19456 15436 19508
rect 5816 19388 5868 19440
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 3608 19320 3660 19372
rect 4068 19320 4120 19372
rect 4436 19363 4488 19372
rect 4436 19329 4445 19363
rect 4445 19329 4479 19363
rect 4479 19329 4488 19363
rect 4436 19320 4488 19329
rect 4528 19320 4580 19372
rect 5172 19320 5224 19372
rect 6092 19320 6144 19372
rect 3424 19252 3476 19304
rect 4344 19252 4396 19304
rect 4804 19252 4856 19304
rect 10416 19388 10468 19440
rect 10876 19388 10928 19440
rect 8392 19363 8444 19372
rect 8392 19329 8426 19363
rect 8426 19329 8444 19363
rect 8392 19320 8444 19329
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 11336 19363 11388 19372
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 12808 19320 12860 19372
rect 13176 19320 13228 19372
rect 13636 19320 13688 19372
rect 13912 19363 13964 19372
rect 13912 19329 13921 19363
rect 13921 19329 13955 19363
rect 13955 19329 13964 19363
rect 13912 19320 13964 19329
rect 14372 19320 14424 19372
rect 15568 19388 15620 19440
rect 16396 19456 16448 19508
rect 16672 19499 16724 19508
rect 16672 19465 16681 19499
rect 16681 19465 16715 19499
rect 16715 19465 16724 19499
rect 16672 19456 16724 19465
rect 18328 19456 18380 19508
rect 19616 19499 19668 19508
rect 19616 19465 19625 19499
rect 19625 19465 19659 19499
rect 19659 19465 19668 19499
rect 19616 19456 19668 19465
rect 21088 19499 21140 19508
rect 21088 19465 21097 19499
rect 21097 19465 21131 19499
rect 21131 19465 21140 19499
rect 21088 19456 21140 19465
rect 21364 19456 21416 19508
rect 21456 19456 21508 19508
rect 16028 19388 16080 19440
rect 16764 19388 16816 19440
rect 17592 19388 17644 19440
rect 14740 19363 14792 19372
rect 14740 19329 14774 19363
rect 14774 19329 14792 19363
rect 15936 19363 15988 19372
rect 3240 19184 3292 19236
rect 3516 19116 3568 19168
rect 7748 19159 7800 19168
rect 7748 19125 7757 19159
rect 7757 19125 7791 19159
rect 7791 19125 7800 19159
rect 7748 19116 7800 19125
rect 8484 19116 8536 19168
rect 13728 19252 13780 19304
rect 14188 19252 14240 19304
rect 14740 19320 14792 19329
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 16120 19320 16172 19372
rect 16396 19363 16448 19372
rect 16396 19329 16405 19363
rect 16405 19329 16439 19363
rect 16439 19329 16448 19363
rect 16396 19320 16448 19329
rect 16488 19320 16540 19372
rect 19432 19320 19484 19372
rect 20444 19388 20496 19440
rect 20904 19320 20956 19372
rect 21272 19363 21324 19372
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21272 19320 21324 19329
rect 24124 19388 24176 19440
rect 22836 19363 22888 19372
rect 16764 19252 16816 19304
rect 15200 19116 15252 19168
rect 15384 19116 15436 19168
rect 15660 19116 15712 19168
rect 18512 19116 18564 19168
rect 21272 19116 21324 19168
rect 22836 19329 22845 19363
rect 22845 19329 22879 19363
rect 22879 19329 22888 19363
rect 22836 19320 22888 19329
rect 21732 19252 21784 19304
rect 22468 19295 22520 19304
rect 22468 19261 22477 19295
rect 22477 19261 22511 19295
rect 22511 19261 22520 19295
rect 22468 19252 22520 19261
rect 23112 19252 23164 19304
rect 21833 19227 21885 19236
rect 21833 19193 21867 19227
rect 21867 19193 21885 19227
rect 21833 19184 21885 19193
rect 21640 19116 21692 19168
rect 21732 19116 21784 19168
rect 23112 19116 23164 19168
rect 3749 19014 3801 19066
rect 3813 19014 3865 19066
rect 3877 19014 3929 19066
rect 3941 19014 3993 19066
rect 4005 19014 4057 19066
rect 9347 19014 9399 19066
rect 9411 19014 9463 19066
rect 9475 19014 9527 19066
rect 9539 19014 9591 19066
rect 9603 19014 9655 19066
rect 14945 19014 14997 19066
rect 15009 19014 15061 19066
rect 15073 19014 15125 19066
rect 15137 19014 15189 19066
rect 15201 19014 15253 19066
rect 20543 19014 20595 19066
rect 20607 19014 20659 19066
rect 20671 19014 20723 19066
rect 20735 19014 20787 19066
rect 20799 19014 20851 19066
rect 3516 18912 3568 18964
rect 4160 18912 4212 18964
rect 4804 18912 4856 18964
rect 3608 18887 3660 18896
rect 3608 18853 3617 18887
rect 3617 18853 3651 18887
rect 3651 18853 3660 18887
rect 3608 18844 3660 18853
rect 6368 18912 6420 18964
rect 8760 18955 8812 18964
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 11796 18912 11848 18964
rect 12808 18912 12860 18964
rect 14096 18912 14148 18964
rect 15292 18912 15344 18964
rect 17040 18955 17092 18964
rect 3424 18776 3476 18828
rect 5816 18819 5868 18828
rect 5816 18785 5825 18819
rect 5825 18785 5859 18819
rect 5859 18785 5868 18819
rect 5816 18776 5868 18785
rect 8576 18776 8628 18828
rect 10968 18776 11020 18828
rect 5172 18708 5224 18760
rect 5724 18708 5776 18760
rect 7380 18751 7432 18760
rect 7380 18717 7389 18751
rect 7389 18717 7423 18751
rect 7423 18717 7432 18751
rect 7380 18708 7432 18717
rect 9680 18708 9732 18760
rect 9864 18751 9916 18760
rect 9864 18717 9898 18751
rect 9898 18717 9916 18751
rect 9864 18708 9916 18717
rect 3240 18683 3292 18692
rect 3240 18649 3249 18683
rect 3249 18649 3283 18683
rect 3283 18649 3292 18683
rect 3240 18640 3292 18649
rect 7012 18683 7064 18692
rect 2964 18572 3016 18624
rect 3516 18572 3568 18624
rect 5356 18572 5408 18624
rect 7012 18649 7030 18683
rect 7030 18649 7064 18683
rect 7012 18640 7064 18649
rect 8300 18640 8352 18692
rect 10876 18640 10928 18692
rect 14188 18708 14240 18760
rect 11428 18640 11480 18692
rect 15384 18708 15436 18760
rect 15568 18751 15620 18760
rect 15568 18717 15577 18751
rect 15577 18717 15611 18751
rect 15611 18717 15620 18751
rect 15568 18708 15620 18717
rect 16396 18708 16448 18760
rect 14924 18640 14976 18692
rect 6000 18572 6052 18624
rect 7104 18572 7156 18624
rect 7748 18572 7800 18624
rect 12992 18572 13044 18624
rect 13084 18572 13136 18624
rect 16028 18640 16080 18692
rect 16120 18572 16172 18624
rect 17040 18921 17049 18955
rect 17049 18921 17083 18955
rect 17083 18921 17092 18955
rect 17040 18912 17092 18921
rect 18052 18912 18104 18964
rect 18144 18912 18196 18964
rect 18696 18912 18748 18964
rect 19616 18912 19668 18964
rect 20996 18844 21048 18896
rect 16948 18708 17000 18760
rect 18328 18708 18380 18760
rect 18880 18708 18932 18760
rect 22744 18819 22796 18828
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 19340 18708 19392 18760
rect 20536 18708 20588 18760
rect 20720 18708 20772 18760
rect 23020 18751 23072 18760
rect 23020 18717 23029 18751
rect 23029 18717 23063 18751
rect 23063 18717 23072 18751
rect 23020 18708 23072 18717
rect 17500 18640 17552 18692
rect 18604 18640 18656 18692
rect 17592 18572 17644 18624
rect 19616 18572 19668 18624
rect 20352 18683 20404 18692
rect 20352 18649 20392 18683
rect 20392 18649 20404 18683
rect 20352 18640 20404 18649
rect 21916 18572 21968 18624
rect 22284 18572 22336 18624
rect 6548 18470 6600 18522
rect 6612 18470 6664 18522
rect 6676 18470 6728 18522
rect 6740 18470 6792 18522
rect 6804 18470 6856 18522
rect 12146 18470 12198 18522
rect 12210 18470 12262 18522
rect 12274 18470 12326 18522
rect 12338 18470 12390 18522
rect 12402 18470 12454 18522
rect 17744 18470 17796 18522
rect 17808 18470 17860 18522
rect 17872 18470 17924 18522
rect 17936 18470 17988 18522
rect 18000 18470 18052 18522
rect 2872 18368 2924 18420
rect 3332 18368 3384 18420
rect 3516 18300 3568 18352
rect 4804 18368 4856 18420
rect 7104 18300 7156 18352
rect 7380 18368 7432 18420
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 10232 18368 10284 18420
rect 10876 18368 10928 18420
rect 9036 18300 9088 18352
rect 3240 18232 3292 18284
rect 3424 18232 3476 18284
rect 2964 18207 3016 18216
rect 2964 18173 2973 18207
rect 2973 18173 3007 18207
rect 3007 18173 3016 18207
rect 2964 18164 3016 18173
rect 3884 18164 3936 18216
rect 3424 18096 3476 18148
rect 4160 18164 4212 18216
rect 4620 18164 4672 18216
rect 5264 18164 5316 18216
rect 6460 18232 6512 18284
rect 9772 18232 9824 18284
rect 10508 18232 10560 18284
rect 14004 18368 14056 18420
rect 14740 18368 14792 18420
rect 17316 18368 17368 18420
rect 17592 18368 17644 18420
rect 22284 18411 22336 18420
rect 22284 18377 22293 18411
rect 22293 18377 22327 18411
rect 22327 18377 22336 18411
rect 22284 18368 22336 18377
rect 22744 18411 22796 18420
rect 22744 18377 22753 18411
rect 22753 18377 22787 18411
rect 22787 18377 22796 18411
rect 22744 18368 22796 18377
rect 12072 18300 12124 18352
rect 12624 18300 12676 18352
rect 5356 18096 5408 18148
rect 6184 18164 6236 18216
rect 14280 18275 14332 18284
rect 15568 18300 15620 18352
rect 16212 18300 16264 18352
rect 14280 18241 14298 18275
rect 14298 18241 14332 18275
rect 14280 18232 14332 18241
rect 3056 18028 3108 18080
rect 4988 18028 5040 18080
rect 6092 18071 6144 18080
rect 6092 18037 6101 18071
rect 6101 18037 6135 18071
rect 6135 18037 6144 18071
rect 8300 18096 8352 18148
rect 11428 18096 11480 18148
rect 13084 18139 13136 18148
rect 13084 18105 13093 18139
rect 13093 18105 13127 18139
rect 13127 18105 13136 18139
rect 13084 18096 13136 18105
rect 13176 18139 13228 18148
rect 13176 18105 13185 18139
rect 13185 18105 13219 18139
rect 13219 18105 13228 18139
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 16396 18164 16448 18216
rect 17132 18300 17184 18352
rect 17040 18232 17092 18284
rect 18052 18300 18104 18352
rect 18604 18300 18656 18352
rect 19340 18300 19392 18352
rect 20168 18300 20220 18352
rect 20628 18300 20680 18352
rect 21732 18300 21784 18352
rect 19432 18232 19484 18284
rect 19892 18232 19944 18284
rect 18236 18207 18288 18216
rect 18236 18173 18245 18207
rect 18245 18173 18279 18207
rect 18279 18173 18288 18207
rect 18236 18164 18288 18173
rect 13176 18096 13228 18105
rect 6092 18028 6144 18037
rect 8852 18028 8904 18080
rect 11244 18028 11296 18080
rect 11704 18028 11756 18080
rect 14648 18028 14700 18080
rect 18328 18096 18380 18148
rect 16120 18028 16172 18080
rect 16396 18071 16448 18080
rect 16396 18037 16405 18071
rect 16405 18037 16439 18071
rect 16439 18037 16448 18071
rect 16396 18028 16448 18037
rect 17592 18028 17644 18080
rect 18144 18028 18196 18080
rect 18788 18028 18840 18080
rect 20996 18232 21048 18284
rect 20076 18164 20128 18216
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 20168 18139 20220 18148
rect 20168 18105 20177 18139
rect 20177 18105 20211 18139
rect 20211 18105 20220 18139
rect 20168 18096 20220 18105
rect 21272 18096 21324 18148
rect 20260 18028 20312 18080
rect 21548 18028 21600 18080
rect 21916 18028 21968 18080
rect 3749 17926 3801 17978
rect 3813 17926 3865 17978
rect 3877 17926 3929 17978
rect 3941 17926 3993 17978
rect 4005 17926 4057 17978
rect 9347 17926 9399 17978
rect 9411 17926 9463 17978
rect 9475 17926 9527 17978
rect 9539 17926 9591 17978
rect 9603 17926 9655 17978
rect 14945 17926 14997 17978
rect 15009 17926 15061 17978
rect 15073 17926 15125 17978
rect 15137 17926 15189 17978
rect 15201 17926 15253 17978
rect 20543 17926 20595 17978
rect 20607 17926 20659 17978
rect 20671 17926 20723 17978
rect 20735 17926 20787 17978
rect 20799 17926 20851 17978
rect 3148 17824 3200 17876
rect 5908 17867 5960 17876
rect 5908 17833 5917 17867
rect 5917 17833 5951 17867
rect 5951 17833 5960 17867
rect 5908 17824 5960 17833
rect 6276 17824 6328 17876
rect 11244 17824 11296 17876
rect 13176 17824 13228 17876
rect 14464 17824 14516 17876
rect 16580 17824 16632 17876
rect 18972 17824 19024 17876
rect 19524 17824 19576 17876
rect 19984 17824 20036 17876
rect 20444 17824 20496 17876
rect 19248 17799 19300 17808
rect 19248 17765 19257 17799
rect 19257 17765 19291 17799
rect 19291 17765 19300 17799
rect 19248 17756 19300 17765
rect 21364 17824 21416 17876
rect 21732 17867 21784 17876
rect 21732 17833 21741 17867
rect 21741 17833 21775 17867
rect 21775 17833 21784 17867
rect 21732 17824 21784 17833
rect 22468 17824 22520 17876
rect 23204 17824 23256 17876
rect 2872 17688 2924 17740
rect 3424 17688 3476 17740
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 3608 17620 3660 17672
rect 6092 17620 6144 17672
rect 9128 17620 9180 17672
rect 11060 17663 11112 17672
rect 11060 17629 11069 17663
rect 11069 17629 11103 17663
rect 11103 17629 11112 17663
rect 11060 17620 11112 17629
rect 12992 17620 13044 17672
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 14096 17663 14148 17672
rect 13728 17620 13780 17629
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 16396 17620 16448 17672
rect 17132 17663 17184 17672
rect 17132 17629 17141 17663
rect 17141 17629 17175 17663
rect 17175 17629 17184 17663
rect 17132 17620 17184 17629
rect 21364 17688 21416 17740
rect 22100 17688 22152 17740
rect 19340 17620 19392 17672
rect 4712 17595 4764 17604
rect 4068 17484 4120 17536
rect 4712 17561 4746 17595
rect 4746 17561 4764 17595
rect 4712 17552 4764 17561
rect 4804 17552 4856 17604
rect 5724 17552 5776 17604
rect 6000 17552 6052 17604
rect 7196 17552 7248 17604
rect 10232 17552 10284 17604
rect 12532 17595 12584 17604
rect 12532 17561 12566 17595
rect 12566 17561 12584 17595
rect 12532 17552 12584 17561
rect 5080 17484 5132 17536
rect 7380 17527 7432 17536
rect 7380 17493 7389 17527
rect 7389 17493 7423 17527
rect 7423 17493 7432 17527
rect 7380 17484 7432 17493
rect 7472 17484 7524 17536
rect 10324 17484 10376 17536
rect 14188 17484 14240 17536
rect 14556 17484 14608 17536
rect 14832 17484 14884 17536
rect 16672 17595 16724 17604
rect 16672 17561 16690 17595
rect 16690 17561 16724 17595
rect 16672 17552 16724 17561
rect 17408 17484 17460 17536
rect 18052 17552 18104 17604
rect 18144 17552 18196 17604
rect 18604 17552 18656 17604
rect 19616 17552 19668 17604
rect 20168 17552 20220 17604
rect 20352 17595 20404 17604
rect 20352 17561 20370 17595
rect 20370 17561 20404 17595
rect 20352 17552 20404 17561
rect 20720 17620 20772 17672
rect 21548 17663 21600 17672
rect 21548 17629 21557 17663
rect 21557 17629 21591 17663
rect 21591 17629 21600 17663
rect 21548 17620 21600 17629
rect 22284 17552 22336 17604
rect 21088 17527 21140 17536
rect 21088 17493 21097 17527
rect 21097 17493 21131 17527
rect 21131 17493 21140 17527
rect 21088 17484 21140 17493
rect 21272 17484 21324 17536
rect 22192 17527 22244 17536
rect 22192 17493 22201 17527
rect 22201 17493 22235 17527
rect 22235 17493 22244 17527
rect 22192 17484 22244 17493
rect 22468 17484 22520 17536
rect 23112 17527 23164 17536
rect 23112 17493 23121 17527
rect 23121 17493 23155 17527
rect 23155 17493 23164 17527
rect 23112 17484 23164 17493
rect 6548 17382 6600 17434
rect 6612 17382 6664 17434
rect 6676 17382 6728 17434
rect 6740 17382 6792 17434
rect 6804 17382 6856 17434
rect 12146 17382 12198 17434
rect 12210 17382 12262 17434
rect 12274 17382 12326 17434
rect 12338 17382 12390 17434
rect 12402 17382 12454 17434
rect 17744 17382 17796 17434
rect 17808 17382 17860 17434
rect 17872 17382 17924 17434
rect 17936 17382 17988 17434
rect 18000 17382 18052 17434
rect 4620 17280 4672 17332
rect 6276 17280 6328 17332
rect 8024 17280 8076 17332
rect 9036 17323 9088 17332
rect 9036 17289 9045 17323
rect 9045 17289 9079 17323
rect 9079 17289 9088 17323
rect 9036 17280 9088 17289
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 11060 17323 11112 17332
rect 11060 17289 11069 17323
rect 11069 17289 11103 17323
rect 11103 17289 11112 17323
rect 11060 17280 11112 17289
rect 11520 17280 11572 17332
rect 15292 17280 15344 17332
rect 16212 17323 16264 17332
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 17500 17280 17552 17332
rect 18328 17280 18380 17332
rect 18604 17323 18656 17332
rect 18604 17289 18613 17323
rect 18613 17289 18647 17323
rect 18647 17289 18656 17323
rect 18604 17280 18656 17289
rect 19432 17280 19484 17332
rect 19800 17280 19852 17332
rect 20168 17280 20220 17332
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 4896 17212 4948 17264
rect 5540 17212 5592 17264
rect 6184 17212 6236 17264
rect 4528 17144 4580 17196
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 6828 17119 6880 17128
rect 4804 17076 4856 17085
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 8944 17212 8996 17264
rect 7748 17144 7800 17196
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 4160 17008 4212 17060
rect 4712 16940 4764 16992
rect 5540 16940 5592 16992
rect 7288 17008 7340 17060
rect 6552 16940 6604 16992
rect 9036 17076 9088 17128
rect 12716 17187 12768 17196
rect 12716 17153 12734 17187
rect 12734 17153 12768 17187
rect 12716 17144 12768 17153
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 14096 17212 14148 17264
rect 12992 17144 13044 17153
rect 14004 17187 14056 17196
rect 14004 17153 14013 17187
rect 14013 17153 14047 17187
rect 14047 17153 14056 17187
rect 14004 17144 14056 17153
rect 14464 17144 14516 17196
rect 16396 17212 16448 17264
rect 14648 17144 14700 17196
rect 16028 17187 16080 17196
rect 16028 17153 16037 17187
rect 16037 17153 16071 17187
rect 16071 17153 16080 17187
rect 16028 17144 16080 17153
rect 17316 17212 17368 17264
rect 17776 17255 17828 17264
rect 17776 17221 17794 17255
rect 17794 17221 17828 17255
rect 17776 17212 17828 17221
rect 18788 17212 18840 17264
rect 20076 17212 20128 17264
rect 20720 17212 20772 17264
rect 23020 17323 23072 17332
rect 23020 17289 23029 17323
rect 23029 17289 23063 17323
rect 23063 17289 23072 17323
rect 23020 17280 23072 17289
rect 21364 17255 21416 17264
rect 21364 17221 21373 17255
rect 21373 17221 21407 17255
rect 21407 17221 21416 17255
rect 21364 17212 21416 17221
rect 22100 17212 22152 17264
rect 22468 17212 22520 17264
rect 10232 17008 10284 17060
rect 11888 16940 11940 16992
rect 13820 17008 13872 17060
rect 14004 17008 14056 17060
rect 14464 17051 14516 17060
rect 14464 17017 14473 17051
rect 14473 17017 14507 17051
rect 14507 17017 14516 17051
rect 14464 17008 14516 17017
rect 16948 17076 17000 17128
rect 15660 17008 15712 17060
rect 18144 17144 18196 17196
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 19800 17187 19852 17196
rect 19800 17153 19818 17187
rect 19818 17153 19852 17187
rect 19800 17144 19852 17153
rect 19984 17144 20036 17196
rect 20996 17144 21048 17196
rect 22560 17144 22612 17196
rect 23296 17144 23348 17196
rect 19064 17076 19116 17128
rect 20076 17119 20128 17128
rect 20076 17085 20085 17119
rect 20085 17085 20119 17119
rect 20119 17085 20128 17119
rect 20076 17076 20128 17085
rect 21364 17076 21416 17128
rect 22100 17119 22152 17128
rect 22100 17085 22109 17119
rect 22109 17085 22143 17119
rect 22143 17085 22152 17119
rect 22100 17076 22152 17085
rect 18328 17008 18380 17060
rect 18512 17008 18564 17060
rect 20904 17008 20956 17060
rect 21640 17008 21692 17060
rect 22928 17051 22980 17060
rect 22928 17017 22937 17051
rect 22937 17017 22971 17051
rect 22971 17017 22980 17051
rect 22928 17008 22980 17017
rect 15936 16983 15988 16992
rect 15936 16949 15945 16983
rect 15945 16949 15979 16983
rect 15979 16949 15988 16983
rect 15936 16940 15988 16949
rect 16028 16940 16080 16992
rect 16396 16940 16448 16992
rect 16672 16940 16724 16992
rect 21088 16940 21140 16992
rect 21364 16940 21416 16992
rect 22008 16940 22060 16992
rect 22744 16940 22796 16992
rect 3749 16838 3801 16890
rect 3813 16838 3865 16890
rect 3877 16838 3929 16890
rect 3941 16838 3993 16890
rect 4005 16838 4057 16890
rect 9347 16838 9399 16890
rect 9411 16838 9463 16890
rect 9475 16838 9527 16890
rect 9539 16838 9591 16890
rect 9603 16838 9655 16890
rect 14945 16838 14997 16890
rect 15009 16838 15061 16890
rect 15073 16838 15125 16890
rect 15137 16838 15189 16890
rect 15201 16838 15253 16890
rect 20543 16838 20595 16890
rect 20607 16838 20659 16890
rect 20671 16838 20723 16890
rect 20735 16838 20787 16890
rect 20799 16838 20851 16890
rect 4160 16779 4212 16788
rect 4160 16745 4169 16779
rect 4169 16745 4203 16779
rect 4203 16745 4212 16779
rect 4160 16736 4212 16745
rect 4804 16736 4856 16788
rect 6552 16736 6604 16788
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 9680 16736 9732 16788
rect 12716 16736 12768 16788
rect 5172 16711 5224 16720
rect 5172 16677 5181 16711
rect 5181 16677 5215 16711
rect 5215 16677 5224 16711
rect 5172 16668 5224 16677
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 11612 16668 11664 16720
rect 16212 16736 16264 16788
rect 17776 16736 17828 16788
rect 18604 16736 18656 16788
rect 14096 16711 14148 16720
rect 14096 16677 14105 16711
rect 14105 16677 14139 16711
rect 14139 16677 14148 16711
rect 14096 16668 14148 16677
rect 8944 16600 8996 16652
rect 6276 16575 6328 16584
rect 6276 16541 6294 16575
rect 6294 16541 6328 16575
rect 6276 16532 6328 16541
rect 6460 16464 6512 16516
rect 6828 16464 6880 16516
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 8116 16439 8168 16448
rect 4620 16396 4672 16405
rect 8116 16405 8125 16439
rect 8125 16405 8159 16439
rect 8159 16405 8168 16439
rect 10232 16464 10284 16516
rect 10692 16464 10744 16516
rect 13636 16507 13688 16516
rect 13636 16473 13654 16507
rect 13654 16473 13688 16507
rect 13636 16464 13688 16473
rect 14096 16464 14148 16516
rect 14280 16464 14332 16516
rect 16672 16575 16724 16584
rect 16672 16541 16690 16575
rect 16690 16541 16724 16575
rect 16672 16532 16724 16541
rect 16580 16464 16632 16516
rect 17592 16532 17644 16584
rect 20444 16736 20496 16788
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 19524 16575 19576 16584
rect 19524 16541 19558 16575
rect 19558 16541 19576 16575
rect 19524 16532 19576 16541
rect 19800 16532 19852 16584
rect 20904 16736 20956 16788
rect 21364 16600 21416 16652
rect 21272 16532 21324 16584
rect 22192 16736 22244 16788
rect 23020 16779 23072 16788
rect 23020 16745 23029 16779
rect 23029 16745 23063 16779
rect 23063 16745 23072 16779
rect 23020 16736 23072 16745
rect 22560 16668 22612 16720
rect 22008 16600 22060 16652
rect 22560 16532 22612 16584
rect 8116 16396 8168 16405
rect 9220 16439 9272 16448
rect 9220 16405 9229 16439
rect 9229 16405 9263 16439
rect 9263 16405 9272 16439
rect 9220 16396 9272 16405
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 15384 16396 15436 16448
rect 15568 16439 15620 16448
rect 15568 16405 15577 16439
rect 15577 16405 15611 16439
rect 15611 16405 15620 16439
rect 20628 16464 20680 16516
rect 21916 16464 21968 16516
rect 15568 16396 15620 16405
rect 20996 16396 21048 16448
rect 21732 16396 21784 16448
rect 22376 16396 22428 16448
rect 22652 16396 22704 16448
rect 6548 16294 6600 16346
rect 6612 16294 6664 16346
rect 6676 16294 6728 16346
rect 6740 16294 6792 16346
rect 6804 16294 6856 16346
rect 12146 16294 12198 16346
rect 12210 16294 12262 16346
rect 12274 16294 12326 16346
rect 12338 16294 12390 16346
rect 12402 16294 12454 16346
rect 17744 16294 17796 16346
rect 17808 16294 17860 16346
rect 17872 16294 17924 16346
rect 17936 16294 17988 16346
rect 18000 16294 18052 16346
rect 3608 16192 3660 16244
rect 12440 16192 12492 16244
rect 16764 16192 16816 16244
rect 4528 16124 4580 16176
rect 4804 16124 4856 16176
rect 5540 16056 5592 16108
rect 5908 16099 5960 16108
rect 6920 16124 6972 16176
rect 5908 16065 5926 16099
rect 5926 16065 5960 16099
rect 5908 16056 5960 16065
rect 3516 15920 3568 15972
rect 4344 15988 4396 16040
rect 8116 16099 8168 16108
rect 8116 16065 8125 16099
rect 8125 16065 8159 16099
rect 8159 16065 8168 16099
rect 8116 16056 8168 16065
rect 8208 16056 8260 16108
rect 8852 15988 8904 16040
rect 4620 15920 4672 15972
rect 4896 15920 4948 15972
rect 6368 15920 6420 15972
rect 7656 15852 7708 15904
rect 9036 16031 9088 16040
rect 9036 15997 9045 16031
rect 9045 15997 9079 16031
rect 9079 15997 9088 16031
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 11428 16056 11480 16108
rect 12808 16056 12860 16108
rect 15568 16124 15620 16176
rect 16028 16124 16080 16176
rect 16488 16124 16540 16176
rect 17040 16124 17092 16176
rect 18236 16192 18288 16244
rect 18512 16192 18564 16244
rect 19984 16192 20036 16244
rect 20352 16192 20404 16244
rect 15752 16056 15804 16108
rect 16580 16056 16632 16108
rect 20168 16124 20220 16176
rect 21088 16192 21140 16244
rect 22284 16192 22336 16244
rect 22560 16235 22612 16244
rect 22560 16201 22569 16235
rect 22569 16201 22603 16235
rect 22603 16201 22612 16235
rect 22560 16192 22612 16201
rect 9036 15988 9088 15997
rect 16488 15963 16540 15972
rect 16488 15929 16497 15963
rect 16497 15929 16531 15963
rect 16531 15929 16540 15963
rect 16488 15920 16540 15929
rect 19064 15988 19116 16040
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 18696 15920 18748 15972
rect 20444 15988 20496 16040
rect 20904 16056 20956 16108
rect 21272 16056 21324 16108
rect 21916 16056 21968 16108
rect 22376 16124 22428 16176
rect 23204 16124 23256 16176
rect 21732 15988 21784 16040
rect 22468 16056 22520 16108
rect 22928 16099 22980 16108
rect 22928 16065 22937 16099
rect 22937 16065 22971 16099
rect 22971 16065 22980 16099
rect 22928 16056 22980 16065
rect 22376 15988 22428 16040
rect 21916 15920 21968 15972
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 12256 15852 12308 15861
rect 12624 15852 12676 15904
rect 14280 15852 14332 15904
rect 14556 15895 14608 15904
rect 14556 15861 14565 15895
rect 14565 15861 14599 15895
rect 14599 15861 14608 15895
rect 14556 15852 14608 15861
rect 15108 15852 15160 15904
rect 16672 15852 16724 15904
rect 17316 15852 17368 15904
rect 19156 15852 19208 15904
rect 19340 15852 19392 15904
rect 22928 15920 22980 15972
rect 22468 15852 22520 15904
rect 23112 15895 23164 15904
rect 23112 15861 23121 15895
rect 23121 15861 23155 15895
rect 23155 15861 23164 15895
rect 23112 15852 23164 15861
rect 3749 15750 3801 15802
rect 3813 15750 3865 15802
rect 3877 15750 3929 15802
rect 3941 15750 3993 15802
rect 4005 15750 4057 15802
rect 9347 15750 9399 15802
rect 9411 15750 9463 15802
rect 9475 15750 9527 15802
rect 9539 15750 9591 15802
rect 9603 15750 9655 15802
rect 14945 15750 14997 15802
rect 15009 15750 15061 15802
rect 15073 15750 15125 15802
rect 15137 15750 15189 15802
rect 15201 15750 15253 15802
rect 20543 15750 20595 15802
rect 20607 15750 20659 15802
rect 20671 15750 20723 15802
rect 20735 15750 20787 15802
rect 20799 15750 20851 15802
rect 4436 15648 4488 15700
rect 4804 15648 4856 15700
rect 4344 15512 4396 15564
rect 6460 15648 6512 15700
rect 9128 15648 9180 15700
rect 11796 15648 11848 15700
rect 12440 15648 12492 15700
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 14648 15648 14700 15700
rect 15476 15648 15528 15700
rect 16212 15691 16264 15700
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 17408 15648 17460 15700
rect 6276 15580 6328 15632
rect 15660 15580 15712 15632
rect 15844 15580 15896 15632
rect 18328 15648 18380 15700
rect 19524 15648 19576 15700
rect 20352 15648 20404 15700
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 8208 15444 8260 15496
rect 10692 15512 10744 15564
rect 11336 15444 11388 15496
rect 14832 15512 14884 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 15936 15512 15988 15564
rect 18236 15512 18288 15564
rect 20536 15580 20588 15632
rect 19248 15555 19300 15564
rect 19248 15521 19257 15555
rect 19257 15521 19291 15555
rect 19291 15521 19300 15555
rect 19248 15512 19300 15521
rect 21272 15512 21324 15564
rect 5356 15376 5408 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 7748 15376 7800 15428
rect 9312 15376 9364 15428
rect 13452 15376 13504 15428
rect 15660 15376 15712 15428
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 16948 15376 17000 15428
rect 9220 15308 9272 15360
rect 10784 15308 10836 15360
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 16672 15351 16724 15360
rect 16672 15317 16681 15351
rect 16681 15317 16715 15351
rect 16715 15317 16724 15351
rect 16672 15308 16724 15317
rect 17040 15308 17092 15360
rect 18144 15487 18196 15496
rect 18144 15453 18153 15487
rect 18153 15453 18187 15487
rect 18187 15453 18196 15487
rect 21824 15648 21876 15700
rect 22376 15691 22428 15700
rect 22376 15657 22385 15691
rect 22385 15657 22419 15691
rect 22419 15657 22428 15691
rect 22376 15648 22428 15657
rect 22008 15580 22060 15632
rect 22100 15580 22152 15632
rect 21824 15512 21876 15564
rect 18144 15444 18196 15453
rect 18604 15419 18656 15428
rect 18604 15385 18613 15419
rect 18613 15385 18647 15419
rect 18647 15385 18656 15419
rect 18604 15376 18656 15385
rect 19064 15376 19116 15428
rect 21640 15444 21692 15496
rect 22744 15444 22796 15496
rect 20444 15376 20496 15428
rect 20536 15376 20588 15428
rect 20904 15308 20956 15360
rect 21088 15351 21140 15360
rect 21088 15317 21097 15351
rect 21097 15317 21131 15351
rect 21131 15317 21140 15351
rect 21088 15308 21140 15317
rect 21180 15351 21232 15360
rect 21180 15317 21189 15351
rect 21189 15317 21223 15351
rect 21223 15317 21232 15351
rect 21180 15308 21232 15317
rect 21824 15308 21876 15360
rect 21916 15351 21968 15360
rect 21916 15317 21925 15351
rect 21925 15317 21959 15351
rect 21959 15317 21968 15351
rect 22744 15351 22796 15360
rect 21916 15308 21968 15317
rect 22744 15317 22753 15351
rect 22753 15317 22787 15351
rect 22787 15317 22796 15351
rect 22744 15308 22796 15317
rect 6548 15206 6600 15258
rect 6612 15206 6664 15258
rect 6676 15206 6728 15258
rect 6740 15206 6792 15258
rect 6804 15206 6856 15258
rect 12146 15206 12198 15258
rect 12210 15206 12262 15258
rect 12274 15206 12326 15258
rect 12338 15206 12390 15258
rect 12402 15206 12454 15258
rect 17744 15206 17796 15258
rect 17808 15206 17860 15258
rect 17872 15206 17924 15258
rect 17936 15206 17988 15258
rect 18000 15206 18052 15258
rect 5080 15104 5132 15156
rect 5724 15036 5776 15088
rect 7380 15036 7432 15088
rect 4896 15011 4948 15020
rect 4896 14977 4905 15011
rect 4905 14977 4939 15011
rect 4939 14977 4948 15011
rect 4896 14968 4948 14977
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 6276 14968 6328 15020
rect 6920 14968 6972 15020
rect 8208 15104 8260 15156
rect 11796 15104 11848 15156
rect 13452 15147 13504 15156
rect 13452 15113 13461 15147
rect 13461 15113 13495 15147
rect 13495 15113 13504 15147
rect 13452 15104 13504 15113
rect 10784 14968 10836 15020
rect 11336 15011 11388 15020
rect 11336 14977 11345 15011
rect 11345 14977 11379 15011
rect 11379 14977 11388 15011
rect 11336 14968 11388 14977
rect 5540 14900 5592 14952
rect 5908 14900 5960 14952
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 4712 14764 4764 14816
rect 6368 14764 6420 14816
rect 6644 14764 6696 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 11060 14764 11112 14816
rect 13636 15036 13688 15088
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 15568 15104 15620 15156
rect 17224 15104 17276 15156
rect 19340 15104 19392 15156
rect 21640 15147 21692 15156
rect 15476 15011 15528 15020
rect 15476 14977 15494 15011
rect 15494 14977 15528 15011
rect 15476 14968 15528 14977
rect 15660 14968 15712 15020
rect 16212 14968 16264 15020
rect 16764 14968 16816 15020
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 11796 14900 11848 14952
rect 12440 14900 12492 14952
rect 15844 14832 15896 14884
rect 16488 14832 16540 14884
rect 19156 14900 19208 14952
rect 21640 15113 21649 15147
rect 21649 15113 21683 15147
rect 21683 15113 21692 15147
rect 21640 15104 21692 15113
rect 22468 15147 22520 15156
rect 22468 15113 22477 15147
rect 22477 15113 22511 15147
rect 22511 15113 22520 15147
rect 22468 15104 22520 15113
rect 22744 15104 22796 15156
rect 21916 15036 21968 15088
rect 19616 14968 19668 15020
rect 21732 14968 21784 15020
rect 23204 14968 23256 15020
rect 19524 14875 19576 14884
rect 19524 14841 19533 14875
rect 19533 14841 19567 14875
rect 19567 14841 19576 14875
rect 19524 14832 19576 14841
rect 12624 14764 12676 14816
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 13360 14764 13412 14816
rect 15752 14764 15804 14816
rect 16120 14764 16172 14816
rect 19340 14764 19392 14816
rect 19432 14764 19484 14816
rect 20076 14764 20128 14816
rect 21088 14900 21140 14952
rect 21548 14764 21600 14816
rect 22008 14807 22060 14816
rect 22008 14773 22017 14807
rect 22017 14773 22051 14807
rect 22051 14773 22060 14807
rect 22008 14764 22060 14773
rect 22468 14764 22520 14816
rect 23020 14764 23072 14816
rect 3749 14662 3801 14714
rect 3813 14662 3865 14714
rect 3877 14662 3929 14714
rect 3941 14662 3993 14714
rect 4005 14662 4057 14714
rect 9347 14662 9399 14714
rect 9411 14662 9463 14714
rect 9475 14662 9527 14714
rect 9539 14662 9591 14714
rect 9603 14662 9655 14714
rect 14945 14662 14997 14714
rect 15009 14662 15061 14714
rect 15073 14662 15125 14714
rect 15137 14662 15189 14714
rect 15201 14662 15253 14714
rect 20543 14662 20595 14714
rect 20607 14662 20659 14714
rect 20671 14662 20723 14714
rect 20735 14662 20787 14714
rect 20799 14662 20851 14714
rect 5080 14467 5132 14476
rect 5080 14433 5089 14467
rect 5089 14433 5123 14467
rect 5123 14433 5132 14467
rect 5080 14424 5132 14433
rect 5632 14560 5684 14612
rect 5816 14560 5868 14612
rect 7012 14560 7064 14612
rect 8116 14560 8168 14612
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 11612 14603 11664 14612
rect 11612 14569 11621 14603
rect 11621 14569 11655 14603
rect 11655 14569 11664 14603
rect 11612 14560 11664 14569
rect 12808 14560 12860 14612
rect 16948 14603 17000 14612
rect 9680 14492 9732 14544
rect 11888 14492 11940 14544
rect 16212 14535 16264 14544
rect 6920 14356 6972 14408
rect 10324 14356 10376 14408
rect 6644 14288 6696 14340
rect 4896 14220 4948 14272
rect 5080 14220 5132 14272
rect 5816 14220 5868 14272
rect 6460 14220 6512 14272
rect 9772 14288 9824 14340
rect 11428 14288 11480 14340
rect 12440 14356 12492 14408
rect 13360 14424 13412 14476
rect 13728 14467 13780 14476
rect 13728 14433 13737 14467
rect 13737 14433 13771 14467
rect 13771 14433 13780 14467
rect 13728 14424 13780 14433
rect 16212 14501 16221 14535
rect 16221 14501 16255 14535
rect 16255 14501 16264 14535
rect 16212 14492 16264 14501
rect 16948 14569 16957 14603
rect 16957 14569 16991 14603
rect 16991 14569 17000 14603
rect 16948 14560 17000 14569
rect 17592 14560 17644 14612
rect 18144 14560 18196 14612
rect 18788 14603 18840 14612
rect 18788 14569 18797 14603
rect 18797 14569 18831 14603
rect 18831 14569 18840 14603
rect 18788 14560 18840 14569
rect 19432 14560 19484 14612
rect 18880 14535 18932 14544
rect 18880 14501 18889 14535
rect 18889 14501 18923 14535
rect 18923 14501 18932 14535
rect 18880 14492 18932 14501
rect 20444 14560 20496 14612
rect 21088 14492 21140 14544
rect 22744 14492 22796 14544
rect 21272 14467 21324 14476
rect 21272 14433 21281 14467
rect 21281 14433 21315 14467
rect 21315 14433 21324 14467
rect 21272 14424 21324 14433
rect 22468 14467 22520 14476
rect 22468 14433 22477 14467
rect 22477 14433 22511 14467
rect 22511 14433 22520 14467
rect 22468 14424 22520 14433
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 17316 14356 17368 14408
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 10968 14220 11020 14272
rect 11244 14220 11296 14272
rect 11796 14220 11848 14272
rect 12900 14288 12952 14340
rect 13636 14331 13688 14340
rect 13636 14297 13645 14331
rect 13645 14297 13679 14331
rect 13679 14297 13688 14331
rect 13636 14288 13688 14297
rect 15476 14288 15528 14340
rect 14648 14220 14700 14272
rect 15200 14220 15252 14272
rect 15384 14220 15436 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 17224 14288 17276 14340
rect 19156 14356 19208 14408
rect 19524 14399 19576 14408
rect 19524 14365 19558 14399
rect 19558 14365 19576 14399
rect 19524 14356 19576 14365
rect 21456 14356 21508 14408
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 22100 14356 22152 14408
rect 23020 14399 23072 14408
rect 23020 14365 23029 14399
rect 23029 14365 23063 14399
rect 23063 14365 23072 14399
rect 23020 14356 23072 14365
rect 19892 14288 19944 14340
rect 21180 14220 21232 14272
rect 22468 14288 22520 14340
rect 22376 14263 22428 14272
rect 22376 14229 22385 14263
rect 22385 14229 22419 14263
rect 22419 14229 22428 14263
rect 22376 14220 22428 14229
rect 22928 14263 22980 14272
rect 22928 14229 22937 14263
rect 22937 14229 22971 14263
rect 22971 14229 22980 14263
rect 22928 14220 22980 14229
rect 6548 14118 6600 14170
rect 6612 14118 6664 14170
rect 6676 14118 6728 14170
rect 6740 14118 6792 14170
rect 6804 14118 6856 14170
rect 12146 14118 12198 14170
rect 12210 14118 12262 14170
rect 12274 14118 12326 14170
rect 12338 14118 12390 14170
rect 12402 14118 12454 14170
rect 17744 14118 17796 14170
rect 17808 14118 17860 14170
rect 17872 14118 17924 14170
rect 17936 14118 17988 14170
rect 18000 14118 18052 14170
rect 1676 14016 1728 14068
rect 6460 14016 6512 14068
rect 6920 14016 6972 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 11244 14059 11296 14068
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 11336 14016 11388 14068
rect 5080 13948 5132 14000
rect 4344 13923 4396 13932
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 5540 13812 5592 13864
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 5908 13855 5960 13864
rect 5908 13821 5917 13855
rect 5917 13821 5951 13855
rect 5951 13821 5960 13855
rect 5908 13812 5960 13821
rect 6920 13923 6972 13932
rect 6920 13889 6954 13923
rect 6954 13889 6972 13923
rect 8116 13923 8168 13932
rect 6920 13880 6972 13889
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 8392 13923 8444 13932
rect 8392 13889 8426 13923
rect 8426 13889 8444 13923
rect 8392 13880 8444 13889
rect 9772 13948 9824 14000
rect 10876 13948 10928 14000
rect 13636 14016 13688 14068
rect 14648 14059 14700 14068
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 16212 14016 16264 14068
rect 17040 14059 17092 14068
rect 17040 14025 17049 14059
rect 17049 14025 17083 14059
rect 17083 14025 17092 14059
rect 17040 14016 17092 14025
rect 19616 14059 19668 14068
rect 11888 13948 11940 14000
rect 14280 13948 14332 14000
rect 15016 13991 15068 14000
rect 15016 13957 15025 13991
rect 15025 13957 15059 13991
rect 15059 13957 15068 13991
rect 15016 13948 15068 13957
rect 18144 13948 18196 14000
rect 19616 14025 19625 14059
rect 19625 14025 19659 14059
rect 19659 14025 19668 14059
rect 19616 14016 19668 14025
rect 20904 14016 20956 14068
rect 22836 14059 22888 14068
rect 22836 14025 22845 14059
rect 22845 14025 22879 14059
rect 22879 14025 22888 14059
rect 22836 14016 22888 14025
rect 19800 13948 19852 14000
rect 21272 13948 21324 14000
rect 21916 13948 21968 14000
rect 22008 13948 22060 14000
rect 15200 13880 15252 13932
rect 16120 13880 16172 13932
rect 4160 13719 4212 13728
rect 4160 13685 4169 13719
rect 4169 13685 4203 13719
rect 4203 13685 4212 13719
rect 4160 13676 4212 13685
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 14924 13812 14976 13864
rect 16488 13812 16540 13864
rect 15292 13744 15344 13796
rect 16028 13744 16080 13796
rect 16856 13812 16908 13864
rect 16948 13812 17000 13864
rect 17316 13855 17368 13864
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 18512 13923 18564 13932
rect 18512 13889 18546 13923
rect 18546 13889 18564 13923
rect 18144 13812 18196 13864
rect 18512 13880 18564 13889
rect 19984 13923 20036 13932
rect 19984 13889 20018 13923
rect 20018 13889 20036 13923
rect 19984 13880 20036 13889
rect 21456 13880 21508 13932
rect 21916 13855 21968 13864
rect 5264 13676 5316 13685
rect 7012 13676 7064 13728
rect 8024 13719 8076 13728
rect 8024 13685 8033 13719
rect 8033 13685 8067 13719
rect 8067 13685 8076 13719
rect 8024 13676 8076 13685
rect 9220 13676 9272 13728
rect 18604 13676 18656 13728
rect 21548 13787 21600 13796
rect 21548 13753 21557 13787
rect 21557 13753 21591 13787
rect 21591 13753 21600 13787
rect 21548 13744 21600 13753
rect 21916 13821 21925 13855
rect 21925 13821 21959 13855
rect 21959 13821 21968 13855
rect 21916 13812 21968 13821
rect 23848 13812 23900 13864
rect 20076 13676 20128 13728
rect 22008 13676 22060 13728
rect 22560 13719 22612 13728
rect 22560 13685 22569 13719
rect 22569 13685 22603 13719
rect 22603 13685 22612 13719
rect 22560 13676 22612 13685
rect 3749 13574 3801 13626
rect 3813 13574 3865 13626
rect 3877 13574 3929 13626
rect 3941 13574 3993 13626
rect 4005 13574 4057 13626
rect 9347 13574 9399 13626
rect 9411 13574 9463 13626
rect 9475 13574 9527 13626
rect 9539 13574 9591 13626
rect 9603 13574 9655 13626
rect 14945 13574 14997 13626
rect 15009 13574 15061 13626
rect 15073 13574 15125 13626
rect 15137 13574 15189 13626
rect 15201 13574 15253 13626
rect 20543 13574 20595 13626
rect 20607 13574 20659 13626
rect 20671 13574 20723 13626
rect 20735 13574 20787 13626
rect 20799 13574 20851 13626
rect 3424 13472 3476 13524
rect 4344 13472 4396 13524
rect 6920 13472 6972 13524
rect 8116 13515 8168 13524
rect 8116 13481 8125 13515
rect 8125 13481 8159 13515
rect 8159 13481 8168 13515
rect 8116 13472 8168 13481
rect 8300 13472 8352 13524
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 14280 13472 14332 13524
rect 15384 13515 15436 13524
rect 15384 13481 15393 13515
rect 15393 13481 15427 13515
rect 15427 13481 15436 13515
rect 15384 13472 15436 13481
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 18420 13472 18472 13524
rect 4344 13379 4396 13388
rect 4344 13345 4353 13379
rect 4353 13345 4387 13379
rect 4387 13345 4396 13379
rect 4344 13336 4396 13345
rect 4988 13336 5040 13388
rect 5356 13336 5408 13388
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 15108 13447 15160 13456
rect 15108 13413 15117 13447
rect 15117 13413 15151 13447
rect 15151 13413 15160 13447
rect 15108 13404 15160 13413
rect 21640 13472 21692 13524
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 21456 13336 21508 13388
rect 21824 13336 21876 13388
rect 4436 13268 4488 13320
rect 5264 13268 5316 13320
rect 8024 13268 8076 13320
rect 13176 13311 13228 13320
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 7012 13200 7064 13252
rect 8208 13200 8260 13252
rect 8300 13200 8352 13252
rect 9036 13243 9088 13252
rect 9036 13209 9045 13243
rect 9045 13209 9079 13243
rect 9079 13209 9088 13243
rect 9036 13200 9088 13209
rect 10968 13200 11020 13252
rect 4252 13132 4304 13141
rect 5816 13132 5868 13184
rect 9220 13132 9272 13184
rect 9404 13175 9456 13184
rect 9404 13141 9413 13175
rect 9413 13141 9447 13175
rect 9447 13141 9456 13175
rect 9404 13132 9456 13141
rect 10508 13132 10560 13184
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 19340 13268 19392 13320
rect 20076 13268 20128 13320
rect 22560 13336 22612 13388
rect 22928 13379 22980 13388
rect 22928 13345 22937 13379
rect 22937 13345 22971 13379
rect 22971 13345 22980 13379
rect 22928 13336 22980 13345
rect 22192 13268 22244 13320
rect 16028 13243 16080 13252
rect 16028 13209 16062 13243
rect 16062 13209 16080 13243
rect 16028 13200 16080 13209
rect 12808 13132 12860 13184
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 17040 13132 17092 13184
rect 19156 13200 19208 13252
rect 19432 13200 19484 13252
rect 20904 13200 20956 13252
rect 21088 13243 21140 13252
rect 21088 13209 21097 13243
rect 21097 13209 21131 13243
rect 21131 13209 21140 13243
rect 21088 13200 21140 13209
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 19616 13132 19668 13184
rect 19708 13132 19760 13184
rect 21548 13132 21600 13184
rect 6548 13030 6600 13082
rect 6612 13030 6664 13082
rect 6676 13030 6728 13082
rect 6740 13030 6792 13082
rect 6804 13030 6856 13082
rect 12146 13030 12198 13082
rect 12210 13030 12262 13082
rect 12274 13030 12326 13082
rect 12338 13030 12390 13082
rect 12402 13030 12454 13082
rect 17744 13030 17796 13082
rect 17808 13030 17860 13082
rect 17872 13030 17924 13082
rect 17936 13030 17988 13082
rect 18000 13030 18052 13082
rect 3240 12928 3292 12980
rect 4160 12928 4212 12980
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 5172 12928 5224 12980
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 9404 12928 9456 12980
rect 11060 12928 11112 12980
rect 11336 12928 11388 12980
rect 11612 12928 11664 12980
rect 16212 12971 16264 12980
rect 4896 12903 4948 12912
rect 4896 12869 4905 12903
rect 4905 12869 4939 12903
rect 4939 12869 4948 12903
rect 4896 12860 4948 12869
rect 3332 12792 3384 12844
rect 9036 12860 9088 12912
rect 4344 12724 4396 12776
rect 4988 12724 5040 12776
rect 5356 12724 5408 12776
rect 6092 12767 6144 12776
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 6368 12724 6420 12776
rect 9404 12792 9456 12844
rect 4896 12588 4948 12640
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 8392 12588 8444 12640
rect 10784 12656 10836 12708
rect 11060 12699 11112 12708
rect 11060 12665 11069 12699
rect 11069 12665 11103 12699
rect 11103 12665 11112 12699
rect 11060 12656 11112 12665
rect 12808 12860 12860 12912
rect 16212 12937 16221 12971
rect 16221 12937 16255 12971
rect 16255 12937 16264 12971
rect 16212 12928 16264 12937
rect 17316 12928 17368 12980
rect 18328 12971 18380 12980
rect 18328 12937 18337 12971
rect 18337 12937 18371 12971
rect 18371 12937 18380 12971
rect 18328 12928 18380 12937
rect 11796 12792 11848 12844
rect 16304 12860 16356 12912
rect 16488 12860 16540 12912
rect 13820 12792 13872 12844
rect 14280 12792 14332 12844
rect 15384 12792 15436 12844
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 22376 12928 22428 12980
rect 19340 12792 19392 12844
rect 20352 12792 20404 12844
rect 18604 12724 18656 12776
rect 21640 12792 21692 12844
rect 22008 12792 22060 12844
rect 23112 12835 23164 12844
rect 23112 12801 23121 12835
rect 23121 12801 23155 12835
rect 23155 12801 23164 12835
rect 23112 12792 23164 12801
rect 11428 12588 11480 12640
rect 12716 12656 12768 12708
rect 16028 12699 16080 12708
rect 16028 12665 16037 12699
rect 16037 12665 16071 12699
rect 16071 12665 16080 12699
rect 16028 12656 16080 12665
rect 19984 12656 20036 12708
rect 12164 12588 12216 12640
rect 15384 12588 15436 12640
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 17132 12588 17184 12640
rect 18420 12588 18472 12640
rect 19064 12588 19116 12640
rect 22008 12588 22060 12640
rect 22928 12631 22980 12640
rect 22928 12597 22937 12631
rect 22937 12597 22971 12631
rect 22971 12597 22980 12631
rect 22928 12588 22980 12597
rect 3749 12486 3801 12538
rect 3813 12486 3865 12538
rect 3877 12486 3929 12538
rect 3941 12486 3993 12538
rect 4005 12486 4057 12538
rect 9347 12486 9399 12538
rect 9411 12486 9463 12538
rect 9475 12486 9527 12538
rect 9539 12486 9591 12538
rect 9603 12486 9655 12538
rect 14945 12486 14997 12538
rect 15009 12486 15061 12538
rect 15073 12486 15125 12538
rect 15137 12486 15189 12538
rect 15201 12486 15253 12538
rect 20543 12486 20595 12538
rect 20607 12486 20659 12538
rect 20671 12486 20723 12538
rect 20735 12486 20787 12538
rect 20799 12486 20851 12538
rect 6368 12384 6420 12436
rect 8392 12384 8444 12436
rect 5080 12248 5132 12300
rect 6000 12248 6052 12300
rect 10508 12384 10560 12436
rect 11612 12384 11664 12436
rect 12164 12427 12216 12436
rect 5448 12112 5500 12164
rect 6460 12112 6512 12164
rect 8944 12180 8996 12232
rect 10784 12316 10836 12368
rect 12164 12393 12173 12427
rect 12173 12393 12207 12427
rect 12207 12393 12216 12427
rect 12164 12384 12216 12393
rect 12808 12384 12860 12436
rect 13912 12384 13964 12436
rect 16580 12427 16632 12436
rect 12256 12316 12308 12368
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 12164 12248 12216 12300
rect 14280 12316 14332 12368
rect 15108 12316 15160 12368
rect 12716 12291 12768 12300
rect 12716 12257 12725 12291
rect 12725 12257 12759 12291
rect 12759 12257 12768 12291
rect 12716 12248 12768 12257
rect 13728 12248 13780 12300
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 16488 12359 16540 12368
rect 16488 12325 16497 12359
rect 16497 12325 16531 12359
rect 16531 12325 16540 12359
rect 16488 12316 16540 12325
rect 18512 12384 18564 12436
rect 21456 12427 21508 12436
rect 13176 12180 13228 12232
rect 7196 12112 7248 12164
rect 8024 12112 8076 12164
rect 3148 12044 3200 12096
rect 4988 12044 5040 12096
rect 7012 12044 7064 12096
rect 10416 12112 10468 12164
rect 12256 12112 12308 12164
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 15108 12180 15160 12189
rect 16856 12248 16908 12300
rect 17960 12248 18012 12300
rect 17224 12180 17276 12232
rect 18328 12180 18380 12232
rect 18604 12223 18656 12232
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 21456 12393 21465 12427
rect 21465 12393 21499 12427
rect 21499 12393 21508 12427
rect 21456 12384 21508 12393
rect 21916 12384 21968 12436
rect 21364 12248 21416 12300
rect 18604 12180 18656 12189
rect 15476 12112 15528 12164
rect 16488 12112 16540 12164
rect 18696 12112 18748 12164
rect 19340 12180 19392 12232
rect 19984 12180 20036 12232
rect 19616 12112 19668 12164
rect 11980 12044 12032 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 16948 12044 17000 12096
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 17408 12044 17460 12096
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 18236 12044 18288 12096
rect 18788 12087 18840 12096
rect 18788 12053 18797 12087
rect 18797 12053 18831 12087
rect 18831 12053 18840 12087
rect 18788 12044 18840 12053
rect 19800 12044 19852 12096
rect 20260 12044 20312 12096
rect 21732 12180 21784 12232
rect 22652 12316 22704 12368
rect 22928 12316 22980 12368
rect 22192 12291 22244 12300
rect 22192 12257 22201 12291
rect 22201 12257 22235 12291
rect 22235 12257 22244 12291
rect 22192 12248 22244 12257
rect 22376 12248 22428 12300
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 22008 12180 22060 12232
rect 22744 12180 22796 12232
rect 21640 12112 21692 12164
rect 22008 12087 22060 12096
rect 22008 12053 22017 12087
rect 22017 12053 22051 12087
rect 22051 12053 22060 12087
rect 22008 12044 22060 12053
rect 22560 12044 22612 12096
rect 22744 12087 22796 12096
rect 22744 12053 22753 12087
rect 22753 12053 22787 12087
rect 22787 12053 22796 12087
rect 22744 12044 22796 12053
rect 6548 11942 6600 11994
rect 6612 11942 6664 11994
rect 6676 11942 6728 11994
rect 6740 11942 6792 11994
rect 6804 11942 6856 11994
rect 12146 11942 12198 11994
rect 12210 11942 12262 11994
rect 12274 11942 12326 11994
rect 12338 11942 12390 11994
rect 12402 11942 12454 11994
rect 17744 11942 17796 11994
rect 17808 11942 17860 11994
rect 17872 11942 17924 11994
rect 17936 11942 17988 11994
rect 18000 11942 18052 11994
rect 3332 11883 3384 11892
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 3332 11840 3384 11849
rect 4252 11840 4304 11892
rect 4528 11840 4580 11892
rect 4896 11883 4948 11892
rect 4896 11849 4905 11883
rect 4905 11849 4939 11883
rect 4939 11849 4948 11883
rect 4896 11840 4948 11849
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 5448 11883 5500 11892
rect 4988 11840 5040 11849
rect 5448 11849 5457 11883
rect 5457 11849 5491 11883
rect 5491 11849 5500 11883
rect 5448 11840 5500 11849
rect 6460 11840 6512 11892
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 11796 11840 11848 11892
rect 13176 11840 13228 11892
rect 13544 11840 13596 11892
rect 14280 11883 14332 11892
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 14372 11840 14424 11892
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 15660 11840 15712 11892
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 16672 11840 16724 11892
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 18328 11883 18380 11892
rect 18328 11849 18337 11883
rect 18337 11849 18371 11883
rect 18371 11849 18380 11883
rect 18328 11840 18380 11849
rect 18604 11840 18656 11892
rect 19984 11840 20036 11892
rect 20352 11840 20404 11892
rect 21088 11840 21140 11892
rect 4160 11772 4212 11824
rect 4344 11772 4396 11824
rect 7380 11772 7432 11824
rect 11336 11772 11388 11824
rect 12992 11772 13044 11824
rect 13268 11772 13320 11824
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 3148 11704 3200 11713
rect 3608 11704 3660 11756
rect 4252 11704 4304 11756
rect 10324 11704 10376 11756
rect 12808 11704 12860 11756
rect 13084 11704 13136 11756
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 4160 11636 4212 11688
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 6092 11679 6144 11688
rect 6092 11645 6101 11679
rect 6101 11645 6135 11679
rect 6135 11645 6144 11679
rect 6092 11636 6144 11645
rect 11520 11679 11572 11688
rect 8024 11500 8076 11552
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 15936 11772 15988 11824
rect 13636 11704 13688 11756
rect 13728 11636 13780 11688
rect 16212 11704 16264 11756
rect 18236 11772 18288 11824
rect 18788 11772 18840 11824
rect 20996 11772 21048 11824
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17960 11704 18012 11756
rect 11796 11500 11848 11552
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 16948 11636 17000 11688
rect 18328 11704 18380 11756
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 19248 11704 19300 11756
rect 21640 11772 21692 11824
rect 22284 11772 22336 11824
rect 22652 11815 22704 11824
rect 22652 11781 22661 11815
rect 22661 11781 22695 11815
rect 22695 11781 22704 11815
rect 22652 11772 22704 11781
rect 16764 11500 16816 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 18604 11543 18656 11552
rect 18604 11509 18613 11543
rect 18613 11509 18647 11543
rect 18647 11509 18656 11543
rect 18604 11500 18656 11509
rect 21272 11747 21324 11756
rect 21272 11713 21290 11747
rect 21290 11713 21324 11747
rect 21548 11747 21600 11756
rect 21272 11704 21324 11713
rect 21548 11713 21557 11747
rect 21557 11713 21591 11747
rect 21591 11713 21600 11747
rect 21548 11704 21600 11713
rect 20352 11500 20404 11552
rect 21640 11500 21692 11552
rect 22376 11679 22428 11688
rect 22376 11645 22385 11679
rect 22385 11645 22419 11679
rect 22419 11645 22428 11679
rect 22376 11636 22428 11645
rect 22560 11500 22612 11552
rect 3749 11398 3801 11450
rect 3813 11398 3865 11450
rect 3877 11398 3929 11450
rect 3941 11398 3993 11450
rect 4005 11398 4057 11450
rect 9347 11398 9399 11450
rect 9411 11398 9463 11450
rect 9475 11398 9527 11450
rect 9539 11398 9591 11450
rect 9603 11398 9655 11450
rect 14945 11398 14997 11450
rect 15009 11398 15061 11450
rect 15073 11398 15125 11450
rect 15137 11398 15189 11450
rect 15201 11398 15253 11450
rect 20543 11398 20595 11450
rect 20607 11398 20659 11450
rect 20671 11398 20723 11450
rect 20735 11398 20787 11450
rect 20799 11398 20851 11450
rect 7196 11339 7248 11348
rect 7196 11305 7205 11339
rect 7205 11305 7239 11339
rect 7239 11305 7248 11339
rect 7196 11296 7248 11305
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 11980 11339 12032 11348
rect 11980 11305 11989 11339
rect 11989 11305 12023 11339
rect 12023 11305 12032 11339
rect 11980 11296 12032 11305
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 16856 11296 16908 11348
rect 17040 11296 17092 11348
rect 17960 11296 18012 11348
rect 19248 11339 19300 11348
rect 5724 11271 5776 11280
rect 5724 11237 5733 11271
rect 5733 11237 5767 11271
rect 5767 11237 5776 11271
rect 5724 11228 5776 11237
rect 10324 11271 10376 11280
rect 10324 11237 10333 11271
rect 10333 11237 10367 11271
rect 10367 11237 10376 11271
rect 10324 11228 10376 11237
rect 4344 11160 4396 11212
rect 4712 11160 4764 11212
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 8024 11092 8076 11144
rect 9680 11092 9732 11144
rect 12072 11092 12124 11144
rect 13452 11160 13504 11212
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19064 11228 19116 11280
rect 19340 11228 19392 11280
rect 15108 11160 15160 11212
rect 15660 11160 15712 11212
rect 17316 11160 17368 11212
rect 14648 11092 14700 11144
rect 5448 11024 5500 11076
rect 6460 11024 6512 11076
rect 7012 11024 7064 11076
rect 11980 11024 12032 11076
rect 13084 11067 13136 11076
rect 13084 11033 13102 11067
rect 13102 11033 13136 11067
rect 13084 11024 13136 11033
rect 16672 11024 16724 11076
rect 19340 11092 19392 11144
rect 20352 11135 20404 11144
rect 20352 11101 20370 11135
rect 20370 11101 20404 11135
rect 20628 11135 20680 11144
rect 20352 11092 20404 11101
rect 17592 11067 17644 11076
rect 17592 11033 17601 11067
rect 17601 11033 17635 11067
rect 17635 11033 17644 11067
rect 17592 11024 17644 11033
rect 19248 11024 19300 11076
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 20628 11092 20680 11101
rect 22008 11296 22060 11348
rect 22284 11271 22336 11280
rect 22284 11237 22293 11271
rect 22293 11237 22327 11271
rect 22327 11237 22336 11271
rect 22284 11228 22336 11237
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 22836 11203 22888 11212
rect 22836 11169 22845 11203
rect 22845 11169 22879 11203
rect 22879 11169 22888 11203
rect 22836 11160 22888 11169
rect 23020 11203 23072 11212
rect 23020 11169 23029 11203
rect 23029 11169 23063 11203
rect 23063 11169 23072 11203
rect 23020 11160 23072 11169
rect 21364 11092 21416 11144
rect 21272 11024 21324 11076
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 4528 10956 4580 11008
rect 4988 10956 5040 11008
rect 7748 10956 7800 11008
rect 10324 10956 10376 11008
rect 18512 10956 18564 11008
rect 18972 10956 19024 11008
rect 19156 10956 19208 11008
rect 22376 10999 22428 11008
rect 22376 10965 22385 10999
rect 22385 10965 22419 10999
rect 22419 10965 22428 10999
rect 22376 10956 22428 10965
rect 6548 10854 6600 10906
rect 6612 10854 6664 10906
rect 6676 10854 6728 10906
rect 6740 10854 6792 10906
rect 6804 10854 6856 10906
rect 12146 10854 12198 10906
rect 12210 10854 12262 10906
rect 12274 10854 12326 10906
rect 12338 10854 12390 10906
rect 12402 10854 12454 10906
rect 17744 10854 17796 10906
rect 17808 10854 17860 10906
rect 17872 10854 17924 10906
rect 17936 10854 17988 10906
rect 18000 10854 18052 10906
rect 4344 10752 4396 10804
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 4988 10752 5040 10761
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 6828 10684 6880 10736
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 7932 10727 7984 10736
rect 7932 10693 7950 10727
rect 7950 10693 7984 10727
rect 7932 10684 7984 10693
rect 8116 10684 8168 10736
rect 11796 10727 11848 10736
rect 11796 10693 11830 10727
rect 11830 10693 11848 10727
rect 11796 10684 11848 10693
rect 13084 10752 13136 10804
rect 13268 10795 13320 10804
rect 13268 10761 13277 10795
rect 13277 10761 13311 10795
rect 13311 10761 13320 10795
rect 13268 10752 13320 10761
rect 14832 10752 14884 10804
rect 15108 10752 15160 10804
rect 22560 10795 22612 10804
rect 15384 10684 15436 10736
rect 10508 10659 10560 10668
rect 4712 10548 4764 10600
rect 4252 10480 4304 10532
rect 5080 10480 5132 10532
rect 6828 10523 6880 10532
rect 6828 10489 6837 10523
rect 6837 10489 6871 10523
rect 6871 10489 6880 10523
rect 6828 10480 6880 10489
rect 5908 10412 5960 10464
rect 7104 10412 7156 10464
rect 8208 10412 8260 10464
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 12072 10616 12124 10668
rect 13636 10616 13688 10668
rect 13452 10548 13504 10600
rect 13820 10616 13872 10668
rect 15660 10616 15712 10668
rect 16120 10659 16172 10668
rect 16120 10625 16138 10659
rect 16138 10625 16172 10659
rect 16120 10616 16172 10625
rect 17224 10616 17276 10668
rect 19432 10684 19484 10736
rect 20628 10684 20680 10736
rect 21548 10727 21600 10736
rect 21548 10693 21557 10727
rect 21557 10693 21591 10727
rect 21591 10693 21600 10727
rect 21548 10684 21600 10693
rect 19156 10616 19208 10668
rect 20352 10659 20404 10668
rect 20352 10625 20386 10659
rect 20386 10625 20404 10659
rect 22560 10761 22569 10795
rect 22569 10761 22603 10795
rect 22603 10761 22612 10795
rect 22560 10752 22612 10761
rect 22100 10727 22152 10736
rect 22100 10693 22109 10727
rect 22109 10693 22143 10727
rect 22143 10693 22152 10727
rect 22100 10684 22152 10693
rect 23388 10684 23440 10736
rect 20352 10616 20404 10625
rect 21732 10548 21784 10600
rect 22284 10616 22336 10668
rect 10508 10412 10560 10464
rect 13176 10412 13228 10464
rect 13360 10412 13412 10464
rect 19800 10412 19852 10464
rect 21272 10412 21324 10464
rect 21456 10455 21508 10464
rect 21456 10421 21465 10455
rect 21465 10421 21499 10455
rect 21499 10421 21508 10455
rect 21456 10412 21508 10421
rect 21548 10412 21600 10464
rect 22100 10412 22152 10464
rect 3749 10310 3801 10362
rect 3813 10310 3865 10362
rect 3877 10310 3929 10362
rect 3941 10310 3993 10362
rect 4005 10310 4057 10362
rect 9347 10310 9399 10362
rect 9411 10310 9463 10362
rect 9475 10310 9527 10362
rect 9539 10310 9591 10362
rect 9603 10310 9655 10362
rect 14945 10310 14997 10362
rect 15009 10310 15061 10362
rect 15073 10310 15125 10362
rect 15137 10310 15189 10362
rect 15201 10310 15253 10362
rect 20543 10310 20595 10362
rect 20607 10310 20659 10362
rect 20671 10310 20723 10362
rect 20735 10310 20787 10362
rect 20799 10310 20851 10362
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 4620 10208 4672 10260
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 10508 10251 10560 10260
rect 7288 10208 7340 10217
rect 4160 10072 4212 10124
rect 5356 10072 5408 10124
rect 5908 10115 5960 10124
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 5908 10072 5960 10081
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 5080 10004 5132 10056
rect 3792 9936 3844 9988
rect 4436 9936 4488 9988
rect 6184 9979 6236 9988
rect 6184 9945 6218 9979
rect 6218 9945 6236 9979
rect 6184 9936 6236 9945
rect 8208 10004 8260 10056
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 10324 10140 10376 10192
rect 11612 10072 11664 10124
rect 13176 10140 13228 10192
rect 13820 10183 13872 10192
rect 13360 10072 13412 10124
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 13820 10149 13829 10183
rect 13829 10149 13863 10183
rect 13863 10149 13872 10183
rect 13820 10140 13872 10149
rect 15384 10140 15436 10192
rect 15660 10183 15712 10192
rect 15660 10149 15669 10183
rect 15669 10149 15703 10183
rect 15703 10149 15712 10183
rect 15660 10140 15712 10149
rect 16120 10140 16172 10192
rect 18420 10140 18472 10192
rect 10508 10004 10560 10056
rect 12992 10004 13044 10056
rect 13820 10004 13872 10056
rect 16856 10072 16908 10124
rect 17040 10004 17092 10056
rect 20352 10208 20404 10260
rect 3516 9868 3568 9920
rect 5080 9911 5132 9920
rect 5080 9877 5089 9911
rect 5089 9877 5123 9911
rect 5123 9877 5132 9911
rect 5080 9868 5132 9877
rect 6460 9868 6512 9920
rect 12072 9868 12124 9920
rect 13268 9936 13320 9988
rect 18328 9936 18380 9988
rect 19340 10004 19392 10056
rect 19524 10047 19576 10056
rect 19524 10013 19558 10047
rect 19558 10013 19576 10047
rect 19524 10004 19576 10013
rect 19800 10004 19852 10056
rect 20720 10183 20772 10192
rect 20720 10149 20729 10183
rect 20729 10149 20763 10183
rect 20763 10149 20772 10183
rect 20720 10140 20772 10149
rect 21456 10004 21508 10056
rect 22100 10047 22152 10056
rect 22100 10013 22109 10047
rect 22109 10013 22143 10047
rect 22143 10013 22152 10047
rect 22652 10047 22704 10056
rect 22100 10004 22152 10013
rect 13360 9911 13412 9920
rect 13360 9877 13369 9911
rect 13369 9877 13403 9911
rect 13403 9877 13412 9911
rect 13360 9868 13412 9877
rect 13452 9911 13504 9920
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 16948 9911 17000 9920
rect 13452 9868 13504 9877
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17132 9868 17184 9920
rect 17224 9868 17276 9920
rect 22284 9936 22336 9988
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 20444 9868 20496 9920
rect 22008 9868 22060 9920
rect 22100 9868 22152 9920
rect 22376 9868 22428 9920
rect 23480 9868 23532 9920
rect 6548 9766 6600 9818
rect 6612 9766 6664 9818
rect 6676 9766 6728 9818
rect 6740 9766 6792 9818
rect 6804 9766 6856 9818
rect 12146 9766 12198 9818
rect 12210 9766 12262 9818
rect 12274 9766 12326 9818
rect 12338 9766 12390 9818
rect 12402 9766 12454 9818
rect 17744 9766 17796 9818
rect 17808 9766 17860 9818
rect 17872 9766 17924 9818
rect 17936 9766 17988 9818
rect 18000 9766 18052 9818
rect 3516 9707 3568 9716
rect 3516 9673 3525 9707
rect 3525 9673 3559 9707
rect 3559 9673 3568 9707
rect 3516 9664 3568 9673
rect 3792 9707 3844 9716
rect 3792 9673 3801 9707
rect 3801 9673 3835 9707
rect 3835 9673 3844 9707
rect 3792 9664 3844 9673
rect 6920 9664 6972 9716
rect 7932 9664 7984 9716
rect 7288 9596 7340 9648
rect 7380 9596 7432 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 4528 9528 4580 9580
rect 6184 9528 6236 9580
rect 6644 9528 6696 9580
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 6276 9392 6328 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3148 9324 3200 9376
rect 4436 9324 4488 9376
rect 6460 9324 6512 9376
rect 10508 9664 10560 9716
rect 11796 9664 11848 9716
rect 13268 9707 13320 9716
rect 13268 9673 13277 9707
rect 13277 9673 13311 9707
rect 13311 9673 13320 9707
rect 13268 9664 13320 9673
rect 13360 9664 13412 9716
rect 15660 9664 15712 9716
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 9036 9324 9088 9376
rect 17040 9664 17092 9716
rect 19340 9664 19392 9716
rect 13452 9528 13504 9580
rect 15476 9528 15528 9580
rect 17040 9528 17092 9580
rect 17500 9528 17552 9580
rect 17776 9528 17828 9580
rect 18972 9596 19024 9648
rect 19156 9596 19208 9648
rect 21272 9664 21324 9716
rect 19616 9596 19668 9648
rect 13360 9460 13412 9512
rect 17224 9460 17276 9512
rect 19984 9571 20036 9580
rect 19984 9537 20002 9571
rect 20002 9537 20036 9571
rect 19984 9528 20036 9537
rect 18972 9460 19024 9512
rect 22100 9596 22152 9648
rect 22836 9639 22888 9648
rect 22836 9605 22845 9639
rect 22845 9605 22879 9639
rect 22879 9605 22888 9639
rect 22836 9596 22888 9605
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 21088 9460 21140 9512
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 11336 9324 11388 9376
rect 13544 9324 13596 9376
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 17776 9324 17828 9376
rect 18972 9324 19024 9376
rect 19340 9324 19392 9376
rect 20260 9324 20312 9376
rect 22284 9460 22336 9512
rect 22652 9324 22704 9376
rect 23020 9367 23072 9376
rect 23020 9333 23029 9367
rect 23029 9333 23063 9367
rect 23063 9333 23072 9367
rect 23020 9324 23072 9333
rect 3749 9222 3801 9274
rect 3813 9222 3865 9274
rect 3877 9222 3929 9274
rect 3941 9222 3993 9274
rect 4005 9222 4057 9274
rect 9347 9222 9399 9274
rect 9411 9222 9463 9274
rect 9475 9222 9527 9274
rect 9539 9222 9591 9274
rect 9603 9222 9655 9274
rect 14945 9222 14997 9274
rect 15009 9222 15061 9274
rect 15073 9222 15125 9274
rect 15137 9222 15189 9274
rect 15201 9222 15253 9274
rect 20543 9222 20595 9274
rect 20607 9222 20659 9274
rect 20671 9222 20723 9274
rect 20735 9222 20787 9274
rect 20799 9222 20851 9274
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 4344 9120 4396 9172
rect 5356 9120 5408 9172
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 10876 9120 10928 9172
rect 13820 9163 13872 9172
rect 13820 9129 13829 9163
rect 13829 9129 13863 9163
rect 13863 9129 13872 9163
rect 13820 9120 13872 9129
rect 3332 9052 3384 9104
rect 4160 9052 4212 9104
rect 3148 9027 3200 9036
rect 3148 8993 3157 9027
rect 3157 8993 3191 9027
rect 3191 8993 3200 9027
rect 3148 8984 3200 8993
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 6644 9052 6696 9104
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 16212 9120 16264 9172
rect 18604 9120 18656 9172
rect 20260 9120 20312 9172
rect 20628 9120 20680 9172
rect 22100 9120 22152 9172
rect 19064 9095 19116 9104
rect 19064 9061 19073 9095
rect 19073 9061 19107 9095
rect 19107 9061 19116 9095
rect 19064 9052 19116 9061
rect 23204 9052 23256 9104
rect 19432 8984 19484 9036
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 22744 9027 22796 9036
rect 22744 8993 22753 9027
rect 22753 8993 22787 9027
rect 22787 8993 22796 9027
rect 22744 8984 22796 8993
rect 4160 8916 4212 8968
rect 5080 8916 5132 8968
rect 6920 8916 6972 8968
rect 4528 8848 4580 8900
rect 5724 8848 5776 8900
rect 3240 8823 3292 8832
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 4436 8780 4488 8832
rect 4896 8780 4948 8832
rect 7288 8780 7340 8832
rect 10048 8916 10100 8968
rect 10600 8916 10652 8968
rect 14832 8959 14884 8968
rect 14832 8925 14866 8959
rect 14866 8925 14884 8959
rect 14832 8916 14884 8925
rect 18144 8916 18196 8968
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 11428 8780 11480 8789
rect 16120 8780 16172 8832
rect 17960 8848 18012 8900
rect 18328 8848 18380 8900
rect 18236 8780 18288 8832
rect 20260 8848 20312 8900
rect 21088 8916 21140 8968
rect 23020 8916 23072 8968
rect 20444 8848 20496 8900
rect 20536 8848 20588 8900
rect 19800 8780 19852 8832
rect 19892 8780 19944 8832
rect 20628 8780 20680 8832
rect 21824 8891 21876 8900
rect 21824 8857 21842 8891
rect 21842 8857 21876 8891
rect 22560 8891 22612 8900
rect 21824 8848 21876 8857
rect 22560 8857 22569 8891
rect 22569 8857 22603 8891
rect 22603 8857 22612 8891
rect 22560 8848 22612 8857
rect 23020 8823 23072 8832
rect 23020 8789 23029 8823
rect 23029 8789 23063 8823
rect 23063 8789 23072 8823
rect 23020 8780 23072 8789
rect 6548 8678 6600 8730
rect 6612 8678 6664 8730
rect 6676 8678 6728 8730
rect 6740 8678 6792 8730
rect 6804 8678 6856 8730
rect 12146 8678 12198 8730
rect 12210 8678 12262 8730
rect 12274 8678 12326 8730
rect 12338 8678 12390 8730
rect 12402 8678 12454 8730
rect 17744 8678 17796 8730
rect 17808 8678 17860 8730
rect 17872 8678 17924 8730
rect 17936 8678 17988 8730
rect 18000 8678 18052 8730
rect 3700 8576 3752 8628
rect 4896 8576 4948 8628
rect 6184 8619 6236 8628
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 6920 8576 6972 8628
rect 10600 8576 10652 8628
rect 16764 8576 16816 8628
rect 18420 8576 18472 8628
rect 19156 8576 19208 8628
rect 19524 8619 19576 8628
rect 19524 8585 19533 8619
rect 19533 8585 19567 8619
rect 19567 8585 19576 8619
rect 19524 8576 19576 8585
rect 20352 8576 20404 8628
rect 4436 8508 4488 8560
rect 3608 8440 3660 8492
rect 6460 8508 6512 8560
rect 3884 8372 3936 8424
rect 3424 8304 3476 8356
rect 3700 8304 3752 8356
rect 4160 8415 4212 8424
rect 4160 8381 4169 8415
rect 4169 8381 4203 8415
rect 4203 8381 4212 8415
rect 8484 8508 8536 8560
rect 10048 8508 10100 8560
rect 4160 8372 4212 8381
rect 4252 8304 4304 8356
rect 7104 8483 7156 8492
rect 7104 8449 7138 8483
rect 7138 8449 7156 8483
rect 7104 8440 7156 8449
rect 4344 8236 4396 8288
rect 8116 8304 8168 8356
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 10692 8440 10744 8492
rect 11520 8440 11572 8492
rect 16120 8440 16172 8492
rect 16764 8440 16816 8492
rect 17040 8508 17092 8560
rect 19248 8440 19300 8492
rect 6460 8279 6512 8288
rect 6460 8245 6469 8279
rect 6469 8245 6503 8279
rect 6503 8245 6512 8279
rect 6460 8236 6512 8245
rect 15936 8347 15988 8356
rect 15936 8313 15945 8347
rect 15945 8313 15979 8347
rect 15979 8313 15988 8347
rect 15936 8304 15988 8313
rect 18144 8415 18196 8424
rect 18144 8381 18153 8415
rect 18153 8381 18187 8415
rect 18187 8381 18196 8415
rect 18144 8372 18196 8381
rect 19156 8372 19208 8424
rect 21180 8483 21232 8492
rect 21180 8449 21189 8483
rect 21189 8449 21223 8483
rect 21223 8449 21232 8483
rect 21180 8440 21232 8449
rect 21548 8440 21600 8492
rect 22008 8440 22060 8492
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 22284 8415 22336 8424
rect 22284 8381 22293 8415
rect 22293 8381 22327 8415
rect 22327 8381 22336 8415
rect 22284 8372 22336 8381
rect 19616 8236 19668 8288
rect 20260 8236 20312 8288
rect 20628 8236 20680 8288
rect 21272 8304 21324 8356
rect 21824 8347 21876 8356
rect 21824 8313 21833 8347
rect 21833 8313 21867 8347
rect 21867 8313 21876 8347
rect 21824 8304 21876 8313
rect 22100 8236 22152 8288
rect 23572 8372 23624 8424
rect 3749 8134 3801 8186
rect 3813 8134 3865 8186
rect 3877 8134 3929 8186
rect 3941 8134 3993 8186
rect 4005 8134 4057 8186
rect 9347 8134 9399 8186
rect 9411 8134 9463 8186
rect 9475 8134 9527 8186
rect 9539 8134 9591 8186
rect 9603 8134 9655 8186
rect 14945 8134 14997 8186
rect 15009 8134 15061 8186
rect 15073 8134 15125 8186
rect 15137 8134 15189 8186
rect 15201 8134 15253 8186
rect 20543 8134 20595 8186
rect 20607 8134 20659 8186
rect 20671 8134 20723 8186
rect 20735 8134 20787 8186
rect 20799 8134 20851 8186
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 19524 7964 19576 8016
rect 9680 7896 9732 7948
rect 11336 7896 11388 7948
rect 20996 8032 21048 8084
rect 21088 7964 21140 8016
rect 5540 7828 5592 7880
rect 5356 7760 5408 7812
rect 6920 7760 6972 7812
rect 5724 7692 5776 7744
rect 5908 7735 5960 7744
rect 5908 7701 5917 7735
rect 5917 7701 5951 7735
rect 5951 7701 5960 7735
rect 8484 7803 8536 7812
rect 8484 7769 8502 7803
rect 8502 7769 8536 7803
rect 8484 7760 8536 7769
rect 5908 7692 5960 7701
rect 8668 7692 8720 7744
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 11428 7828 11480 7880
rect 14648 7828 14700 7880
rect 16212 7828 16264 7880
rect 12808 7803 12860 7812
rect 12808 7769 12842 7803
rect 12842 7769 12860 7803
rect 12808 7760 12860 7769
rect 12900 7760 12952 7812
rect 18880 7828 18932 7880
rect 21180 7896 21232 7948
rect 21732 7939 21784 7948
rect 21732 7905 21744 7939
rect 21744 7905 21778 7939
rect 21778 7905 21784 7939
rect 21732 7896 21784 7905
rect 20260 7760 20312 7812
rect 8944 7692 8996 7701
rect 11152 7735 11204 7744
rect 11152 7701 11161 7735
rect 11161 7701 11195 7735
rect 11195 7701 11204 7735
rect 11152 7692 11204 7701
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 12072 7692 12124 7744
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 16764 7692 16816 7744
rect 16948 7735 17000 7744
rect 16948 7701 16957 7735
rect 16957 7701 16991 7735
rect 16991 7701 17000 7735
rect 16948 7692 17000 7701
rect 17040 7735 17092 7744
rect 17040 7701 17049 7735
rect 17049 7701 17083 7735
rect 17083 7701 17092 7735
rect 17040 7692 17092 7701
rect 18052 7692 18104 7744
rect 18328 7692 18380 7744
rect 18696 7692 18748 7744
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 19616 7692 19668 7744
rect 21364 7828 21416 7880
rect 22376 7828 22428 7880
rect 20812 7760 20864 7812
rect 22008 7692 22060 7744
rect 23112 7735 23164 7744
rect 23112 7701 23121 7735
rect 23121 7701 23155 7735
rect 23155 7701 23164 7735
rect 23112 7692 23164 7701
rect 6548 7590 6600 7642
rect 6612 7590 6664 7642
rect 6676 7590 6728 7642
rect 6740 7590 6792 7642
rect 6804 7590 6856 7642
rect 12146 7590 12198 7642
rect 12210 7590 12262 7642
rect 12274 7590 12326 7642
rect 12338 7590 12390 7642
rect 12402 7590 12454 7642
rect 17744 7590 17796 7642
rect 17808 7590 17860 7642
rect 17872 7590 17924 7642
rect 17936 7590 17988 7642
rect 18000 7590 18052 7642
rect 3240 7488 3292 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 9680 7488 9732 7540
rect 11428 7488 11480 7540
rect 13452 7488 13504 7540
rect 14464 7488 14516 7540
rect 17960 7488 18012 7540
rect 18236 7488 18288 7540
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 21640 7488 21692 7540
rect 22100 7531 22152 7540
rect 22100 7497 22109 7531
rect 22109 7497 22143 7531
rect 22143 7497 22152 7531
rect 22100 7488 22152 7497
rect 22284 7488 22336 7540
rect 5540 7420 5592 7472
rect 6460 7463 6512 7472
rect 6460 7429 6469 7463
rect 6469 7429 6503 7463
rect 6503 7429 6512 7463
rect 6460 7420 6512 7429
rect 4344 7284 4396 7336
rect 5632 7352 5684 7404
rect 8944 7420 8996 7472
rect 9864 7420 9916 7472
rect 13912 7420 13964 7472
rect 14556 7420 14608 7472
rect 17040 7420 17092 7472
rect 18788 7420 18840 7472
rect 19432 7420 19484 7472
rect 22836 7463 22888 7472
rect 22836 7429 22845 7463
rect 22845 7429 22879 7463
rect 22879 7429 22888 7463
rect 22836 7420 22888 7429
rect 5816 7284 5868 7336
rect 8760 7395 8812 7404
rect 8760 7361 8794 7395
rect 8794 7361 8812 7395
rect 8760 7352 8812 7361
rect 10232 7395 10284 7404
rect 10232 7361 10266 7395
rect 10266 7361 10284 7395
rect 10232 7352 10284 7361
rect 11796 7352 11848 7404
rect 11980 7395 12032 7404
rect 11980 7361 12014 7395
rect 12014 7361 12032 7395
rect 11980 7352 12032 7361
rect 15936 7352 15988 7404
rect 18880 7352 18932 7404
rect 14648 7284 14700 7336
rect 19616 7327 19668 7336
rect 8760 7148 8812 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 14280 7148 14332 7200
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 18144 7259 18196 7268
rect 18144 7225 18153 7259
rect 18153 7225 18187 7259
rect 18187 7225 18196 7259
rect 18144 7216 18196 7225
rect 22284 7352 22336 7404
rect 22928 7352 22980 7404
rect 21824 7284 21876 7336
rect 17592 7148 17644 7200
rect 19156 7148 19208 7200
rect 21456 7148 21508 7200
rect 22100 7216 22152 7268
rect 22652 7259 22704 7268
rect 22652 7225 22661 7259
rect 22661 7225 22695 7259
rect 22695 7225 22704 7259
rect 22652 7216 22704 7225
rect 22376 7148 22428 7200
rect 22836 7148 22888 7200
rect 23020 7191 23072 7200
rect 23020 7157 23029 7191
rect 23029 7157 23063 7191
rect 23063 7157 23072 7191
rect 23020 7148 23072 7157
rect 3749 7046 3801 7098
rect 3813 7046 3865 7098
rect 3877 7046 3929 7098
rect 3941 7046 3993 7098
rect 4005 7046 4057 7098
rect 9347 7046 9399 7098
rect 9411 7046 9463 7098
rect 9475 7046 9527 7098
rect 9539 7046 9591 7098
rect 9603 7046 9655 7098
rect 14945 7046 14997 7098
rect 15009 7046 15061 7098
rect 15073 7046 15125 7098
rect 15137 7046 15189 7098
rect 15201 7046 15253 7098
rect 20543 7046 20595 7098
rect 20607 7046 20659 7098
rect 20671 7046 20723 7098
rect 20735 7046 20787 7098
rect 20799 7046 20851 7098
rect 5632 6987 5684 6996
rect 5632 6953 5641 6987
rect 5641 6953 5675 6987
rect 5675 6953 5684 6987
rect 5632 6944 5684 6953
rect 8484 6987 8536 6996
rect 8484 6953 8493 6987
rect 8493 6953 8527 6987
rect 8527 6953 8536 6987
rect 8484 6944 8536 6953
rect 12072 6944 12124 6996
rect 11796 6876 11848 6928
rect 12624 6944 12676 6996
rect 13912 6944 13964 6996
rect 14648 6944 14700 6996
rect 16212 6944 16264 6996
rect 18696 6944 18748 6996
rect 19248 6944 19300 6996
rect 22376 6944 22428 6996
rect 23112 6944 23164 6996
rect 1584 6740 1636 6792
rect 6184 6740 6236 6792
rect 6276 6672 6328 6724
rect 8392 6740 8444 6792
rect 9956 6740 10008 6792
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 17592 6740 17644 6792
rect 18328 6808 18380 6860
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 20536 6876 20588 6928
rect 20720 6808 20772 6860
rect 21088 6808 21140 6860
rect 9864 6672 9916 6724
rect 11152 6672 11204 6724
rect 12072 6672 12124 6724
rect 3608 6604 3660 6656
rect 9772 6604 9824 6656
rect 10232 6604 10284 6656
rect 13268 6604 13320 6656
rect 15200 6672 15252 6724
rect 16028 6672 16080 6724
rect 16948 6672 17000 6724
rect 14188 6604 14240 6656
rect 14740 6604 14792 6656
rect 15844 6604 15896 6656
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 17500 6604 17552 6656
rect 18604 6715 18656 6724
rect 18604 6681 18613 6715
rect 18613 6681 18647 6715
rect 18647 6681 18656 6715
rect 18604 6672 18656 6681
rect 19156 6740 19208 6792
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 19800 6740 19852 6792
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 21640 6851 21692 6860
rect 21640 6817 21652 6851
rect 21652 6817 21686 6851
rect 21686 6817 21692 6851
rect 21640 6808 21692 6817
rect 22284 6808 22336 6860
rect 23388 6808 23440 6860
rect 22560 6740 22612 6792
rect 19340 6672 19392 6724
rect 19616 6672 19668 6724
rect 20168 6672 20220 6724
rect 20812 6672 20864 6724
rect 18328 6604 18380 6656
rect 19156 6604 19208 6656
rect 20628 6604 20680 6656
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 21548 6604 21600 6656
rect 22652 6604 22704 6656
rect 6548 6502 6600 6554
rect 6612 6502 6664 6554
rect 6676 6502 6728 6554
rect 6740 6502 6792 6554
rect 6804 6502 6856 6554
rect 12146 6502 12198 6554
rect 12210 6502 12262 6554
rect 12274 6502 12326 6554
rect 12338 6502 12390 6554
rect 12402 6502 12454 6554
rect 17744 6502 17796 6554
rect 17808 6502 17860 6554
rect 17872 6502 17924 6554
rect 17936 6502 17988 6554
rect 18000 6502 18052 6554
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 9864 6400 9916 6452
rect 11244 6400 11296 6452
rect 5908 6332 5960 6384
rect 2136 6264 2188 6316
rect 8760 6332 8812 6384
rect 9772 6375 9824 6384
rect 9772 6341 9781 6375
rect 9781 6341 9815 6375
rect 9815 6341 9824 6375
rect 9772 6332 9824 6341
rect 10876 6332 10928 6384
rect 8944 6196 8996 6248
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 8024 6103 8076 6112
rect 8024 6069 8033 6103
rect 8033 6069 8067 6103
rect 8067 6069 8076 6103
rect 8024 6060 8076 6069
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9220 6060 9272 6112
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 11336 6264 11388 6316
rect 13176 6332 13228 6384
rect 13268 6375 13320 6384
rect 13268 6341 13286 6375
rect 13286 6341 13320 6375
rect 13268 6332 13320 6341
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 12532 6196 12584 6248
rect 13912 6443 13964 6452
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 16580 6400 16632 6452
rect 18144 6400 18196 6452
rect 18696 6400 18748 6452
rect 14280 6332 14332 6384
rect 14648 6264 14700 6316
rect 14280 6196 14332 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 16672 6332 16724 6384
rect 17132 6332 17184 6384
rect 20720 6400 20772 6452
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 21180 6400 21232 6452
rect 23020 6400 23072 6452
rect 14832 6264 14884 6316
rect 14556 6196 14608 6205
rect 11520 6128 11572 6180
rect 11980 6128 12032 6180
rect 15384 6128 15436 6180
rect 11888 6060 11940 6112
rect 12900 6060 12952 6112
rect 13544 6060 13596 6112
rect 14096 6060 14148 6112
rect 15476 6060 15528 6112
rect 17592 6264 17644 6316
rect 18696 6264 18748 6316
rect 20536 6332 20588 6384
rect 22192 6375 22244 6384
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 18512 6196 18564 6248
rect 19248 6264 19300 6316
rect 17132 6060 17184 6112
rect 22192 6341 22201 6375
rect 22201 6341 22235 6375
rect 22235 6341 22244 6375
rect 22192 6332 22244 6341
rect 22284 6375 22336 6384
rect 22284 6341 22293 6375
rect 22293 6341 22327 6375
rect 22327 6341 22336 6375
rect 22284 6332 22336 6341
rect 23480 6332 23532 6384
rect 21364 6239 21416 6248
rect 18788 6060 18840 6112
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 19984 6060 20036 6112
rect 20168 6060 20220 6112
rect 21364 6205 21373 6239
rect 21373 6205 21407 6239
rect 21407 6205 21416 6239
rect 21364 6196 21416 6205
rect 23296 6264 23348 6316
rect 21824 6196 21876 6248
rect 21732 6128 21784 6180
rect 22376 6239 22428 6248
rect 22376 6205 22385 6239
rect 22385 6205 22419 6239
rect 22419 6205 22428 6239
rect 22376 6196 22428 6205
rect 22836 6128 22888 6180
rect 23112 6128 23164 6180
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 3749 5958 3801 6010
rect 3813 5958 3865 6010
rect 3877 5958 3929 6010
rect 3941 5958 3993 6010
rect 4005 5958 4057 6010
rect 9347 5958 9399 6010
rect 9411 5958 9463 6010
rect 9475 5958 9527 6010
rect 9539 5958 9591 6010
rect 9603 5958 9655 6010
rect 14945 5958 14997 6010
rect 15009 5958 15061 6010
rect 15073 5958 15125 6010
rect 15137 5958 15189 6010
rect 15201 5958 15253 6010
rect 20543 5958 20595 6010
rect 20607 5958 20659 6010
rect 20671 5958 20723 6010
rect 20735 5958 20787 6010
rect 20799 5958 20851 6010
rect 5356 5763 5408 5772
rect 5356 5729 5365 5763
rect 5365 5729 5399 5763
rect 5399 5729 5408 5763
rect 5356 5720 5408 5729
rect 8392 5856 8444 5908
rect 8668 5856 8720 5908
rect 11704 5856 11756 5908
rect 7012 5788 7064 5840
rect 5724 5652 5776 5704
rect 5816 5652 5868 5704
rect 6552 5652 6604 5704
rect 5632 5584 5684 5636
rect 9128 5720 9180 5772
rect 9220 5720 9272 5772
rect 9588 5720 9640 5772
rect 10784 5788 10836 5840
rect 11428 5831 11480 5840
rect 11428 5797 11437 5831
rect 11437 5797 11471 5831
rect 11471 5797 11480 5831
rect 11428 5788 11480 5797
rect 12624 5856 12676 5908
rect 14556 5856 14608 5908
rect 16948 5856 17000 5908
rect 13176 5720 13228 5772
rect 13544 5720 13596 5772
rect 14096 5763 14148 5772
rect 14096 5729 14105 5763
rect 14105 5729 14139 5763
rect 14139 5729 14148 5763
rect 14096 5720 14148 5729
rect 14556 5761 14608 5772
rect 14556 5727 14568 5761
rect 14568 5727 14602 5761
rect 14602 5727 14608 5761
rect 14556 5720 14608 5727
rect 14740 5720 14792 5772
rect 17224 5788 17276 5840
rect 19064 5831 19116 5840
rect 19064 5797 19073 5831
rect 19073 5797 19107 5831
rect 19107 5797 19116 5831
rect 19064 5788 19116 5797
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 17500 5720 17552 5772
rect 19984 5856 20036 5908
rect 20904 5856 20956 5908
rect 21732 5856 21784 5908
rect 22100 5856 22152 5908
rect 23020 5899 23072 5908
rect 23020 5865 23029 5899
rect 23029 5865 23063 5899
rect 23063 5865 23072 5899
rect 23020 5856 23072 5865
rect 20444 5788 20496 5840
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 9036 5652 9088 5704
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 11704 5652 11756 5704
rect 16580 5652 16632 5704
rect 17132 5652 17184 5704
rect 17592 5652 17644 5704
rect 18604 5652 18656 5704
rect 6920 5516 6972 5568
rect 7104 5516 7156 5568
rect 16212 5584 16264 5636
rect 20076 5695 20128 5704
rect 20076 5661 20085 5695
rect 20085 5661 20119 5695
rect 20119 5661 20128 5695
rect 20076 5652 20128 5661
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 14372 5516 14424 5568
rect 16304 5559 16356 5568
rect 16304 5525 16313 5559
rect 16313 5525 16347 5559
rect 16347 5525 16356 5559
rect 16304 5516 16356 5525
rect 16856 5516 16908 5568
rect 20168 5584 20220 5636
rect 19156 5516 19208 5568
rect 20076 5516 20128 5568
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 21916 5720 21968 5772
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 21180 5668 21232 5720
rect 23664 5720 23716 5772
rect 22836 5695 22888 5704
rect 22836 5661 22845 5695
rect 22845 5661 22879 5695
rect 22879 5661 22888 5695
rect 22836 5652 22888 5661
rect 21456 5516 21508 5568
rect 22560 5559 22612 5568
rect 22560 5525 22569 5559
rect 22569 5525 22603 5559
rect 22603 5525 22612 5559
rect 22560 5516 22612 5525
rect 6548 5414 6600 5466
rect 6612 5414 6664 5466
rect 6676 5414 6728 5466
rect 6740 5414 6792 5466
rect 6804 5414 6856 5466
rect 12146 5414 12198 5466
rect 12210 5414 12262 5466
rect 12274 5414 12326 5466
rect 12338 5414 12390 5466
rect 12402 5414 12454 5466
rect 17744 5414 17796 5466
rect 17808 5414 17860 5466
rect 17872 5414 17924 5466
rect 17936 5414 17988 5466
rect 18000 5414 18052 5466
rect 5816 5355 5868 5364
rect 5816 5321 5825 5355
rect 5825 5321 5859 5355
rect 5859 5321 5868 5355
rect 5816 5312 5868 5321
rect 8024 5312 8076 5364
rect 5908 5244 5960 5296
rect 6920 5244 6972 5296
rect 7012 5176 7064 5228
rect 8484 5176 8536 5228
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7840 5108 7892 5160
rect 8392 5108 8444 5160
rect 9588 5312 9640 5364
rect 8944 5176 8996 5228
rect 11060 5312 11112 5364
rect 13544 5355 13596 5364
rect 13544 5321 13553 5355
rect 13553 5321 13587 5355
rect 13587 5321 13596 5355
rect 13544 5312 13596 5321
rect 16212 5312 16264 5364
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 17500 5355 17552 5364
rect 17500 5321 17509 5355
rect 17509 5321 17543 5355
rect 17543 5321 17552 5355
rect 17500 5312 17552 5321
rect 19156 5312 19208 5364
rect 10876 5244 10928 5296
rect 14372 5287 14424 5296
rect 14372 5253 14381 5287
rect 14381 5253 14415 5287
rect 14415 5253 14424 5287
rect 14372 5244 14424 5253
rect 16396 5244 16448 5296
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 16028 5176 16080 5228
rect 17316 5176 17368 5228
rect 10140 5108 10192 5160
rect 10784 5108 10836 5160
rect 14832 5108 14884 5160
rect 15384 5108 15436 5160
rect 15936 5108 15988 5160
rect 18788 5244 18840 5296
rect 20076 5312 20128 5364
rect 20260 5312 20312 5364
rect 20996 5355 21048 5364
rect 20996 5321 21005 5355
rect 21005 5321 21039 5355
rect 21039 5321 21048 5355
rect 20996 5312 21048 5321
rect 21364 5312 21416 5364
rect 22284 5355 22336 5364
rect 22284 5321 22293 5355
rect 22293 5321 22327 5355
rect 22327 5321 22336 5355
rect 22284 5312 22336 5321
rect 22652 5312 22704 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 20536 5287 20588 5296
rect 20536 5253 20545 5287
rect 20545 5253 20579 5287
rect 20579 5253 20588 5287
rect 20536 5244 20588 5253
rect 22192 5244 22244 5296
rect 19984 5176 20036 5228
rect 21548 5219 21600 5228
rect 21548 5185 21557 5219
rect 21557 5185 21591 5219
rect 21591 5185 21600 5219
rect 21548 5176 21600 5185
rect 20168 5108 20220 5160
rect 22560 5176 22612 5228
rect 10048 5040 10100 5092
rect 14372 5040 14424 5092
rect 7472 4972 7524 5024
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 7840 4972 7892 5024
rect 10692 4972 10744 5024
rect 16120 4972 16172 5024
rect 18696 5015 18748 5024
rect 18696 4981 18705 5015
rect 18705 4981 18739 5015
rect 18739 4981 18748 5015
rect 18696 4972 18748 4981
rect 19708 4972 19760 5024
rect 20444 4972 20496 5024
rect 3749 4870 3801 4922
rect 3813 4870 3865 4922
rect 3877 4870 3929 4922
rect 3941 4870 3993 4922
rect 4005 4870 4057 4922
rect 9347 4870 9399 4922
rect 9411 4870 9463 4922
rect 9475 4870 9527 4922
rect 9539 4870 9591 4922
rect 9603 4870 9655 4922
rect 14945 4870 14997 4922
rect 15009 4870 15061 4922
rect 15073 4870 15125 4922
rect 15137 4870 15189 4922
rect 15201 4870 15253 4922
rect 20543 4870 20595 4922
rect 20607 4870 20659 4922
rect 20671 4870 20723 4922
rect 20735 4870 20787 4922
rect 20799 4870 20851 4922
rect 6920 4768 6972 4820
rect 7472 4700 7524 4752
rect 8392 4743 8444 4752
rect 7656 4632 7708 4684
rect 8392 4709 8401 4743
rect 8401 4709 8435 4743
rect 8435 4709 8444 4743
rect 8392 4700 8444 4709
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 17592 4768 17644 4820
rect 19984 4768 20036 4820
rect 21640 4768 21692 4820
rect 10416 4632 10468 4684
rect 15476 4632 15528 4684
rect 16304 4675 16356 4684
rect 7748 4564 7800 4616
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 16304 4641 16313 4675
rect 16313 4641 16347 4675
rect 16347 4641 16356 4675
rect 16304 4632 16356 4641
rect 18236 4632 18288 4684
rect 18880 4675 18932 4684
rect 18880 4641 18889 4675
rect 18889 4641 18923 4675
rect 18923 4641 18932 4675
rect 18880 4632 18932 4641
rect 17408 4564 17460 4616
rect 18696 4564 18748 4616
rect 20076 4564 20128 4616
rect 20812 4564 20864 4616
rect 21180 4607 21232 4616
rect 21180 4573 21189 4607
rect 21189 4573 21223 4607
rect 21223 4573 21232 4607
rect 21180 4564 21232 4573
rect 21824 4632 21876 4684
rect 23296 4700 23348 4752
rect 22100 4632 22152 4684
rect 22652 4675 22704 4684
rect 22284 4564 22336 4616
rect 22652 4641 22661 4675
rect 22661 4641 22695 4675
rect 22695 4641 22704 4675
rect 22652 4632 22704 4641
rect 23388 4564 23440 4616
rect 18236 4496 18288 4548
rect 19340 4496 19392 4548
rect 20168 4496 20220 4548
rect 20260 4496 20312 4548
rect 20536 4496 20588 4548
rect 10876 4428 10928 4480
rect 16212 4428 16264 4480
rect 16580 4428 16632 4480
rect 18696 4471 18748 4480
rect 18696 4437 18705 4471
rect 18705 4437 18739 4471
rect 18739 4437 18748 4471
rect 18696 4428 18748 4437
rect 18972 4428 19024 4480
rect 19708 4428 19760 4480
rect 19800 4428 19852 4480
rect 22100 4471 22152 4480
rect 22100 4437 22109 4471
rect 22109 4437 22143 4471
rect 22143 4437 22152 4471
rect 22100 4428 22152 4437
rect 6548 4326 6600 4378
rect 6612 4326 6664 4378
rect 6676 4326 6728 4378
rect 6740 4326 6792 4378
rect 6804 4326 6856 4378
rect 12146 4326 12198 4378
rect 12210 4326 12262 4378
rect 12274 4326 12326 4378
rect 12338 4326 12390 4378
rect 12402 4326 12454 4378
rect 17744 4326 17796 4378
rect 17808 4326 17860 4378
rect 17872 4326 17924 4378
rect 17936 4326 17988 4378
rect 18000 4326 18052 4378
rect 6920 4224 6972 4276
rect 15936 4224 15988 4276
rect 18696 4224 18748 4276
rect 19800 4267 19852 4276
rect 19800 4233 19809 4267
rect 19809 4233 19843 4267
rect 19843 4233 19852 4267
rect 19800 4224 19852 4233
rect 20444 4224 20496 4276
rect 22100 4267 22152 4276
rect 22100 4233 22109 4267
rect 22109 4233 22143 4267
rect 22143 4233 22152 4267
rect 22100 4224 22152 4233
rect 14832 4156 14884 4208
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 16028 4156 16080 4208
rect 17316 4156 17368 4208
rect 16304 4088 16356 4140
rect 15660 4020 15712 4072
rect 16396 4020 16448 4072
rect 16120 3952 16172 4004
rect 16304 3952 16356 4004
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 12532 3884 12584 3936
rect 15844 3884 15896 3936
rect 16488 3884 16540 3936
rect 16672 4020 16724 4072
rect 16948 4131 17000 4140
rect 16948 4097 16957 4131
rect 16957 4097 16991 4131
rect 16991 4097 17000 4131
rect 16948 4088 17000 4097
rect 17224 4088 17276 4140
rect 20536 4088 20588 4140
rect 21272 4131 21324 4140
rect 17040 4020 17092 4072
rect 18420 4063 18472 4072
rect 18420 4029 18429 4063
rect 18429 4029 18463 4063
rect 18463 4029 18472 4063
rect 18420 4020 18472 4029
rect 19524 4063 19576 4072
rect 19524 4029 19533 4063
rect 19533 4029 19567 4063
rect 19567 4029 19576 4063
rect 19524 4020 19576 4029
rect 20444 4020 20496 4072
rect 21272 4097 21281 4131
rect 21281 4097 21315 4131
rect 21315 4097 21324 4131
rect 21272 4088 21324 4097
rect 21364 4131 21416 4140
rect 21364 4097 21373 4131
rect 21373 4097 21407 4131
rect 21407 4097 21416 4131
rect 21364 4088 21416 4097
rect 22100 4088 22152 4140
rect 23572 4088 23624 4140
rect 22744 4020 22796 4072
rect 21364 3952 21416 4004
rect 23756 4020 23808 4072
rect 23204 3952 23256 4004
rect 18052 3884 18104 3936
rect 19984 3884 20036 3936
rect 20260 3927 20312 3936
rect 20260 3893 20269 3927
rect 20269 3893 20303 3927
rect 20303 3893 20312 3927
rect 21548 3927 21600 3936
rect 20260 3884 20312 3893
rect 21548 3893 21557 3927
rect 21557 3893 21591 3927
rect 21591 3893 21600 3927
rect 21548 3884 21600 3893
rect 22468 3884 22520 3936
rect 22652 3927 22704 3936
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 3749 3782 3801 3834
rect 3813 3782 3865 3834
rect 3877 3782 3929 3834
rect 3941 3782 3993 3834
rect 4005 3782 4057 3834
rect 9347 3782 9399 3834
rect 9411 3782 9463 3834
rect 9475 3782 9527 3834
rect 9539 3782 9591 3834
rect 9603 3782 9655 3834
rect 14945 3782 14997 3834
rect 15009 3782 15061 3834
rect 15073 3782 15125 3834
rect 15137 3782 15189 3834
rect 15201 3782 15253 3834
rect 20543 3782 20595 3834
rect 20607 3782 20659 3834
rect 20671 3782 20723 3834
rect 20735 3782 20787 3834
rect 20799 3782 20851 3834
rect 9772 3680 9824 3732
rect 17224 3723 17276 3732
rect 12900 3612 12952 3664
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 19340 3723 19392 3732
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 20076 3680 20128 3732
rect 12532 3587 12584 3596
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 14372 3544 14424 3596
rect 15936 3544 15988 3596
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 16488 3544 16540 3596
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 18144 3544 18196 3596
rect 19156 3544 19208 3596
rect 5080 3476 5132 3528
rect 10600 3476 10652 3528
rect 15476 3476 15528 3528
rect 16028 3476 16080 3528
rect 18328 3476 18380 3528
rect 19340 3476 19392 3528
rect 20260 3612 20312 3664
rect 21364 3680 21416 3732
rect 22376 3680 22428 3732
rect 23020 3723 23072 3732
rect 23020 3689 23029 3723
rect 23029 3689 23063 3723
rect 23063 3689 23072 3723
rect 23020 3680 23072 3689
rect 19708 3544 19760 3596
rect 21088 3544 21140 3596
rect 22284 3587 22336 3596
rect 22284 3553 22293 3587
rect 22293 3553 22327 3587
rect 22327 3553 22336 3587
rect 22284 3544 22336 3553
rect 20168 3476 20220 3528
rect 20904 3476 20956 3528
rect 22836 3612 22888 3664
rect 22744 3519 22796 3528
rect 22744 3485 22753 3519
rect 22753 3485 22787 3519
rect 22787 3485 22796 3519
rect 22744 3476 22796 3485
rect 21088 3408 21140 3460
rect 22284 3408 22336 3460
rect 22468 3408 22520 3460
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 16212 3340 16264 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 18512 3383 18564 3392
rect 17316 3340 17368 3349
rect 18512 3349 18521 3383
rect 18521 3349 18555 3383
rect 18555 3349 18564 3383
rect 18512 3340 18564 3349
rect 19156 3340 19208 3392
rect 20444 3340 20496 3392
rect 21272 3340 21324 3392
rect 22560 3340 22612 3392
rect 6548 3238 6600 3290
rect 6612 3238 6664 3290
rect 6676 3238 6728 3290
rect 6740 3238 6792 3290
rect 6804 3238 6856 3290
rect 12146 3238 12198 3290
rect 12210 3238 12262 3290
rect 12274 3238 12326 3290
rect 12338 3238 12390 3290
rect 12402 3238 12454 3290
rect 17744 3238 17796 3290
rect 17808 3238 17860 3290
rect 17872 3238 17924 3290
rect 17936 3238 17988 3290
rect 18000 3238 18052 3290
rect 12992 3136 13044 3188
rect 17316 3136 17368 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 5080 3068 5132 3120
rect 4528 2796 4580 2848
rect 11060 3000 11112 3052
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 20352 3136 20404 3188
rect 20444 3136 20496 3188
rect 23112 3136 23164 3188
rect 19432 3068 19484 3120
rect 19800 3111 19852 3120
rect 19800 3077 19809 3111
rect 19809 3077 19843 3111
rect 19843 3077 19852 3111
rect 19800 3068 19852 3077
rect 19524 3000 19576 3052
rect 19984 3000 20036 3052
rect 20904 3000 20956 3052
rect 21180 3000 21232 3052
rect 22652 3043 22704 3052
rect 19340 2932 19392 2984
rect 20168 2932 20220 2984
rect 16396 2864 16448 2916
rect 19432 2864 19484 2916
rect 19524 2907 19576 2916
rect 19524 2873 19533 2907
rect 19533 2873 19567 2907
rect 19567 2873 19576 2907
rect 19524 2864 19576 2873
rect 19892 2864 19944 2916
rect 20536 2864 20588 2916
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 22744 3000 22796 3052
rect 22192 2932 22244 2984
rect 10600 2796 10652 2848
rect 14188 2796 14240 2848
rect 19340 2796 19392 2848
rect 19984 2796 20036 2848
rect 20352 2796 20404 2848
rect 21088 2839 21140 2848
rect 21088 2805 21097 2839
rect 21097 2805 21131 2839
rect 21131 2805 21140 2839
rect 21088 2796 21140 2805
rect 3749 2694 3801 2746
rect 3813 2694 3865 2746
rect 3877 2694 3929 2746
rect 3941 2694 3993 2746
rect 4005 2694 4057 2746
rect 9347 2694 9399 2746
rect 9411 2694 9463 2746
rect 9475 2694 9527 2746
rect 9539 2694 9591 2746
rect 9603 2694 9655 2746
rect 14945 2694 14997 2746
rect 15009 2694 15061 2746
rect 15073 2694 15125 2746
rect 15137 2694 15189 2746
rect 15201 2694 15253 2746
rect 20543 2694 20595 2746
rect 20607 2694 20659 2746
rect 20671 2694 20723 2746
rect 20735 2694 20787 2746
rect 20799 2694 20851 2746
rect 19340 2635 19392 2644
rect 19340 2601 19349 2635
rect 19349 2601 19383 2635
rect 19383 2601 19392 2635
rect 19340 2592 19392 2601
rect 19984 2592 20036 2644
rect 20168 2635 20220 2644
rect 20168 2601 20177 2635
rect 20177 2601 20211 2635
rect 20211 2601 20220 2635
rect 20168 2592 20220 2601
rect 19248 2524 19300 2576
rect 20444 2592 20496 2644
rect 22652 2592 22704 2644
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 19524 2499 19576 2508
rect 19524 2465 19533 2499
rect 19533 2465 19567 2499
rect 19567 2465 19576 2499
rect 19524 2456 19576 2465
rect 22100 2499 22152 2508
rect 22100 2465 22109 2499
rect 22109 2465 22143 2499
rect 22143 2465 22152 2499
rect 22468 2524 22520 2576
rect 23848 2524 23900 2576
rect 22100 2456 22152 2465
rect 22744 2456 22796 2508
rect 4528 2388 4580 2440
rect 6184 2388 6236 2440
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 19800 2388 19852 2440
rect 20904 2388 20956 2440
rect 22008 2388 22060 2440
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 22468 2431 22520 2440
rect 22468 2397 22477 2431
rect 22477 2397 22511 2431
rect 22511 2397 22520 2431
rect 22468 2388 22520 2397
rect 2136 2252 2188 2304
rect 10232 2252 10284 2304
rect 15476 2252 15528 2304
rect 20352 2320 20404 2372
rect 22192 2252 22244 2304
rect 22376 2295 22428 2304
rect 22376 2261 22385 2295
rect 22385 2261 22419 2295
rect 22419 2261 22428 2295
rect 22376 2252 22428 2261
rect 22652 2295 22704 2304
rect 22652 2261 22661 2295
rect 22661 2261 22695 2295
rect 22695 2261 22704 2295
rect 22652 2252 22704 2261
rect 6548 2150 6600 2202
rect 6612 2150 6664 2202
rect 6676 2150 6728 2202
rect 6740 2150 6792 2202
rect 6804 2150 6856 2202
rect 12146 2150 12198 2202
rect 12210 2150 12262 2202
rect 12274 2150 12326 2202
rect 12338 2150 12390 2202
rect 12402 2150 12454 2202
rect 17744 2150 17796 2202
rect 17808 2150 17860 2202
rect 17872 2150 17924 2202
rect 17936 2150 17988 2202
rect 18000 2150 18052 2202
<< metal2 >>
rect 294 23800 350 24600
rect 938 23800 994 24600
rect 1582 23800 1638 24600
rect 2226 23800 2282 24600
rect 2870 23800 2926 24600
rect 3514 23800 3570 24600
rect 4158 23800 4214 24600
rect 4802 23800 4858 24600
rect 5446 23800 5502 24600
rect 6090 23800 6146 24600
rect 6734 23800 6790 24600
rect 7378 23800 7434 24600
rect 8022 23800 8078 24600
rect 8666 23800 8722 24600
rect 9310 23800 9366 24600
rect 9954 23800 10010 24600
rect 10598 23800 10654 24600
rect 11242 23800 11298 24600
rect 11886 23800 11942 24600
rect 12530 23800 12586 24600
rect 13174 23800 13230 24600
rect 13818 23800 13874 24600
rect 14462 23800 14518 24600
rect 14568 23854 15056 23882
rect 308 21690 336 23800
rect 296 21684 348 21690
rect 296 21626 348 21632
rect 952 21418 980 23800
rect 1596 21894 1624 23800
rect 2240 21894 2268 23800
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2332 21729 2360 22034
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 2318 21720 2374 21729
rect 2318 21655 2374 21664
rect 2332 21554 2360 21655
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 940 21412 992 21418
rect 940 21354 992 21360
rect 2044 20936 2096 20942
rect 2042 20904 2044 20913
rect 2096 20904 2098 20913
rect 2042 20839 2098 20848
rect 2332 20602 2360 21490
rect 2608 21418 2636 21966
rect 2688 21956 2740 21962
rect 2688 21898 2740 21904
rect 2700 21690 2728 21898
rect 2884 21894 2912 23800
rect 3330 22536 3386 22545
rect 3330 22471 3386 22480
rect 2962 22128 3018 22137
rect 2962 22063 3018 22072
rect 3148 22092 3200 22098
rect 2872 21888 2924 21894
rect 2778 21856 2834 21865
rect 2872 21830 2924 21836
rect 2778 21791 2834 21800
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2516 21146 2544 21286
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 2700 20913 2728 21490
rect 2792 21146 2820 21791
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 2780 21140 2832 21146
rect 2780 21082 2832 21088
rect 2686 20904 2742 20913
rect 2686 20839 2742 20848
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 2792 18329 2820 20742
rect 2884 20602 2912 21422
rect 2976 20874 3004 22063
rect 3148 22034 3200 22040
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3068 21729 3096 21966
rect 3054 21720 3110 21729
rect 3054 21655 3110 21664
rect 3160 21622 3188 22034
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3252 21690 3280 21966
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3148 21616 3200 21622
rect 3148 21558 3200 21564
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3068 20942 3096 21490
rect 3252 21146 3280 21490
rect 3344 21332 3372 22471
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3528 21842 3556 23800
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 3608 22704 3660 22710
rect 3608 22646 3660 22652
rect 3620 22094 3648 22646
rect 4080 22386 4108 22714
rect 4080 22358 4120 22386
rect 3749 22332 4057 22341
rect 3749 22330 3755 22332
rect 3811 22330 3835 22332
rect 3891 22330 3915 22332
rect 3971 22330 3995 22332
rect 4051 22330 4057 22332
rect 3811 22278 3813 22330
rect 3993 22278 3995 22330
rect 3749 22276 3755 22278
rect 3811 22276 3835 22278
rect 3891 22276 3915 22278
rect 3971 22276 3995 22278
rect 4051 22276 4057 22278
rect 3749 22267 4057 22276
rect 4092 22250 4120 22358
rect 4080 22222 4120 22250
rect 3790 22128 3846 22137
rect 3620 22066 3740 22094
rect 3608 22024 3660 22030
rect 3606 21992 3608 22001
rect 3660 21992 3662 22001
rect 3606 21927 3662 21936
rect 3608 21888 3660 21894
rect 3528 21836 3608 21842
rect 3528 21830 3660 21836
rect 3436 21457 3464 21830
rect 3528 21814 3648 21830
rect 3516 21548 3568 21554
rect 3712 21536 3740 22066
rect 4080 22094 4108 22222
rect 3790 22063 3846 22072
rect 3988 22066 4108 22094
rect 3804 21554 3832 22063
rect 3988 21554 4016 22066
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 21690 4108 21966
rect 4172 21894 4200 23800
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4434 22264 4490 22273
rect 4434 22199 4490 22208
rect 4344 22024 4396 22030
rect 4344 21966 4396 21972
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4356 21570 4384 21966
rect 3516 21490 3568 21496
rect 3620 21508 3740 21536
rect 3792 21548 3844 21554
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3528 21332 3556 21490
rect 3344 21304 3556 21332
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3422 21040 3478 21049
rect 3148 21004 3200 21010
rect 3422 20975 3478 20984
rect 3148 20946 3200 20952
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 3160 20641 3188 20946
rect 3436 20942 3464 20975
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3146 20632 3202 20641
rect 2872 20596 2924 20602
rect 3146 20567 3202 20576
rect 2872 20538 2924 20544
rect 3238 20496 3294 20505
rect 3238 20431 3294 20440
rect 3332 20460 3384 20466
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 3068 19514 3096 19654
rect 3252 19514 3280 20431
rect 3332 20402 3384 20408
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2884 17746 2912 18362
rect 2976 18222 3004 18566
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 3068 17678 3096 18022
rect 3160 17882 3188 19314
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 3252 18698 3280 19178
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3344 18426 3372 20402
rect 3436 20262 3464 20742
rect 3528 20602 3556 21304
rect 3620 21026 3648 21508
rect 3976 21548 4028 21554
rect 3792 21490 3844 21496
rect 3896 21508 3976 21536
rect 3896 21350 3924 21508
rect 3976 21490 4028 21496
rect 4080 21542 4384 21570
rect 4080 21350 4108 21542
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 3749 21244 4057 21253
rect 3749 21242 3755 21244
rect 3811 21242 3835 21244
rect 3891 21242 3915 21244
rect 3971 21242 3995 21244
rect 4051 21242 4057 21244
rect 3811 21190 3813 21242
rect 3993 21190 3995 21242
rect 3749 21188 3755 21190
rect 3811 21188 3835 21190
rect 3891 21188 3915 21190
rect 3971 21188 3995 21190
rect 4051 21188 4057 21190
rect 3749 21179 4057 21188
rect 3792 21072 3844 21078
rect 3620 20998 3740 21026
rect 3792 21014 3844 21020
rect 3712 20942 3740 20998
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3620 20788 3648 20878
rect 3804 20788 3832 21014
rect 3620 20760 3832 20788
rect 4172 20618 4200 21422
rect 4448 21418 4476 22199
rect 4632 22030 4660 22510
rect 4816 22094 4844 23800
rect 5460 22778 5488 23800
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 4816 22066 4936 22094
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4526 21856 4582 21865
rect 4526 21791 4582 21800
rect 4540 21554 4568 21791
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4436 21412 4488 21418
rect 4436 21354 4488 21360
rect 4252 21344 4304 21350
rect 4252 21286 4304 21292
rect 4344 21344 4396 21350
rect 4540 21321 4568 21490
rect 4344 21286 4396 21292
rect 4526 21312 4582 21321
rect 4264 20913 4292 21286
rect 4356 20942 4384 21286
rect 4526 21247 4582 21256
rect 4344 20936 4396 20942
rect 4250 20904 4306 20913
rect 4344 20878 4396 20884
rect 4250 20839 4306 20848
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3804 20590 4200 20618
rect 3804 20398 3832 20590
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3436 19310 3464 20198
rect 3620 19854 3648 20198
rect 3749 20156 4057 20165
rect 3749 20154 3755 20156
rect 3811 20154 3835 20156
rect 3891 20154 3915 20156
rect 3971 20154 3995 20156
rect 4051 20154 4057 20156
rect 3811 20102 3813 20154
rect 3993 20102 3995 20154
rect 3749 20100 3755 20102
rect 3811 20100 3835 20102
rect 3891 20100 3915 20102
rect 3971 20100 3995 20102
rect 4051 20100 4057 20102
rect 3749 20091 4057 20100
rect 4172 20058 4200 20402
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 3608 19848 3660 19854
rect 3608 19790 3660 19796
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3528 19174 3556 19654
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3528 18970 3556 19110
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3620 18902 3648 19314
rect 4080 19122 4108 19314
rect 4080 19094 4200 19122
rect 3749 19068 4057 19077
rect 3749 19066 3755 19068
rect 3811 19066 3835 19068
rect 3891 19066 3915 19068
rect 3971 19066 3995 19068
rect 4051 19066 4057 19068
rect 3811 19014 3813 19066
rect 3993 19014 3995 19066
rect 3749 19012 3755 19014
rect 3811 19012 3835 19014
rect 3891 19012 3915 19014
rect 3971 19012 3995 19014
rect 4051 19012 4057 19014
rect 3749 19003 4057 19012
rect 4172 18970 4200 19094
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 3608 18896 3660 18902
rect 3608 18838 3660 18844
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3436 18465 3464 18770
rect 3514 18728 3570 18737
rect 3514 18663 3570 18672
rect 3528 18630 3556 18663
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3882 18592 3938 18601
rect 3882 18527 3938 18536
rect 3422 18456 3478 18465
rect 3332 18420 3384 18426
rect 3422 18391 3478 18400
rect 3332 18362 3384 18368
rect 3436 18290 3464 18391
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1492 15360 1544 15366
rect 1490 15328 1492 15337
rect 1544 15328 1546 15337
rect 1490 15263 1546 15272
rect 1688 14074 1716 15438
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9217 1440 9522
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1596 6798 1624 9318
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 2148 6322 2176 13806
rect 3252 12986 3280 18226
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3436 17746 3464 18090
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3436 13530 3464 17682
rect 3528 15978 3556 18294
rect 3896 18222 3924 18527
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4172 18057 4200 18158
rect 4158 18048 4214 18057
rect 3749 17980 4057 17989
rect 4158 17983 4214 17992
rect 3749 17978 3755 17980
rect 3811 17978 3835 17980
rect 3891 17978 3915 17980
rect 3971 17978 3995 17980
rect 4051 17978 4057 17980
rect 3811 17926 3813 17978
rect 3993 17926 3995 17978
rect 3749 17924 3755 17926
rect 3811 17924 3835 17926
rect 3891 17924 3915 17926
rect 3971 17924 3995 17926
rect 4051 17924 4057 17926
rect 3749 17915 4057 17924
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 4066 17640 4122 17649
rect 3620 16250 3648 17614
rect 4066 17575 4122 17584
rect 4080 17542 4108 17575
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 3749 16892 4057 16901
rect 3749 16890 3755 16892
rect 3811 16890 3835 16892
rect 3891 16890 3915 16892
rect 3971 16890 3995 16892
rect 4051 16890 4057 16892
rect 3811 16838 3813 16890
rect 3993 16838 3995 16890
rect 3749 16836 3755 16838
rect 3811 16836 3835 16838
rect 3891 16836 3915 16838
rect 3971 16836 3995 16838
rect 4051 16836 4057 16838
rect 3749 16827 4057 16836
rect 4172 16794 4200 17002
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3749 15804 4057 15813
rect 3749 15802 3755 15804
rect 3811 15802 3835 15804
rect 3891 15802 3915 15804
rect 3971 15802 3995 15804
rect 4051 15802 4057 15804
rect 3811 15750 3813 15802
rect 3993 15750 3995 15802
rect 3749 15748 3755 15750
rect 3811 15748 3835 15750
rect 3891 15748 3915 15750
rect 3971 15748 3995 15750
rect 4051 15748 4057 15750
rect 3749 15739 4057 15748
rect 4264 15337 4292 20742
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4356 20058 4384 20538
rect 4632 20534 4660 21966
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 21622 4752 21830
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 4816 21418 4844 21966
rect 4908 21894 4936 22066
rect 4896 21888 4948 21894
rect 4896 21830 4948 21836
rect 5000 21554 5028 22578
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5448 22432 5500 22438
rect 5354 22400 5410 22409
rect 5448 22374 5500 22380
rect 5354 22335 5410 22344
rect 5368 22234 5396 22335
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5172 22160 5224 22166
rect 5172 22102 5224 22108
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5184 22030 5212 22102
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4804 21412 4856 21418
rect 4804 21354 4856 21360
rect 4908 20924 4936 21422
rect 5172 21412 5224 21418
rect 5172 21354 5224 21360
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 5000 20942 5028 21286
rect 4816 20896 4936 20924
rect 4988 20936 5040 20942
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4448 20262 4476 20334
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4356 19514 4384 19790
rect 4632 19514 4660 20334
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4356 16046 4384 19246
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4356 15570 4384 15982
rect 4448 15706 4476 19314
rect 4540 17202 4568 19314
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4632 17338 4660 18158
rect 4724 18034 4752 20742
rect 4816 20641 4844 20896
rect 4988 20878 5040 20884
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4802 20632 4858 20641
rect 4802 20567 4858 20576
rect 4804 20324 4856 20330
rect 4804 20266 4856 20272
rect 4816 19310 4844 20266
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4816 18426 4844 18906
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4724 18006 4844 18034
rect 4816 17762 4844 18006
rect 4724 17734 4844 17762
rect 4724 17610 4752 17734
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4816 17134 4844 17546
rect 4908 17354 4936 20742
rect 5000 20641 5028 20878
rect 4986 20632 5042 20641
rect 4986 20567 5042 20576
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 4986 18184 5042 18193
rect 4986 18119 5042 18128
rect 5000 18086 5028 18119
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5092 17542 5120 19994
rect 5184 19378 5212 21354
rect 5276 21350 5304 22102
rect 5460 22030 5488 22374
rect 5448 22024 5500 22030
rect 5552 22012 5580 22442
rect 5724 22024 5776 22030
rect 5552 21984 5724 22012
rect 5448 21966 5500 21972
rect 5724 21966 5776 21972
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5460 21554 5488 21626
rect 5644 21554 5672 21830
rect 5448 21548 5500 21554
rect 5632 21548 5684 21554
rect 5500 21508 5580 21536
rect 5448 21490 5500 21496
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5368 20942 5396 21354
rect 5552 21350 5580 21508
rect 5632 21490 5684 21496
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5368 19786 5396 19926
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5184 18601 5212 18702
rect 5170 18592 5226 18601
rect 5170 18527 5226 18536
rect 5276 18465 5304 19654
rect 5368 19514 5396 19722
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5460 18873 5488 21286
rect 5736 21146 5764 21966
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 6012 21418 6040 21830
rect 6104 21486 6132 23800
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 6196 22030 6224 22714
rect 6748 22574 6776 23800
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 7208 22273 7236 22510
rect 7194 22264 7250 22273
rect 7194 22199 7250 22208
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6368 22024 6420 22030
rect 6736 22024 6788 22030
rect 6368 21966 6420 21972
rect 6550 21992 6606 22001
rect 6184 21888 6236 21894
rect 6182 21856 6184 21865
rect 6236 21856 6238 21865
rect 6182 21791 6238 21800
rect 6196 21604 6224 21791
rect 6380 21729 6408 21966
rect 6734 21992 6736 22001
rect 6788 21992 6790 22001
rect 6606 21950 6684 21978
rect 6550 21927 6606 21936
rect 6656 21894 6684 21950
rect 6734 21927 6790 21936
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 7010 21856 7066 21865
rect 6366 21720 6422 21729
rect 6366 21655 6422 21664
rect 6196 21576 6316 21604
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 6090 21176 6146 21185
rect 5724 21140 5776 21146
rect 6090 21111 6146 21120
rect 5724 21082 5776 21088
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5724 21004 5776 21010
rect 5724 20946 5776 20952
rect 5446 18864 5502 18873
rect 5446 18799 5502 18808
rect 5552 18680 5580 20946
rect 5736 20618 5764 20946
rect 5908 20800 5960 20806
rect 6104 20777 6132 21111
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 5908 20742 5960 20748
rect 6090 20768 6146 20777
rect 5644 20602 5764 20618
rect 5632 20596 5764 20602
rect 5684 20590 5764 20596
rect 5632 20538 5684 20544
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 5816 20528 5868 20534
rect 5816 20470 5868 20476
rect 5736 19961 5764 20470
rect 5828 20262 5856 20470
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5722 19952 5778 19961
rect 5722 19887 5778 19896
rect 5828 19854 5856 20198
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5630 18864 5686 18873
rect 5630 18799 5686 18808
rect 5543 18652 5580 18680
rect 5356 18624 5408 18630
rect 5543 18612 5571 18652
rect 5543 18584 5580 18612
rect 5356 18566 5408 18572
rect 5262 18456 5318 18465
rect 5262 18391 5318 18400
rect 5276 18222 5304 18391
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5368 18154 5396 18566
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5170 18048 5226 18057
rect 5170 17983 5226 17992
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 4908 17326 5028 17354
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4724 16658 4752 16934
rect 4816 16794 4844 17070
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4540 16182 4568 16390
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4250 15328 4306 15337
rect 4250 15263 4306 15272
rect 3749 14716 4057 14725
rect 3749 14714 3755 14716
rect 3811 14714 3835 14716
rect 3891 14714 3915 14716
rect 3971 14714 3995 14716
rect 4051 14714 4057 14716
rect 3811 14662 3813 14714
rect 3993 14662 3995 14714
rect 3749 14660 3755 14662
rect 3811 14660 3835 14662
rect 3891 14660 3915 14662
rect 3971 14660 3995 14662
rect 4051 14660 4057 14662
rect 3749 14651 4057 14660
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 3749 13628 4057 13637
rect 3749 13626 3755 13628
rect 3811 13626 3835 13628
rect 3891 13626 3915 13628
rect 3971 13626 3995 13628
rect 4051 13626 4057 13628
rect 3811 13574 3813 13626
rect 3993 13574 3995 13626
rect 3749 13572 3755 13574
rect 3811 13572 3835 13574
rect 3891 13572 3915 13574
rect 3971 13572 3995 13574
rect 4051 13572 4057 13574
rect 3749 13563 4057 13572
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 4172 12986 4200 13670
rect 4356 13530 4384 13874
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4158 12880 4214 12889
rect 3332 12844 3384 12850
rect 4158 12815 4214 12824
rect 3332 12786 3384 12792
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11762 3188 12038
rect 3344 11898 3372 12786
rect 3749 12540 4057 12549
rect 3749 12538 3755 12540
rect 3811 12538 3835 12540
rect 3891 12538 3915 12540
rect 3971 12538 3995 12540
rect 4051 12538 4057 12540
rect 3811 12486 3813 12538
rect 3993 12486 3995 12538
rect 3749 12484 3755 12486
rect 3811 12484 3835 12486
rect 3891 12484 3915 12486
rect 3971 12484 3995 12486
rect 4051 12484 4057 12486
rect 3749 12475 4057 12484
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 4172 11830 4200 12815
rect 4264 11898 4292 13126
rect 4356 12782 4384 13330
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4448 12986 4476 13262
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4540 11898 4568 16118
rect 4632 15978 4660 16390
rect 4816 16182 4844 16730
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4160 11824 4212 11830
rect 3882 11792 3938 11801
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3608 11756 3660 11762
rect 4160 11766 4212 11772
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 3882 11727 3938 11736
rect 4252 11756 4304 11762
rect 3608 11698 3660 11704
rect 3620 10266 3648 11698
rect 3896 11694 3924 11727
rect 4252 11698 4304 11704
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 3749 11452 4057 11461
rect 3749 11450 3755 11452
rect 3811 11450 3835 11452
rect 3891 11450 3915 11452
rect 3971 11450 3995 11452
rect 4051 11450 4057 11452
rect 3811 11398 3813 11450
rect 3993 11398 3995 11450
rect 3749 11396 3755 11398
rect 3811 11396 3835 11398
rect 3891 11396 3915 11398
rect 3971 11396 3995 11398
rect 4051 11396 4057 11398
rect 3749 11387 4057 11396
rect 3749 10364 4057 10373
rect 3749 10362 3755 10364
rect 3811 10362 3835 10364
rect 3891 10362 3915 10364
rect 3971 10362 3995 10364
rect 4051 10362 4057 10364
rect 3811 10310 3813 10362
rect 3993 10310 3995 10362
rect 3749 10308 3755 10310
rect 3811 10308 3835 10310
rect 3891 10308 3915 10310
rect 3971 10308 3995 10310
rect 4051 10308 4057 10310
rect 3749 10299 4057 10308
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 4172 10130 4200 11630
rect 4264 10538 4292 11698
rect 4356 11218 4384 11766
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4356 11098 4384 11154
rect 4356 11070 4476 11098
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10810 4384 10950
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4448 10146 4476 11070
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4540 10674 4568 10950
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4632 10266 4660 15914
rect 4816 15706 4844 16118
rect 4908 15978 4936 17206
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4894 15056 4950 15065
rect 4894 14991 4896 15000
rect 4948 14991 4950 15000
rect 4896 14962 4948 14968
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4724 11218 4752 14758
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4908 12918 4936 14214
rect 5000 13394 5028 17326
rect 5184 16726 5212 17983
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 5368 15434 5396 18090
rect 5552 17270 5580 18584
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 16114 5580 16934
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5080 15156 5132 15162
rect 5644 15144 5672 18799
rect 5736 18766 5764 19654
rect 5828 19446 5856 19790
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5828 18834 5856 19382
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5920 18034 5948 20742
rect 6090 20703 6146 20712
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6012 20058 6040 20402
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6104 19922 6132 20198
rect 6196 20058 6224 20946
rect 6288 20806 6316 21576
rect 6472 21536 6500 21830
rect 6548 21788 6856 21797
rect 7010 21791 7066 21800
rect 6548 21786 6554 21788
rect 6610 21786 6634 21788
rect 6690 21786 6714 21788
rect 6770 21786 6794 21788
rect 6850 21786 6856 21788
rect 6610 21734 6612 21786
rect 6792 21734 6794 21786
rect 6548 21732 6554 21734
rect 6610 21732 6634 21734
rect 6690 21732 6714 21734
rect 6770 21732 6794 21734
rect 6850 21732 6856 21734
rect 6548 21723 6856 21732
rect 6380 21508 6500 21536
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6274 20632 6330 20641
rect 6274 20567 6330 20576
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 19786 6132 19858
rect 6092 19780 6144 19786
rect 6092 19722 6144 19728
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6104 18737 6132 19314
rect 6288 18850 6316 20567
rect 6380 18970 6408 21508
rect 7024 21434 7052 21791
rect 7102 21720 7158 21729
rect 7102 21655 7158 21664
rect 6460 21412 6512 21418
rect 6460 21354 6512 21360
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6840 21406 7052 21434
rect 6472 20942 6500 21354
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6552 20936 6604 20942
rect 6656 20913 6684 21354
rect 6840 21078 6868 21406
rect 7012 21344 7064 21350
rect 7116 21321 7144 21655
rect 7012 21286 7064 21292
rect 7102 21312 7158 21321
rect 6828 21072 6880 21078
rect 6828 21014 6880 21020
rect 7024 21010 7052 21286
rect 7102 21247 7158 21256
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6828 20936 6880 20942
rect 6552 20878 6604 20884
rect 6642 20904 6698 20913
rect 6564 20806 6592 20878
rect 6642 20839 6698 20848
rect 6826 20904 6828 20913
rect 6880 20904 6882 20913
rect 6826 20839 6882 20848
rect 7208 20806 7236 22199
rect 7392 22094 7420 23800
rect 8036 22438 8064 23800
rect 8680 22506 8708 23800
rect 9324 22778 9352 23800
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 8668 22500 8720 22506
rect 8668 22442 8720 22448
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8758 22400 8814 22409
rect 8758 22335 8814 22344
rect 8772 22098 8800 22335
rect 9347 22332 9655 22341
rect 9347 22330 9353 22332
rect 9409 22330 9433 22332
rect 9489 22330 9513 22332
rect 9569 22330 9593 22332
rect 9649 22330 9655 22332
rect 9409 22278 9411 22330
rect 9591 22278 9593 22330
rect 9347 22276 9353 22278
rect 9409 22276 9433 22278
rect 9489 22276 9513 22278
rect 9569 22276 9593 22278
rect 9649 22276 9655 22278
rect 9347 22267 9655 22276
rect 9036 22160 9088 22166
rect 9036 22102 9088 22108
rect 7300 22066 7420 22094
rect 8760 22092 8812 22098
rect 7300 21486 7328 22066
rect 8760 22034 8812 22040
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 7392 21554 7420 21898
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 8116 21888 8168 21894
rect 8576 21888 8628 21894
rect 8116 21830 8168 21836
rect 8574 21856 8576 21865
rect 8628 21856 8630 21865
rect 7576 21690 7604 21830
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 7392 21146 7420 21490
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 6548 20700 6856 20709
rect 6548 20698 6554 20700
rect 6610 20698 6634 20700
rect 6690 20698 6714 20700
rect 6770 20698 6794 20700
rect 6850 20698 6856 20700
rect 6610 20646 6612 20698
rect 6792 20646 6794 20698
rect 6548 20644 6554 20646
rect 6610 20644 6634 20646
rect 6690 20644 6714 20646
rect 6770 20644 6794 20646
rect 6850 20644 6856 20646
rect 6548 20635 6856 20644
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6748 20398 6776 20538
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6548 19612 6856 19621
rect 6548 19610 6554 19612
rect 6610 19610 6634 19612
rect 6690 19610 6714 19612
rect 6770 19610 6794 19612
rect 6850 19610 6856 19612
rect 6610 19558 6612 19610
rect 6792 19558 6794 19610
rect 6548 19556 6554 19558
rect 6610 19556 6634 19558
rect 6690 19556 6714 19558
rect 6770 19556 6794 19558
rect 6850 19556 6856 19558
rect 6548 19547 6856 19556
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6288 18822 6408 18850
rect 6090 18728 6146 18737
rect 6146 18686 6316 18714
rect 6090 18663 6146 18672
rect 6000 18624 6052 18630
rect 6104 18603 6132 18663
rect 6000 18566 6052 18572
rect 5828 18006 5948 18034
rect 5724 17604 5776 17610
rect 5828 17592 5856 18006
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 5776 17564 5856 17592
rect 5724 17546 5776 17552
rect 5920 16114 5948 17818
rect 6012 17610 6040 18566
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6104 17678 6132 18022
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 6196 17270 6224 18158
rect 6288 17882 6316 18686
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6288 16590 6316 17274
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 6288 15638 6316 16526
rect 6380 15978 6408 18822
rect 6548 18524 6856 18533
rect 6548 18522 6554 18524
rect 6610 18522 6634 18524
rect 6690 18522 6714 18524
rect 6770 18522 6794 18524
rect 6850 18522 6856 18524
rect 6610 18470 6612 18522
rect 6792 18470 6794 18522
rect 6548 18468 6554 18470
rect 6610 18468 6634 18470
rect 6690 18468 6714 18470
rect 6770 18468 6794 18470
rect 6850 18468 6856 18470
rect 6548 18459 6856 18468
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6472 18057 6500 18226
rect 6458 18048 6514 18057
rect 6458 17983 6514 17992
rect 6932 17785 6960 20742
rect 7300 20369 7328 20810
rect 7286 20360 7342 20369
rect 7286 20295 7342 20304
rect 7576 19786 7604 21422
rect 7944 21146 7972 21830
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 6918 17776 6974 17785
rect 6918 17711 6974 17720
rect 6548 17436 6856 17445
rect 6548 17434 6554 17436
rect 6610 17434 6634 17436
rect 6690 17434 6714 17436
rect 6770 17434 6794 17436
rect 6850 17434 6856 17436
rect 6610 17382 6612 17434
rect 6792 17382 6794 17434
rect 6548 17380 6554 17382
rect 6610 17380 6634 17382
rect 6690 17380 6714 17382
rect 6770 17380 6794 17382
rect 6850 17380 6856 17382
rect 6548 17371 6856 17380
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6564 16794 6592 16934
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6840 16522 6868 17070
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6828 16516 6880 16522
rect 6828 16458 6880 16464
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6472 15706 6500 16458
rect 6548 16348 6856 16357
rect 6548 16346 6554 16348
rect 6610 16346 6634 16348
rect 6690 16346 6714 16348
rect 6770 16346 6794 16348
rect 6850 16346 6856 16348
rect 6610 16294 6612 16346
rect 6792 16294 6794 16346
rect 6548 16292 6554 16294
rect 6610 16292 6634 16294
rect 6690 16292 6714 16294
rect 6770 16292 6794 16294
rect 6850 16292 6856 16294
rect 6548 16283 6856 16292
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6548 15260 6856 15269
rect 6548 15258 6554 15260
rect 6610 15258 6634 15260
rect 6690 15258 6714 15260
rect 6770 15258 6794 15260
rect 6850 15258 6856 15260
rect 6610 15206 6612 15258
rect 6792 15206 6794 15258
rect 6548 15204 6554 15206
rect 6610 15204 6634 15206
rect 6690 15204 6714 15206
rect 6770 15204 6794 15206
rect 6850 15204 6856 15206
rect 6548 15195 6856 15204
rect 5080 15098 5132 15104
rect 5552 15116 5672 15144
rect 5092 14482 5120 15098
rect 5552 14958 5580 15116
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5644 14618 5672 14962
rect 5632 14612 5684 14618
rect 5552 14572 5632 14600
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 14006 5120 14214
rect 5080 14000 5132 14006
rect 5080 13942 5132 13948
rect 5552 13870 5580 14572
rect 5632 14554 5684 14560
rect 5736 13870 5764 15030
rect 6932 15026 6960 16118
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5828 14278 5856 14554
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5920 13870 5948 14894
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5184 12986 5212 13670
rect 5276 13326 5304 13670
rect 5354 13424 5410 13433
rect 6288 13394 6316 14962
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 5354 13359 5356 13368
rect 5408 13359 5410 13368
rect 6276 13388 6328 13394
rect 5356 13330 5408 13336
rect 6276 13330 6328 13336
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 5368 12782 5396 13330
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12986 5856 13126
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 6380 12782 6408 14758
rect 6656 14346 6684 14758
rect 6932 14414 6960 14962
rect 7024 14618 7052 18634
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18358 7144 18566
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7194 18320 7250 18329
rect 7194 18255 7250 18264
rect 7208 17610 7236 18255
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7300 17066 7328 19722
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7392 18426 7420 18702
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7470 17640 7526 17649
rect 7470 17575 7526 17584
rect 7484 17542 7512 17575
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7392 15094 7420 17478
rect 7668 15910 7696 20742
rect 8036 20482 8064 21490
rect 8128 21486 8156 21830
rect 8574 21791 8630 21800
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8128 21350 8156 21422
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8128 21010 8156 21286
rect 8220 21010 8248 21490
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8116 20800 8168 20806
rect 8220 20788 8248 20946
rect 8168 20760 8248 20788
rect 8116 20742 8168 20748
rect 8680 20602 8708 21898
rect 8758 21856 8814 21865
rect 8758 21791 8814 21800
rect 8772 21185 8800 21791
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8758 21176 8814 21185
rect 8758 21111 8814 21120
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8864 20942 8892 21082
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8036 20454 8524 20482
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18630 7788 19110
rect 8312 18698 8340 20334
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8404 19378 8432 19994
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8496 19174 8524 20454
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7760 17202 7788 18566
rect 8312 18154 8340 18634
rect 8496 18426 8524 19110
rect 8588 18834 8616 20402
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8680 18193 8708 20334
rect 8760 19780 8812 19786
rect 8760 19722 8812 19728
rect 8772 18970 8800 19722
rect 8864 19718 8892 20878
rect 8956 20330 8984 21422
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 9048 19530 9076 22102
rect 9968 22094 9996 23800
rect 10230 22264 10286 22273
rect 10230 22199 10286 22208
rect 10244 22098 10272 22199
rect 9876 22066 9996 22094
rect 10232 22092 10284 22098
rect 9128 22024 9180 22030
rect 9876 22001 9904 22066
rect 10232 22034 10284 22040
rect 9128 21966 9180 21972
rect 9862 21992 9918 22001
rect 9140 21457 9168 21966
rect 9862 21927 9918 21936
rect 10046 21992 10102 22001
rect 10046 21927 10102 21936
rect 10140 21956 10192 21962
rect 10060 21894 10088 21927
rect 10140 21898 10192 21904
rect 9312 21888 9364 21894
rect 10048 21888 10100 21894
rect 9312 21830 9364 21836
rect 9402 21856 9458 21865
rect 9324 21690 9352 21830
rect 10048 21830 10100 21836
rect 9402 21791 9458 21800
rect 9416 21690 9444 21791
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9404 21684 9456 21690
rect 9456 21644 9628 21672
rect 9404 21626 9456 21632
rect 9496 21480 9548 21486
rect 9126 21448 9182 21457
rect 9416 21440 9496 21468
rect 9416 21434 9444 21440
rect 9126 21383 9182 21392
rect 9232 21406 9444 21434
rect 9496 21422 9548 21428
rect 9600 21434 9628 21644
rect 10060 21593 10088 21830
rect 10046 21584 10102 21593
rect 10046 21519 10102 21528
rect 9864 21480 9916 21486
rect 9600 21406 9812 21434
rect 10152 21468 10180 21898
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 9916 21440 10180 21468
rect 9864 21422 9916 21428
rect 9126 21176 9182 21185
rect 9232 21146 9260 21406
rect 9680 21344 9732 21350
rect 9784 21321 9812 21406
rect 9680 21286 9732 21292
rect 9770 21312 9826 21321
rect 9347 21244 9655 21253
rect 9347 21242 9353 21244
rect 9409 21242 9433 21244
rect 9489 21242 9513 21244
rect 9569 21242 9593 21244
rect 9649 21242 9655 21244
rect 9409 21190 9411 21242
rect 9591 21190 9593 21242
rect 9347 21188 9353 21190
rect 9409 21188 9433 21190
rect 9489 21188 9513 21190
rect 9569 21188 9593 21190
rect 9649 21188 9655 21190
rect 9347 21179 9655 21188
rect 9126 21111 9182 21120
rect 9220 21140 9272 21146
rect 8864 19502 9076 19530
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8666 18184 8722 18193
rect 8300 18148 8352 18154
rect 8666 18119 8722 18128
rect 8300 18090 8352 18096
rect 8864 18086 8892 19502
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 8036 16794 8064 17274
rect 8024 16788 8076 16794
rect 8076 16748 8248 16776
rect 8024 16730 8076 16736
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8128 16114 8156 16390
rect 8220 16114 8248 16748
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 8128 15570 8156 16050
rect 8864 16046 8892 18022
rect 9048 17338 9076 18294
rect 9140 17762 9168 21111
rect 9220 21082 9272 21088
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9508 20942 9536 21082
rect 9692 21010 9720 21286
rect 9770 21247 9826 21256
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9772 20936 9824 20942
rect 10152 20913 10180 21440
rect 9772 20878 9824 20884
rect 10138 20904 10194 20913
rect 9508 20602 9536 20878
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9784 20534 9812 20878
rect 10138 20839 10194 20848
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9220 20324 9272 20330
rect 9220 20266 9272 20272
rect 9232 19786 9260 20266
rect 9347 20156 9655 20165
rect 9347 20154 9353 20156
rect 9409 20154 9433 20156
rect 9489 20154 9513 20156
rect 9569 20154 9593 20156
rect 9649 20154 9655 20156
rect 9409 20102 9411 20154
rect 9591 20102 9593 20154
rect 9347 20100 9353 20102
rect 9409 20100 9433 20102
rect 9489 20100 9513 20102
rect 9569 20100 9593 20102
rect 9649 20100 9655 20102
rect 9347 20091 9655 20100
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9692 19514 9720 20334
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9588 19372 9640 19378
rect 9640 19332 9720 19360
rect 9588 19314 9640 19320
rect 9347 19068 9655 19077
rect 9347 19066 9353 19068
rect 9409 19066 9433 19068
rect 9489 19066 9513 19068
rect 9569 19066 9593 19068
rect 9649 19066 9655 19068
rect 9409 19014 9411 19066
rect 9591 19014 9593 19066
rect 9347 19012 9353 19014
rect 9409 19012 9433 19014
rect 9489 19012 9513 19014
rect 9569 19012 9593 19014
rect 9649 19012 9655 19014
rect 9347 19003 9655 19012
rect 9692 18766 9720 19332
rect 9876 18766 9904 19450
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9692 18306 9720 18702
rect 9692 18290 9812 18306
rect 9692 18284 9824 18290
rect 9692 18278 9772 18284
rect 9772 18226 9824 18232
rect 9347 17980 9655 17989
rect 9347 17978 9353 17980
rect 9409 17978 9433 17980
rect 9489 17978 9513 17980
rect 9569 17978 9593 17980
rect 9649 17978 9655 17980
rect 9409 17926 9411 17978
rect 9591 17926 9593 17978
rect 9347 17924 9353 17926
rect 9409 17924 9433 17926
rect 9489 17924 9513 17926
rect 9569 17924 9593 17926
rect 9649 17924 9655 17926
rect 9347 17915 9655 17924
rect 9140 17734 9260 17762
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 8956 16658 8984 17206
rect 9048 17134 9076 17274
rect 9140 17202 9168 17614
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8956 16538 8984 16594
rect 9232 16538 9260 17734
rect 9347 16892 9655 16901
rect 9347 16890 9353 16892
rect 9409 16890 9433 16892
rect 9489 16890 9513 16892
rect 9569 16890 9593 16892
rect 9649 16890 9655 16892
rect 9409 16838 9411 16890
rect 9591 16838 9593 16890
rect 9347 16836 9353 16838
rect 9409 16836 9433 16838
rect 9489 16836 9513 16838
rect 9569 16836 9593 16838
rect 9649 16836 9655 16838
rect 9347 16827 9655 16836
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 8956 16510 9076 16538
rect 9048 16046 9076 16510
rect 9140 16510 9260 16538
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6472 14074 6500 14214
rect 6548 14172 6856 14181
rect 6548 14170 6554 14172
rect 6610 14170 6634 14172
rect 6690 14170 6714 14172
rect 6770 14170 6794 14172
rect 6850 14170 6856 14172
rect 6610 14118 6612 14170
rect 6792 14118 6794 14170
rect 6548 14116 6554 14118
rect 6610 14116 6634 14118
rect 6690 14116 6714 14118
rect 6770 14116 6794 14118
rect 6850 14116 6856 14118
rect 6548 14107 6856 14116
rect 6932 14074 6960 14350
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6932 13530 6960 13874
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7024 13258 7052 13670
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6548 13084 6856 13093
rect 6548 13082 6554 13084
rect 6610 13082 6634 13084
rect 6690 13082 6714 13084
rect 6770 13082 6794 13084
rect 6850 13082 6856 13084
rect 6610 13030 6612 13082
rect 6792 13030 6794 13082
rect 6548 13028 6554 13030
rect 6610 13028 6634 13030
rect 6690 13028 6714 13030
rect 6770 13028 6794 13030
rect 6850 13028 6856 13030
rect 6548 13019 6856 13028
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 11898 4936 12582
rect 5000 12434 5028 12718
rect 5000 12406 5120 12434
rect 5092 12306 5120 12406
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 6000 12300 6052 12306
rect 6104 12288 6132 12718
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 6380 12442 6408 12582
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6052 12260 6132 12288
rect 6000 12242 6052 12248
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11898 5028 12038
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5092 11694 5120 12242
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5460 11898 5488 12106
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 6104 11694 6132 12260
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 6472 11898 6500 12106
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6548 11996 6856 12005
rect 6548 11994 6554 11996
rect 6610 11994 6634 11996
rect 6690 11994 6714 11996
rect 6770 11994 6794 11996
rect 6850 11994 6856 11996
rect 6610 11942 6612 11994
rect 6792 11942 6794 11994
rect 6548 11940 6554 11942
rect 6610 11940 6634 11942
rect 6690 11940 6714 11942
rect 6770 11940 6794 11942
rect 6850 11940 6856 11942
rect 6548 11931 6856 11940
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10606 4752 11154
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5000 10810 5028 10950
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 5092 10538 5120 11086
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 10810 5488 11018
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4160 10124 4212 10130
rect 4448 10118 4660 10146
rect 4160 10066 4212 10072
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9042 3188 9318
rect 3344 9110 3372 9522
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 7546 3280 8774
rect 3436 8362 3464 9998
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 9722 3556 9862
rect 3804 9722 3832 9930
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3620 9178 3648 9522
rect 4448 9518 4476 9930
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4436 9512 4488 9518
rect 4356 9460 4436 9466
rect 4356 9454 4488 9460
rect 4356 9438 4476 9454
rect 3749 9276 4057 9285
rect 3749 9274 3755 9276
rect 3811 9274 3835 9276
rect 3891 9274 3915 9276
rect 3971 9274 3995 9276
rect 4051 9274 4057 9276
rect 3811 9222 3813 9274
rect 3993 9222 3995 9274
rect 3749 9220 3755 9222
rect 3811 9220 3835 9222
rect 3891 9220 3915 9222
rect 3971 9220 3995 9222
rect 4051 9220 4057 9222
rect 3749 9211 4057 9220
rect 4356 9178 4384 9438
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4172 8974 4200 9046
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3620 6662 3648 8434
rect 3712 8362 3740 8570
rect 4172 8430 4200 8910
rect 3884 8424 3936 8430
rect 4160 8424 4212 8430
rect 3936 8372 4108 8378
rect 3884 8366 4108 8372
rect 4160 8366 4212 8372
rect 3700 8356 3752 8362
rect 3896 8350 4108 8366
rect 3700 8298 3752 8304
rect 4080 8242 4108 8350
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 8242 4292 8298
rect 4356 8294 4384 9114
rect 4448 9042 4476 9318
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4540 8906 4568 9522
rect 4632 9042 4660 10118
rect 5092 10062 5120 10474
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 5092 8974 5120 9862
rect 5368 9518 5396 10066
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5368 9042 5396 9114
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5736 8906 5764 11222
rect 7024 11082 7052 12038
rect 7208 11354 7236 12106
rect 7392 11830 7420 12582
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 10130 5948 10406
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6196 9586 6224 9930
rect 6472 9926 6500 11018
rect 6548 10908 6856 10917
rect 6548 10906 6554 10908
rect 6610 10906 6634 10908
rect 6690 10906 6714 10908
rect 6770 10906 6794 10908
rect 6850 10906 6856 10908
rect 6610 10854 6612 10906
rect 6792 10854 6794 10906
rect 6548 10852 6554 10854
rect 6610 10852 6634 10854
rect 6690 10852 6714 10854
rect 6770 10852 6794 10854
rect 6850 10852 6856 10854
rect 6548 10843 6856 10852
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6840 10577 6868 10678
rect 6826 10568 6882 10577
rect 6826 10503 6828 10512
rect 6880 10503 6882 10512
rect 6828 10474 6880 10480
rect 7116 10470 7144 11086
rect 7760 11014 7788 15370
rect 8128 14618 8156 15506
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15162 8248 15438
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 9048 14958 9076 15982
rect 9140 15706 9168 16510
rect 9692 16454 9720 16730
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9232 15366 9260 16390
rect 9347 15804 9655 15813
rect 9347 15802 9353 15804
rect 9409 15802 9433 15804
rect 9489 15802 9513 15804
rect 9569 15802 9593 15804
rect 9649 15802 9655 15804
rect 9409 15750 9411 15802
rect 9591 15750 9593 15802
rect 9347 15748 9353 15750
rect 9409 15748 9433 15750
rect 9489 15748 9513 15750
rect 9569 15748 9593 15750
rect 9649 15748 9655 15750
rect 9347 15739 9655 15748
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9324 15178 9352 15370
rect 9232 15150 9352 15178
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8128 13938 8156 14554
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 8036 13326 8064 13670
rect 8128 13530 8156 13874
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8220 13258 8248 14758
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8312 13258 8340 13466
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8404 12646 8432 13874
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12442 8432 12582
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8956 12238 8984 14214
rect 9232 13734 9260 15150
rect 9347 14716 9655 14725
rect 9347 14714 9353 14716
rect 9409 14714 9433 14716
rect 9489 14714 9513 14716
rect 9569 14714 9593 14716
rect 9649 14714 9655 14716
rect 9409 14662 9411 14714
rect 9591 14662 9593 14714
rect 9347 14660 9353 14662
rect 9409 14660 9433 14662
rect 9489 14660 9513 14662
rect 9569 14660 9593 14662
rect 9649 14660 9655 14662
rect 9347 14651 9655 14660
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9692 14074 9720 14486
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9784 14006 9812 14282
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9048 12918 9076 13194
rect 9232 13190 9260 13670
rect 9347 13628 9655 13637
rect 9347 13626 9353 13628
rect 9409 13626 9433 13628
rect 9489 13626 9513 13628
rect 9569 13626 9593 13628
rect 9649 13626 9655 13628
rect 9409 13574 9411 13626
rect 9591 13574 9593 13626
rect 9347 13572 9353 13574
rect 9409 13572 9433 13574
rect 9489 13572 9513 13574
rect 9569 13572 9593 13574
rect 9649 13572 9655 13574
rect 9347 13563 9655 13572
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12986 9444 13126
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9416 12850 9444 12922
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9347 12540 9655 12549
rect 9347 12538 9353 12540
rect 9409 12538 9433 12540
rect 9489 12538 9513 12540
rect 9569 12538 9593 12540
rect 9649 12538 9655 12540
rect 9409 12486 9411 12538
rect 9591 12486 9593 12538
rect 9347 12484 9353 12486
rect 9409 12484 9433 12486
rect 9489 12484 9513 12486
rect 9569 12484 9593 12486
rect 9649 12484 9655 12486
rect 9347 12475 9655 12484
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 8036 11558 8064 12106
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11150 8064 11494
rect 9347 11452 9655 11461
rect 9347 11450 9353 11452
rect 9409 11450 9433 11452
rect 9489 11450 9513 11452
rect 9569 11450 9593 11452
rect 9649 11450 9655 11452
rect 9409 11398 9411 11450
rect 9591 11398 9593 11450
rect 9347 11396 9353 11398
rect 9409 11396 9433 11398
rect 9489 11396 9513 11398
rect 9569 11396 9593 11398
rect 9649 11396 9655 11398
rect 9347 11387 9655 11396
rect 9692 11150 9720 11834
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 8116 10736 8168 10742
rect 8116 10678 8168 10684
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6548 9820 6856 9829
rect 6548 9818 6554 9820
rect 6610 9818 6634 9820
rect 6690 9818 6714 9820
rect 6770 9818 6794 9820
rect 6850 9818 6856 9820
rect 6610 9766 6612 9818
rect 6792 9766 6794 9818
rect 6548 9764 6554 9766
rect 6610 9764 6634 9766
rect 6690 9764 6714 9766
rect 6770 9764 6794 9766
rect 6850 9764 6856 9766
rect 6548 9755 6856 9764
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4448 8566 4476 8774
rect 4908 8634 4936 8774
rect 6196 8634 6224 9522
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 6288 9178 6316 9386
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4080 8214 4292 8242
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 3749 8188 4057 8197
rect 3749 8186 3755 8188
rect 3811 8186 3835 8188
rect 3891 8186 3915 8188
rect 3971 8186 3995 8188
rect 4051 8186 4057 8188
rect 3811 8134 3813 8186
rect 3993 8134 3995 8186
rect 3749 8132 3755 8134
rect 3811 8132 3835 8134
rect 3891 8132 3915 8134
rect 3971 8132 3995 8134
rect 4051 8132 4057 8134
rect 3749 8123 4057 8132
rect 4356 7342 4384 8230
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 3749 7100 4057 7109
rect 3749 7098 3755 7100
rect 3811 7098 3835 7100
rect 3891 7098 3915 7100
rect 3971 7098 3995 7100
rect 4051 7098 4057 7100
rect 3811 7046 3813 7098
rect 3993 7046 3995 7098
rect 3749 7044 3755 7046
rect 3811 7044 3835 7046
rect 3891 7044 3915 7046
rect 3971 7044 3995 7046
rect 4051 7044 4057 7046
rect 3749 7035 4057 7044
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 3749 6012 4057 6021
rect 3749 6010 3755 6012
rect 3811 6010 3835 6012
rect 3891 6010 3915 6012
rect 3971 6010 3995 6012
rect 4051 6010 4057 6012
rect 3811 5958 3813 6010
rect 3993 5958 3995 6010
rect 3749 5956 3755 5958
rect 3811 5956 3835 5958
rect 3891 5956 3915 5958
rect 3971 5956 3995 5958
rect 4051 5956 4057 5958
rect 3749 5947 4057 5956
rect 5368 5778 5396 7754
rect 5552 7478 5580 7822
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 7002 5672 7346
rect 5736 7290 5764 7686
rect 5816 7336 5868 7342
rect 5736 7284 5816 7290
rect 5736 7278 5868 7284
rect 5736 7262 5856 7278
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5736 5710 5764 7262
rect 5920 6390 5948 7686
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6196 6798 6224 7482
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6288 6730 6316 9114
rect 6472 8566 6500 9318
rect 6656 9110 6684 9522
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6932 8974 6960 9658
rect 7300 9654 7328 10202
rect 7944 9722 7972 10678
rect 8128 10577 8156 10678
rect 8114 10568 8170 10577
rect 8114 10503 8170 10512
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10062 8248 10406
rect 9347 10364 9655 10373
rect 9347 10362 9353 10364
rect 9409 10362 9433 10364
rect 9489 10362 9513 10364
rect 9569 10362 9593 10364
rect 9649 10362 9655 10364
rect 9409 10310 9411 10362
rect 9591 10310 9593 10362
rect 9347 10308 9353 10310
rect 9409 10308 9433 10310
rect 9489 10308 9513 10310
rect 9569 10308 9593 10310
rect 9649 10308 9655 10310
rect 9347 10299 9655 10308
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 7288 8832 7340 8838
rect 7392 8786 7420 9590
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 7340 8780 7420 8786
rect 7288 8774 7420 8780
rect 7300 8758 7420 8774
rect 6548 8732 6856 8741
rect 6548 8730 6554 8732
rect 6610 8730 6634 8732
rect 6690 8730 6714 8732
rect 6770 8730 6794 8732
rect 6850 8730 6856 8732
rect 6610 8678 6612 8730
rect 6792 8678 6794 8730
rect 6548 8676 6554 8678
rect 6610 8676 6634 8678
rect 6690 8676 6714 8678
rect 6770 8676 6794 8678
rect 6850 8676 6856 8678
rect 6548 8667 6856 8676
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6472 8294 6500 8502
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6472 7478 6500 8230
rect 6932 7818 6960 8570
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6548 7644 6856 7653
rect 6548 7642 6554 7644
rect 6610 7642 6634 7644
rect 6690 7642 6714 7644
rect 6770 7642 6794 7644
rect 6850 7642 6856 7644
rect 6610 7590 6612 7642
rect 6792 7590 6794 7642
rect 6548 7588 6554 7590
rect 6610 7588 6634 7590
rect 6690 7588 6714 7590
rect 6770 7588 6794 7590
rect 6850 7588 6856 7590
rect 6548 7579 6856 7588
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6548 6556 6856 6565
rect 6548 6554 6554 6556
rect 6610 6554 6634 6556
rect 6690 6554 6714 6556
rect 6770 6554 6794 6556
rect 6850 6554 6856 6556
rect 6610 6502 6612 6554
rect 6792 6502 6794 6554
rect 6548 6500 6554 6502
rect 6610 6500 6634 6502
rect 6690 6500 6714 6502
rect 6770 6500 6794 6502
rect 6850 6500 6856 6502
rect 6548 6491 6856 6500
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5166 5672 5578
rect 5828 5370 5856 5646
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5920 5302 5948 6326
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6564 5710 6592 6054
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6548 5468 6856 5477
rect 6548 5466 6554 5468
rect 6610 5466 6634 5468
rect 6690 5466 6714 5468
rect 6770 5466 6794 5468
rect 6850 5466 6856 5468
rect 6610 5414 6612 5466
rect 6792 5414 6794 5466
rect 6548 5412 6554 5414
rect 6610 5412 6634 5414
rect 6690 5412 6714 5414
rect 6770 5412 6794 5414
rect 6850 5412 6856 5414
rect 6548 5403 6856 5412
rect 6932 5302 6960 5510
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 7024 5234 7052 5782
rect 7116 5574 7144 8434
rect 7392 8090 7420 8758
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 3749 4924 4057 4933
rect 3749 4922 3755 4924
rect 3811 4922 3835 4924
rect 3891 4922 3915 4924
rect 3971 4922 3995 4924
rect 4051 4922 4057 4924
rect 3811 4870 3813 4922
rect 3993 4870 3995 4922
rect 3749 4868 3755 4870
rect 3811 4868 3835 4870
rect 3891 4868 3915 4870
rect 3971 4868 3995 4870
rect 4051 4868 4057 4870
rect 3749 4859 4057 4868
rect 6932 4826 6960 5102
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6548 4380 6856 4389
rect 6548 4378 6554 4380
rect 6610 4378 6634 4380
rect 6690 4378 6714 4380
rect 6770 4378 6794 4380
rect 6850 4378 6856 4380
rect 6610 4326 6612 4378
rect 6792 4326 6794 4378
rect 6548 4324 6554 4326
rect 6610 4324 6634 4326
rect 6690 4324 6714 4326
rect 6770 4324 6794 4326
rect 6850 4324 6856 4326
rect 6548 4315 6856 4324
rect 6932 4282 6960 4762
rect 7484 4758 7512 4966
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7668 4690 7696 4966
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7760 4622 7788 5510
rect 8036 5370 8064 6054
rect 8128 5710 8156 8298
rect 8496 7818 8524 8502
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8496 7002 8524 7754
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8404 6458 8432 6734
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8404 5914 8432 6394
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8496 5234 8524 6054
rect 8680 5914 8708 7686
rect 8956 7478 8984 7686
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8772 7206 8800 7346
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8772 6390 8800 7142
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8956 5234 8984 6190
rect 9048 5710 9076 9318
rect 9347 9276 9655 9285
rect 9347 9274 9353 9276
rect 9409 9274 9433 9276
rect 9489 9274 9513 9276
rect 9569 9274 9593 9276
rect 9649 9274 9655 9276
rect 9409 9222 9411 9274
rect 9591 9222 9593 9274
rect 9347 9220 9353 9222
rect 9409 9220 9433 9222
rect 9489 9220 9513 9222
rect 9569 9220 9593 9222
rect 9649 9220 9655 9222
rect 9347 9211 9655 9220
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8566 10088 8910
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9347 8188 9655 8197
rect 9347 8186 9353 8188
rect 9409 8186 9433 8188
rect 9489 8186 9513 8188
rect 9569 8186 9593 8188
rect 9649 8186 9655 8188
rect 9409 8134 9411 8186
rect 9591 8134 9593 8186
rect 9347 8132 9353 8134
rect 9409 8132 9433 8134
rect 9489 8132 9513 8134
rect 9569 8132 9593 8134
rect 9649 8132 9655 8134
rect 9347 8123 9655 8132
rect 9692 7954 9720 8434
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9347 7100 9655 7109
rect 9347 7098 9353 7100
rect 9409 7098 9433 7100
rect 9489 7098 9513 7100
rect 9569 7098 9593 7100
rect 9649 7098 9655 7100
rect 9409 7046 9411 7098
rect 9591 7046 9593 7098
rect 9347 7044 9353 7046
rect 9409 7044 9433 7046
rect 9489 7044 9513 7046
rect 9569 7044 9593 7046
rect 9649 7044 9655 7046
rect 9347 7035 9655 7044
rect 9692 6322 9720 7482
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9876 7290 9904 7414
rect 9876 7262 9996 7290
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6730 9904 7142
rect 9968 6798 9996 7262
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6390 9812 6598
rect 9876 6458 9904 6666
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5778 9168 6190
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9232 5778 9260 6054
rect 9347 6012 9655 6021
rect 9347 6010 9353 6012
rect 9409 6010 9433 6012
rect 9489 6010 9513 6012
rect 9569 6010 9593 6012
rect 9649 6010 9655 6012
rect 9409 5958 9411 6010
rect 9591 5958 9593 6010
rect 9347 5956 9353 5958
rect 9409 5956 9433 5958
rect 9489 5956 9513 5958
rect 9569 5956 9593 5958
rect 9649 5956 9655 5958
rect 9347 5947 9655 5956
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9600 5370 9628 5714
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 10152 5166 10180 20839
rect 10244 20058 10272 21626
rect 10428 21486 10456 21830
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10336 20466 10364 21422
rect 10428 20806 10456 21422
rect 10520 20942 10548 21626
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10612 20602 10640 23800
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10888 22030 10916 22442
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10704 21078 10732 21490
rect 10692 21072 10744 21078
rect 10692 21014 10744 21020
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10244 18426 10272 19994
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10244 17066 10272 17546
rect 10336 17542 10364 20402
rect 10612 19854 10640 20538
rect 10704 20448 10732 20742
rect 10784 20460 10836 20466
rect 10704 20420 10784 20448
rect 10784 20402 10836 20408
rect 10888 19854 10916 20742
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 10428 19446 10456 19654
rect 10416 19440 10468 19446
rect 10416 19382 10468 19388
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10520 17338 10548 18226
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10244 16522 10272 17002
rect 10704 16522 10732 19654
rect 10888 19446 10916 19790
rect 10980 19514 11008 22170
rect 11256 22094 11284 23800
rect 11900 22778 11928 23800
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11072 22066 11284 22094
rect 11072 21468 11100 22066
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11164 21622 11192 21966
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11072 21440 11192 21468
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11072 20398 11100 21286
rect 11164 20534 11192 21440
rect 11348 21146 11376 21830
rect 11440 21457 11468 22714
rect 12164 22704 12216 22710
rect 12164 22646 12216 22652
rect 11520 22500 11572 22506
rect 11520 22442 11572 22448
rect 11426 21448 11482 21457
rect 11426 21383 11482 21392
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 11164 19786 11192 20334
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11164 19514 11192 19722
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10888 18698 10916 19382
rect 10980 18834 11008 19450
rect 11334 19408 11390 19417
rect 11334 19343 11336 19352
rect 11388 19343 11390 19352
rect 11336 19314 11388 19320
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 11428 18692 11480 18698
rect 11428 18634 11480 18640
rect 10888 18426 10916 18634
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 11440 18154 11468 18634
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11256 17882 11284 18022
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11426 17776 11482 17785
rect 11426 17711 11482 17720
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11334 17640 11390 17649
rect 11072 17338 11100 17614
rect 11334 17575 11390 17584
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11150 16552 11206 16561
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10692 16516 10744 16522
rect 11150 16487 11206 16496
rect 10692 16458 10744 16464
rect 10704 16153 10732 16458
rect 10690 16144 10746 16153
rect 11164 16114 11192 16487
rect 11348 16114 11376 17575
rect 11440 16114 11468 17711
rect 11532 17338 11560 22442
rect 12176 22438 12204 22646
rect 12544 22506 12572 23800
rect 12532 22500 12584 22506
rect 12532 22442 12584 22448
rect 12716 22500 12768 22506
rect 12716 22442 12768 22448
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12176 22098 12204 22374
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11624 16726 11652 21490
rect 11716 21010 11744 21830
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11704 21004 11756 21010
rect 11704 20946 11756 20952
rect 11808 18970 11836 21422
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11796 18964 11848 18970
rect 11716 18924 11796 18952
rect 11716 18086 11744 18924
rect 11796 18906 11848 18912
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11900 16998 11928 20878
rect 11992 20074 12020 21830
rect 12084 21690 12112 22034
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 12146 21788 12454 21797
rect 12146 21786 12152 21788
rect 12208 21786 12232 21788
rect 12288 21786 12312 21788
rect 12368 21786 12392 21788
rect 12448 21786 12454 21788
rect 12208 21734 12210 21786
rect 12390 21734 12392 21786
rect 12146 21732 12152 21734
rect 12208 21732 12232 21734
rect 12288 21732 12312 21734
rect 12368 21732 12392 21734
rect 12448 21732 12454 21734
rect 12146 21723 12454 21732
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12084 20584 12112 21286
rect 12544 20806 12572 21558
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12146 20700 12454 20709
rect 12146 20698 12152 20700
rect 12208 20698 12232 20700
rect 12288 20698 12312 20700
rect 12368 20698 12392 20700
rect 12448 20698 12454 20700
rect 12208 20646 12210 20698
rect 12390 20646 12392 20698
rect 12146 20644 12152 20646
rect 12208 20644 12232 20646
rect 12288 20644 12312 20646
rect 12368 20644 12392 20646
rect 12448 20644 12454 20646
rect 12146 20635 12454 20644
rect 12084 20556 12296 20584
rect 12268 20398 12296 20556
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 11992 20046 12204 20074
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11980 19780 12032 19786
rect 11980 19722 12032 19728
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 10690 16079 10746 16088
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15570 10732 15846
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10796 15026 10824 15302
rect 11348 15026 11376 15438
rect 11808 15162 11836 15642
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10336 12306 10364 14350
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10888 13530 10916 13942
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10980 13258 11008 14214
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10520 12442 10548 13126
rect 11072 12986 11100 14758
rect 11348 14618 11376 14962
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 14074 11284 14214
rect 11348 14074 11376 14554
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11058 12744 11114 12753
rect 10784 12708 10836 12714
rect 11058 12679 11060 12688
rect 10784 12650 10836 12656
rect 11112 12679 11114 12688
rect 11060 12650 11112 12656
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10796 12374 10824 12650
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 11286 10364 11698
rect 10428 11354 10456 12106
rect 11348 11830 11376 12922
rect 11440 12646 11468 14282
rect 11624 12986 11652 14554
rect 11808 14278 11836 14894
rect 11900 14550 11928 14962
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11900 14006 11928 14486
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10198 10364 10950
rect 11532 10674 11560 11630
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 10520 10470 10548 10610
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 10266 10548 10406
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10520 10062 10548 10202
rect 11624 10130 11652 12378
rect 11702 12336 11758 12345
rect 11702 12271 11758 12280
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9722 10548 9998
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 8974 10640 9522
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8634 10640 8910
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10704 8498 10732 9454
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 6662 10272 7346
rect 10782 7304 10838 7313
rect 10782 7239 10838 7248
rect 10690 6896 10746 6905
rect 10690 6831 10746 6840
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 7852 5030 7880 5102
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 8404 4758 8432 5102
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9347 4924 9655 4933
rect 9347 4922 9353 4924
rect 9409 4922 9433 4924
rect 9489 4922 9513 4924
rect 9569 4922 9593 4924
rect 9649 4922 9655 4924
rect 9409 4870 9411 4922
rect 9591 4870 9593 4922
rect 9347 4868 9353 4870
rect 9409 4868 9433 4870
rect 9489 4868 9513 4870
rect 9569 4868 9593 4870
rect 9649 4868 9655 4870
rect 9347 4859 9655 4868
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 3749 3836 4057 3845
rect 3749 3834 3755 3836
rect 3811 3834 3835 3836
rect 3891 3834 3915 3836
rect 3971 3834 3995 3836
rect 4051 3834 4057 3836
rect 3811 3782 3813 3834
rect 3993 3782 3995 3834
rect 3749 3780 3755 3782
rect 3811 3780 3835 3782
rect 3891 3780 3915 3782
rect 3971 3780 3995 3782
rect 4051 3780 4057 3782
rect 3749 3771 4057 3780
rect 9347 3836 9655 3845
rect 9347 3834 9353 3836
rect 9409 3834 9433 3836
rect 9489 3834 9513 3836
rect 9569 3834 9593 3836
rect 9649 3834 9655 3836
rect 9409 3782 9411 3834
rect 9591 3782 9593 3834
rect 9347 3780 9353 3782
rect 9409 3780 9433 3782
rect 9489 3780 9513 3782
rect 9569 3780 9593 3782
rect 9649 3780 9655 3782
rect 9347 3771 9655 3780
rect 9784 3738 9812 4626
rect 10060 4622 10088 5034
rect 10704 5030 10732 6831
rect 10796 6254 10824 7239
rect 10888 6390 10916 9114
rect 11348 7954 11376 9318
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11164 6730 11192 7686
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11256 6458 11284 7686
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 11348 6322 11376 7890
rect 11440 7886 11468 8774
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11428 7540 11480 7546
rect 11532 7528 11560 8434
rect 11480 7500 11560 7528
rect 11428 7482 11480 7488
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10796 5846 10824 6190
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11532 6066 11560 6122
rect 11440 6038 11560 6066
rect 11440 5846 11468 6038
rect 11716 5914 11744 12271
rect 11808 11898 11836 12786
rect 11992 12434 12020 19722
rect 12084 19514 12112 19926
rect 12176 19922 12204 20046
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 12146 19612 12454 19621
rect 12146 19610 12152 19612
rect 12208 19610 12232 19612
rect 12288 19610 12312 19612
rect 12368 19610 12392 19612
rect 12448 19610 12454 19612
rect 12208 19558 12210 19610
rect 12390 19558 12392 19610
rect 12146 19556 12152 19558
rect 12208 19556 12232 19558
rect 12288 19556 12312 19558
rect 12368 19556 12392 19558
rect 12448 19556 12454 19558
rect 12146 19547 12454 19556
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12084 18358 12112 19450
rect 12146 18524 12454 18533
rect 12146 18522 12152 18524
rect 12208 18522 12232 18524
rect 12288 18522 12312 18524
rect 12368 18522 12392 18524
rect 12448 18522 12454 18524
rect 12208 18470 12210 18522
rect 12390 18470 12392 18522
rect 12146 18468 12152 18470
rect 12208 18468 12232 18470
rect 12288 18468 12312 18470
rect 12368 18468 12392 18470
rect 12448 18468 12454 18470
rect 12146 18459 12454 18468
rect 12636 18358 12664 21898
rect 12728 21622 12756 22442
rect 13188 22273 13216 23800
rect 13174 22264 13230 22273
rect 13174 22199 13230 22208
rect 13084 22024 13136 22030
rect 13188 22012 13216 22199
rect 13136 21984 13216 22012
rect 13268 22024 13320 22030
rect 13084 21966 13136 21972
rect 13268 21966 13320 21972
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13832 21978 13860 23800
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 13084 21888 13136 21894
rect 13280 21865 13308 21966
rect 13084 21830 13136 21836
rect 13266 21856 13322 21865
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 19961 12756 21286
rect 12912 20942 12940 21422
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12820 20058 12848 20742
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12714 19952 12770 19961
rect 12714 19887 12770 19896
rect 12808 19916 12860 19922
rect 12728 19854 12756 19887
rect 12808 19858 12860 19864
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12820 19378 12848 19858
rect 12912 19553 12940 20878
rect 12898 19544 12954 19553
rect 12898 19479 12954 19488
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12820 18970 12848 19314
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 13004 18630 13032 20946
rect 13096 20058 13124 21830
rect 13266 21791 13322 21800
rect 13372 21672 13400 21966
rect 13832 21950 13952 21978
rect 13924 21690 13952 21950
rect 13188 21644 13400 21672
rect 13912 21684 13964 21690
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13188 19854 13216 21644
rect 13912 21626 13964 21632
rect 13266 21584 13322 21593
rect 13266 21519 13322 21528
rect 13280 21486 13308 21519
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13280 20942 13308 21422
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13268 20800 13320 20806
rect 13268 20742 13320 20748
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13280 20262 13308 20742
rect 13372 20602 13400 20742
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13464 20330 13492 21422
rect 13728 21072 13780 21078
rect 13726 21040 13728 21049
rect 13820 21072 13872 21078
rect 13780 21040 13782 21049
rect 13820 21014 13872 21020
rect 13726 20975 13782 20984
rect 13634 20632 13690 20641
rect 13634 20567 13690 20576
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13266 19952 13322 19961
rect 13266 19887 13322 19896
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13096 18630 13124 19654
rect 13188 19378 13216 19654
rect 13280 19514 13308 19887
rect 13372 19854 13400 19994
rect 13556 19922 13584 20198
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13648 19514 13676 20567
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13832 19394 13860 21014
rect 13648 19378 13860 19394
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13636 19372 13860 19378
rect 13688 19366 13860 19372
rect 13912 19372 13964 19378
rect 13636 19314 13688 19320
rect 13912 19314 13964 19320
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12624 18352 12676 18358
rect 13004 18329 13032 18566
rect 13082 18456 13138 18465
rect 13082 18391 13138 18400
rect 12624 18294 12676 18300
rect 12990 18320 13046 18329
rect 12990 18255 13046 18264
rect 13096 18154 13124 18391
rect 13740 18204 13768 19246
rect 13740 18176 13860 18204
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13188 17882 13216 18090
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13726 17776 13782 17785
rect 13726 17711 13782 17720
rect 13740 17678 13768 17711
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12146 17436 12454 17445
rect 12146 17434 12152 17436
rect 12208 17434 12232 17436
rect 12288 17434 12312 17436
rect 12368 17434 12392 17436
rect 12448 17434 12454 17436
rect 12208 17382 12210 17434
rect 12390 17382 12392 17434
rect 12146 17380 12152 17382
rect 12208 17380 12232 17382
rect 12288 17380 12312 17382
rect 12368 17380 12392 17382
rect 12448 17380 12454 17382
rect 12146 17371 12454 17380
rect 12146 16348 12454 16357
rect 12146 16346 12152 16348
rect 12208 16346 12232 16348
rect 12288 16346 12312 16348
rect 12368 16346 12392 16348
rect 12448 16346 12454 16348
rect 12208 16294 12210 16346
rect 12390 16294 12392 16346
rect 12146 16292 12152 16294
rect 12208 16292 12232 16294
rect 12288 16292 12312 16294
rect 12368 16292 12392 16294
rect 12448 16292 12454 16294
rect 12146 16283 12454 16292
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 15609 12296 15846
rect 12452 15706 12480 16186
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12254 15600 12310 15609
rect 12254 15535 12310 15544
rect 12146 15260 12454 15269
rect 12146 15258 12152 15260
rect 12208 15258 12232 15260
rect 12288 15258 12312 15260
rect 12368 15258 12392 15260
rect 12448 15258 12454 15260
rect 12208 15206 12210 15258
rect 12390 15206 12392 15258
rect 12146 15204 12152 15206
rect 12208 15204 12232 15206
rect 12288 15204 12312 15206
rect 12368 15204 12392 15206
rect 12448 15204 12454 15206
rect 12146 15195 12454 15204
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14414 12480 14894
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12146 14172 12454 14181
rect 12146 14170 12152 14172
rect 12208 14170 12232 14172
rect 12288 14170 12312 14172
rect 12368 14170 12392 14172
rect 12448 14170 12454 14172
rect 12208 14118 12210 14170
rect 12390 14118 12392 14170
rect 12146 14116 12152 14118
rect 12208 14116 12232 14118
rect 12288 14116 12312 14118
rect 12368 14116 12392 14118
rect 12448 14116 12454 14118
rect 12146 14107 12454 14116
rect 12146 13084 12454 13093
rect 12146 13082 12152 13084
rect 12208 13082 12232 13084
rect 12288 13082 12312 13084
rect 12368 13082 12392 13084
rect 12448 13082 12454 13084
rect 12208 13030 12210 13082
rect 12390 13030 12392 13082
rect 12146 13028 12152 13030
rect 12208 13028 12232 13030
rect 12288 13028 12312 13030
rect 12368 13028 12392 13030
rect 12448 13028 12454 13030
rect 12146 13019 12454 13028
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12442 12204 12582
rect 11900 12406 12020 12434
rect 12164 12436 12216 12442
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 10742 11836 11494
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11808 9722 11836 10678
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11808 6934 11836 7346
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11900 6118 11928 12406
rect 12164 12378 12216 12384
rect 12176 12306 12204 12378
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12268 12170 12296 12310
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11354 12020 12038
rect 12146 11996 12454 12005
rect 12146 11994 12152 11996
rect 12208 11994 12232 11996
rect 12288 11994 12312 11996
rect 12368 11994 12392 11996
rect 12448 11994 12454 11996
rect 12208 11942 12210 11994
rect 12390 11942 12392 11994
rect 12146 11940 12152 11942
rect 12208 11940 12232 11942
rect 12288 11940 12312 11942
rect 12368 11940 12392 11942
rect 12448 11940 12454 11942
rect 12146 11931 12454 11940
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11992 11082 12020 11290
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 12084 10674 12112 11086
rect 12146 10908 12454 10917
rect 12146 10906 12152 10908
rect 12208 10906 12232 10908
rect 12288 10906 12312 10908
rect 12368 10906 12392 10908
rect 12448 10906 12454 10908
rect 12208 10854 12210 10906
rect 12390 10854 12392 10906
rect 12146 10852 12152 10854
rect 12208 10852 12232 10854
rect 12288 10852 12312 10854
rect 12368 10852 12392 10854
rect 12448 10852 12454 10854
rect 12146 10843 12454 10852
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12084 7857 12112 9862
rect 12146 9820 12454 9829
rect 12146 9818 12152 9820
rect 12208 9818 12232 9820
rect 12288 9818 12312 9820
rect 12368 9818 12392 9820
rect 12448 9818 12454 9820
rect 12208 9766 12210 9818
rect 12390 9766 12392 9818
rect 12146 9764 12152 9766
rect 12208 9764 12232 9766
rect 12288 9764 12312 9766
rect 12368 9764 12392 9766
rect 12448 9764 12454 9766
rect 12146 9755 12454 9764
rect 12146 8732 12454 8741
rect 12146 8730 12152 8732
rect 12208 8730 12232 8732
rect 12288 8730 12312 8732
rect 12368 8730 12392 8732
rect 12448 8730 12454 8732
rect 12208 8678 12210 8730
rect 12390 8678 12392 8730
rect 12146 8676 12152 8678
rect 12208 8676 12232 8678
rect 12288 8676 12312 8678
rect 12368 8676 12392 8678
rect 12448 8676 12454 8678
rect 12146 8667 12454 8676
rect 12070 7848 12126 7857
rect 12070 7783 12126 7792
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11992 6186 12020 7346
rect 12084 7002 12112 7686
rect 12146 7644 12454 7653
rect 12146 7642 12152 7644
rect 12208 7642 12232 7644
rect 12288 7642 12312 7644
rect 12368 7642 12392 7644
rect 12448 7642 12454 7644
rect 12208 7590 12210 7642
rect 12390 7590 12392 7642
rect 12146 7588 12152 7590
rect 12208 7588 12232 7590
rect 12288 7588 12312 7590
rect 12368 7588 12392 7590
rect 12448 7588 12454 7590
rect 12146 7579 12454 7588
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12084 6730 12112 6938
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12146 6556 12454 6565
rect 12146 6554 12152 6556
rect 12208 6554 12232 6556
rect 12288 6554 12312 6556
rect 12368 6554 12392 6556
rect 12448 6554 12454 6556
rect 12208 6502 12210 6554
rect 12390 6502 12392 6554
rect 12146 6500 12152 6502
rect 12208 6500 12232 6502
rect 12288 6500 12312 6502
rect 12368 6500 12392 6502
rect 12448 6500 12454 6502
rect 12146 6491 12454 6500
rect 12544 6254 12572 17546
rect 13004 17202 13032 17614
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12728 16794 12756 17138
rect 13832 17066 13860 18176
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 14822 12664 15846
rect 12820 15706 12848 16050
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13464 15162 13492 15370
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13648 15094 13676 16458
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12820 14618 12848 14758
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13280 14385 13308 14758
rect 13372 14482 13400 14758
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13266 14376 13322 14385
rect 12900 14340 12952 14346
rect 13266 14311 13322 14320
rect 13636 14340 13688 14346
rect 12900 14282 12952 14288
rect 13636 14282 13688 14288
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12918 12848 13126
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12728 12306 12756 12650
rect 12820 12442 12848 12854
rect 12808 12436 12860 12442
rect 12912 12434 12940 14282
rect 13648 14074 13676 14282
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 12912 12406 13032 12434
rect 12808 12378 12860 12384
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11762 12848 12038
rect 13004 11830 13032 12406
rect 13188 12238 13216 13262
rect 13740 12434 13768 14418
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12850 13860 13126
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13924 12442 13952 19314
rect 14016 18426 14044 22374
rect 14108 22166 14136 22374
rect 14384 22234 14412 22578
rect 14372 22228 14424 22234
rect 14372 22170 14424 22176
rect 14096 22160 14148 22166
rect 14096 22102 14148 22108
rect 14280 22160 14332 22166
rect 14280 22102 14332 22108
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14108 19922 14136 20402
rect 14200 19990 14228 20742
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14108 18306 14136 18906
rect 14200 18766 14228 19246
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14292 18465 14320 22102
rect 14476 22030 14504 23800
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14384 21010 14412 21422
rect 14372 21004 14424 21010
rect 14372 20946 14424 20952
rect 14476 20942 14504 21490
rect 14568 21078 14596 23854
rect 15028 23746 15056 23854
rect 15106 23800 15162 24600
rect 15750 23800 15806 24600
rect 16394 23800 16450 24600
rect 16776 23854 16988 23882
rect 15120 23746 15148 23800
rect 15028 23718 15148 23746
rect 14945 22332 15253 22341
rect 14945 22330 14951 22332
rect 15007 22330 15031 22332
rect 15087 22330 15111 22332
rect 15167 22330 15191 22332
rect 15247 22330 15253 22332
rect 15007 22278 15009 22330
rect 15189 22278 15191 22330
rect 14945 22276 14951 22278
rect 15007 22276 15031 22278
rect 15087 22276 15111 22278
rect 15167 22276 15191 22278
rect 15247 22276 15253 22278
rect 14945 22267 15253 22276
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 14556 21072 14608 21078
rect 14556 21014 14608 21020
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14476 20777 14504 20878
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14462 20768 14518 20777
rect 14462 20703 14518 20712
rect 14568 19417 14596 20810
rect 14554 19408 14610 19417
rect 14372 19372 14424 19378
rect 14554 19343 14610 19352
rect 14372 19314 14424 19320
rect 14278 18456 14334 18465
rect 14278 18391 14334 18400
rect 14016 18278 14136 18306
rect 14278 18320 14334 18329
rect 14016 17202 14044 18278
rect 14278 18255 14280 18264
rect 14332 18255 14334 18264
rect 14280 18226 14332 18232
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17270 14136 17614
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 13648 12406 13768 12434
rect 13912 12436 13964 12442
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13188 11898 13216 12174
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 10062 13032 11494
rect 13096 11082 13124 11698
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 10810 13124 11018
rect 13280 10810 13308 11766
rect 13556 11354 13584 11834
rect 13648 11762 13676 12406
rect 13912 12378 13964 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13464 10606 13492 11154
rect 13648 10674 13676 11698
rect 13740 11694 13768 12242
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13636 10668 13688 10674
rect 13556 10628 13636 10656
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13188 10198 13216 10406
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13372 10130 13400 10406
rect 13556 10130 13584 10628
rect 13636 10610 13688 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13832 10198 13860 10610
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13832 10062 13860 10134
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13280 9722 13308 9930
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13372 9722 13400 9862
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13372 9518 13400 9658
rect 13464 9586 13492 9862
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 12636 5914 12664 6938
rect 12820 6225 12848 7754
rect 12806 6216 12862 6225
rect 12806 6151 12862 6160
rect 12912 6118 12940 7754
rect 13464 7546 13492 9522
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 9042 13584 9318
rect 13832 9178 13860 9998
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13556 7449 13584 8978
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13924 7478 13952 7686
rect 13912 7472 13964 7478
rect 13542 7440 13598 7449
rect 13912 7414 13964 7420
rect 13542 7375 13598 7384
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 6390 13216 7142
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6390 13308 6598
rect 13924 6458 13952 6938
rect 14016 6474 14044 17002
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 14108 16522 14136 16662
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14200 6662 14228 17478
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 14292 15910 14320 16458
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 14006 14320 14350
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14292 13530 14320 13942
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14292 12850 14320 13466
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14292 12374 14320 12786
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14292 11898 14320 12310
rect 14384 11898 14412 19314
rect 14462 18728 14518 18737
rect 14462 18663 14518 18672
rect 14476 17882 14504 18663
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14568 17542 14596 19343
rect 14660 18086 14688 21966
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15290 21856 15346 21865
rect 14752 21486 14780 21830
rect 15120 21536 15148 21830
rect 15290 21791 15346 21800
rect 14844 21508 15148 21536
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14844 20874 14872 21508
rect 14945 21244 15253 21253
rect 14945 21242 14951 21244
rect 15007 21242 15031 21244
rect 15087 21242 15111 21244
rect 15167 21242 15191 21244
rect 15247 21242 15253 21244
rect 15007 21190 15009 21242
rect 15189 21190 15191 21242
rect 14945 21188 14951 21190
rect 15007 21188 15031 21190
rect 15087 21188 15111 21190
rect 15167 21188 15191 21190
rect 15247 21188 15253 21190
rect 14945 21179 15253 21188
rect 15304 21078 15332 21791
rect 15292 21072 15344 21078
rect 15292 21014 15344 21020
rect 15384 20936 15436 20942
rect 15382 20904 15384 20913
rect 15436 20904 15438 20913
rect 14832 20868 14884 20874
rect 15382 20839 15438 20848
rect 14832 20810 14884 20816
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14752 20398 14780 20742
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14752 20058 14780 20334
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14752 18426 14780 19314
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14844 17542 14872 20266
rect 14936 20262 14964 20742
rect 15488 20482 15516 21966
rect 15580 21350 15608 22034
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15672 21690 15700 21830
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15396 20454 15516 20482
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14945 20156 15253 20165
rect 14945 20154 14951 20156
rect 15007 20154 15031 20156
rect 15087 20154 15111 20156
rect 15167 20154 15191 20156
rect 15247 20154 15253 20156
rect 15007 20102 15009 20154
rect 15189 20102 15191 20154
rect 14945 20100 14951 20102
rect 15007 20100 15031 20102
rect 15087 20100 15111 20102
rect 15167 20100 15191 20102
rect 15247 20100 15253 20102
rect 14945 20091 15253 20100
rect 15200 20052 15252 20058
rect 15304 20040 15332 20334
rect 15252 20012 15332 20040
rect 15200 19994 15252 20000
rect 15212 19174 15240 19994
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14945 19068 15253 19077
rect 14945 19066 14951 19068
rect 15007 19066 15031 19068
rect 15087 19066 15111 19068
rect 15167 19066 15191 19068
rect 15247 19066 15253 19068
rect 15007 19014 15009 19066
rect 15189 19014 15191 19066
rect 14945 19012 14951 19014
rect 15007 19012 15031 19014
rect 15087 19012 15111 19014
rect 15167 19012 15191 19014
rect 15247 19012 15253 19014
rect 14945 19003 15253 19012
rect 15304 18970 15332 19722
rect 15396 19514 15424 20454
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15396 18766 15424 19110
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14936 18465 14964 18634
rect 14922 18456 14978 18465
rect 14922 18391 14978 18400
rect 15290 18320 15346 18329
rect 15290 18255 15346 18264
rect 14945 17980 15253 17989
rect 14945 17978 14951 17980
rect 15007 17978 15031 17980
rect 15087 17978 15111 17980
rect 15167 17978 15191 17980
rect 15247 17978 15253 17980
rect 15007 17926 15009 17978
rect 15189 17926 15191 17978
rect 14945 17924 14951 17926
rect 15007 17924 15031 17926
rect 15087 17924 15111 17926
rect 15167 17924 15191 17926
rect 15247 17924 15253 17926
rect 14945 17915 15253 17924
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14476 17202 14596 17218
rect 14464 17196 14596 17202
rect 14516 17190 14596 17196
rect 14464 17138 14516 17144
rect 14462 17096 14518 17105
rect 14462 17031 14464 17040
rect 14516 17031 14518 17040
rect 14464 17002 14516 17008
rect 14568 15910 14596 17190
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 12434 14596 15846
rect 14660 15706 14688 17138
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14844 15570 14872 17478
rect 15304 17338 15332 18255
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 14945 16892 15253 16901
rect 14945 16890 14951 16892
rect 15007 16890 15031 16892
rect 15087 16890 15111 16892
rect 15167 16890 15191 16892
rect 15247 16890 15253 16892
rect 15007 16838 15009 16890
rect 15189 16838 15191 16890
rect 14945 16836 14951 16838
rect 15007 16836 15031 16838
rect 15087 16836 15111 16838
rect 15167 16836 15191 16838
rect 15247 16836 15253 16838
rect 14945 16827 15253 16836
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15108 15904 15160 15910
rect 15160 15864 15332 15892
rect 15108 15846 15160 15852
rect 14945 15804 15253 15813
rect 14945 15802 14951 15804
rect 15007 15802 15031 15804
rect 15087 15802 15111 15804
rect 15167 15802 15191 15804
rect 15247 15802 15253 15804
rect 15007 15750 15009 15802
rect 15189 15750 15191 15802
rect 14945 15748 14951 15750
rect 15007 15748 15031 15750
rect 15087 15748 15111 15750
rect 15167 15748 15191 15750
rect 15247 15748 15253 15750
rect 14945 15739 15253 15748
rect 15304 15570 15332 15864
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 14945 14716 15253 14725
rect 14945 14714 14951 14716
rect 15007 14714 15031 14716
rect 15087 14714 15111 14716
rect 15167 14714 15191 14716
rect 15247 14714 15253 14716
rect 15007 14662 15009 14714
rect 15189 14662 15191 14714
rect 14945 14660 14951 14662
rect 15007 14660 15031 14662
rect 15087 14660 15111 14662
rect 15167 14660 15191 14662
rect 15247 14660 15253 14662
rect 14945 14651 15253 14660
rect 15014 14512 15070 14521
rect 15014 14447 15070 14456
rect 14648 14272 14700 14278
rect 14700 14232 14964 14260
rect 14648 14214 14700 14220
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14660 13297 14688 14010
rect 14936 13870 14964 14232
rect 15028 14006 15056 14447
rect 15396 14278 15424 16390
rect 15488 15706 15516 20334
rect 15580 20262 15608 21286
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 19854 15608 20198
rect 15672 20097 15700 20266
rect 15658 20088 15714 20097
rect 15658 20023 15714 20032
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15580 19446 15608 19790
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15580 18766 15608 19382
rect 15672 19174 15700 19790
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15580 18358 15608 18702
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15580 16182 15608 16390
rect 15568 16176 15620 16182
rect 15568 16118 15620 16124
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15672 15638 15700 17002
rect 15764 16232 15792 23800
rect 16120 22160 16172 22166
rect 16120 22102 16172 22108
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15844 21888 15896 21894
rect 15948 21865 15976 21898
rect 15844 21830 15896 21836
rect 15934 21856 15990 21865
rect 15856 21729 15884 21830
rect 15934 21791 15990 21800
rect 15842 21720 15898 21729
rect 15898 21678 15976 21706
rect 15842 21655 15898 21664
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 18068 15884 21422
rect 15948 21185 15976 21678
rect 16132 21554 16160 22102
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16304 21888 16356 21894
rect 16224 21848 16304 21876
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 15934 21176 15990 21185
rect 15934 21111 15990 21120
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15948 19854 15976 20742
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16040 19718 16068 20402
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15948 19378 15976 19654
rect 16118 19544 16174 19553
rect 16118 19479 16174 19488
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16040 18698 16068 19382
rect 16132 19378 16160 19479
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16132 18290 16160 18566
rect 16224 18358 16252 21848
rect 16304 21830 16356 21836
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 21593 16344 21626
rect 16302 21584 16358 21593
rect 16302 21519 16358 21528
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16316 21146 16344 21286
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16316 19922 16344 20810
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16120 18080 16172 18086
rect 15856 18040 16120 18068
rect 16120 18022 16172 18028
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16224 17241 16252 17274
rect 16210 17232 16266 17241
rect 16028 17196 16080 17202
rect 16210 17167 16266 17176
rect 16028 17138 16080 17144
rect 16040 16998 16068 17138
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15764 16204 15884 16232
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15488 15026 15516 15506
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15580 15162 15608 15302
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15672 15026 15700 15370
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15764 14822 15792 16050
rect 15856 15638 15884 16204
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15948 15570 15976 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15752 14816 15804 14822
rect 15672 14776 15752 14804
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15016 14000 15068 14006
rect 15212 13977 15240 14214
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15016 13942 15068 13948
rect 15198 13968 15254 13977
rect 15198 13903 15200 13912
rect 15252 13903 15254 13912
rect 15200 13874 15252 13880
rect 14924 13864 14976 13870
rect 15212 13843 15240 13874
rect 14924 13806 14976 13812
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 14945 13628 15253 13637
rect 14945 13626 14951 13628
rect 15007 13626 15031 13628
rect 15087 13626 15111 13628
rect 15167 13626 15191 13628
rect 15247 13626 15253 13628
rect 15007 13574 15009 13626
rect 15189 13574 15191 13626
rect 14945 13572 14951 13574
rect 15007 13572 15031 13574
rect 15087 13572 15111 13574
rect 15167 13572 15191 13574
rect 15247 13572 15253 13574
rect 14945 13563 15253 13572
rect 15108 13456 15160 13462
rect 15106 13424 15108 13433
rect 15160 13424 15162 13433
rect 15106 13359 15162 13368
rect 14646 13288 14702 13297
rect 14646 13223 14702 13232
rect 14476 12406 14596 12434
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14476 7546 14504 12406
rect 14660 11150 14688 13223
rect 14945 12540 15253 12549
rect 14945 12538 14951 12540
rect 15007 12538 15031 12540
rect 15087 12538 15111 12540
rect 15167 12538 15191 12540
rect 15247 12538 15253 12540
rect 15007 12486 15009 12538
rect 15189 12486 15191 12538
rect 14945 12484 14951 12486
rect 15007 12484 15031 12486
rect 15087 12484 15111 12486
rect 15167 12484 15191 12486
rect 15247 12484 15253 12486
rect 14945 12475 15253 12484
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15120 12238 15148 12310
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 14945 11452 15253 11461
rect 14945 11450 14951 11452
rect 15007 11450 15031 11452
rect 15087 11450 15111 11452
rect 15167 11450 15191 11452
rect 15247 11450 15253 11452
rect 15007 11398 15009 11450
rect 15189 11398 15191 11450
rect 14945 11396 14951 11398
rect 15007 11396 15031 11398
rect 15087 11396 15111 11398
rect 15167 11396 15191 11398
rect 15247 11396 15253 11398
rect 14945 11387 15253 11396
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 15120 10810 15148 11154
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 14844 8974 14872 10746
rect 14945 10364 15253 10373
rect 14945 10362 14951 10364
rect 15007 10362 15031 10364
rect 15087 10362 15111 10364
rect 15167 10362 15191 10364
rect 15247 10362 15253 10364
rect 15007 10310 15009 10362
rect 15189 10310 15191 10362
rect 14945 10308 14951 10310
rect 15007 10308 15031 10310
rect 15087 10308 15111 10310
rect 15167 10308 15191 10310
rect 15247 10308 15253 10310
rect 14945 10299 15253 10308
rect 14945 9276 15253 9285
rect 14945 9274 14951 9276
rect 15007 9274 15031 9276
rect 15087 9274 15111 9276
rect 15167 9274 15191 9276
rect 15247 9274 15253 9276
rect 15007 9222 15009 9274
rect 15189 9222 15191 9274
rect 14945 9220 14951 9222
rect 15007 9220 15031 9222
rect 15087 9220 15111 9222
rect 15167 9220 15191 9222
rect 15247 9220 15253 9222
rect 14945 9211 15253 9220
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14945 8188 15253 8197
rect 14945 8186 14951 8188
rect 15007 8186 15031 8188
rect 15087 8186 15111 8188
rect 15167 8186 15191 8188
rect 15247 8186 15253 8188
rect 15007 8134 15009 8186
rect 15189 8134 15191 8186
rect 14945 8132 14951 8134
rect 15007 8132 15031 8134
rect 15087 8132 15111 8134
rect 15167 8132 15191 8134
rect 15247 8132 15253 8134
rect 14945 8123 15253 8132
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 13912 6452 13964 6458
rect 14016 6446 14228 6474
rect 13912 6394 13964 6400
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 10784 5840 10836 5846
rect 11428 5840 11480 5846
rect 10784 5782 10836 5788
rect 11242 5808 11298 5817
rect 11428 5782 11480 5788
rect 11242 5743 11298 5752
rect 11256 5710 11284 5743
rect 11716 5710 11744 5850
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 12146 5468 12454 5477
rect 12146 5466 12152 5468
rect 12208 5466 12232 5468
rect 12288 5466 12312 5468
rect 12368 5466 12392 5468
rect 12448 5466 12454 5468
rect 12208 5414 12210 5466
rect 12390 5414 12392 5466
rect 12146 5412 12152 5414
rect 12208 5412 12232 5414
rect 12288 5412 12312 5414
rect 12368 5412 12392 5414
rect 12448 5412 12454 5414
rect 12146 5403 12454 5412
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10876 5296 10928 5302
rect 10796 5244 10876 5250
rect 10796 5238 10928 5244
rect 10796 5222 10916 5238
rect 10796 5166 10824 5222
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10428 4146 10456 4626
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10888 4146 10916 4422
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 10612 3534 10640 3878
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 3097 1440 3334
rect 5092 3126 5120 3470
rect 6548 3292 6856 3301
rect 6548 3290 6554 3292
rect 6610 3290 6634 3292
rect 6690 3290 6714 3292
rect 6770 3290 6794 3292
rect 6850 3290 6856 3292
rect 6610 3238 6612 3290
rect 6792 3238 6794 3290
rect 6548 3236 6554 3238
rect 6610 3236 6634 3238
rect 6690 3236 6714 3238
rect 6770 3236 6794 3238
rect 6850 3236 6856 3238
rect 6548 3227 6856 3236
rect 5080 3120 5132 3126
rect 1398 3088 1454 3097
rect 5080 3062 5132 3068
rect 11072 3058 11100 5306
rect 12146 4380 12454 4389
rect 12146 4378 12152 4380
rect 12208 4378 12232 4380
rect 12288 4378 12312 4380
rect 12368 4378 12392 4380
rect 12448 4378 12454 4380
rect 12208 4326 12210 4378
rect 12390 4326 12392 4378
rect 12146 4324 12152 4326
rect 12208 4324 12232 4326
rect 12288 4324 12312 4326
rect 12368 4324 12392 4326
rect 12448 4324 12454 4326
rect 12146 4315 12454 4324
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12544 3602 12572 3878
rect 12912 3670 12940 6054
rect 13188 5778 13216 6326
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13556 5778 13584 6054
rect 14108 5778 14136 6054
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13556 5370 13584 5510
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12146 3292 12454 3301
rect 12146 3290 12152 3292
rect 12208 3290 12232 3292
rect 12288 3290 12312 3292
rect 12368 3290 12392 3292
rect 12448 3290 12454 3292
rect 12208 3238 12210 3290
rect 12390 3238 12392 3290
rect 12146 3236 12152 3238
rect 12208 3236 12232 3238
rect 12288 3236 12312 3238
rect 12368 3236 12392 3238
rect 12448 3236 12454 3238
rect 12146 3227 12454 3236
rect 13004 3194 13032 3334
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 1398 3023 1454 3032
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 14200 2854 14228 6446
rect 14292 6390 14320 7142
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14292 6254 14320 6326
rect 14568 6254 14596 7414
rect 14660 7342 14688 7822
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14660 7002 14688 7278
rect 14945 7100 15253 7109
rect 14945 7098 14951 7100
rect 15007 7098 15031 7100
rect 15087 7098 15111 7100
rect 15167 7098 15191 7100
rect 15247 7098 15253 7100
rect 15007 7046 15009 7098
rect 15189 7046 15191 7098
rect 14945 7044 14951 7046
rect 15007 7044 15031 7046
rect 15087 7044 15111 7046
rect 15167 7044 15191 7046
rect 15247 7044 15253 7046
rect 14945 7035 15253 7044
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 15198 6760 15254 6769
rect 15198 6695 15200 6704
rect 15252 6695 15254 6704
rect 15200 6666 15252 6672
rect 14740 6656 14792 6662
rect 14792 6616 14872 6644
rect 14740 6598 14792 6604
rect 14844 6322 14872 6616
rect 14648 6316 14700 6322
rect 14832 6316 14884 6322
rect 14700 6276 14780 6304
rect 14648 6258 14700 6264
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14568 5778 14596 5850
rect 14752 5778 14780 6276
rect 14832 6258 14884 6264
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14384 5302 14412 5510
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14844 5166 14872 6258
rect 14945 6012 15253 6021
rect 14945 6010 14951 6012
rect 15007 6010 15031 6012
rect 15087 6010 15111 6012
rect 15167 6010 15191 6012
rect 15247 6010 15253 6012
rect 15007 5958 15009 6010
rect 15189 5958 15191 6010
rect 14945 5956 14951 5958
rect 15007 5956 15031 5958
rect 15087 5956 15111 5958
rect 15167 5956 15191 5958
rect 15247 5956 15253 5958
rect 14945 5947 15253 5956
rect 15304 5234 15332 13738
rect 15396 13530 15424 14010
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15396 12646 15424 12786
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15396 11898 15424 12582
rect 15488 12170 15516 14282
rect 15672 12434 15700 14776
rect 15752 14758 15804 14764
rect 15856 12434 15884 14826
rect 16040 13802 16068 16118
rect 16224 15706 16252 16730
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16132 13938 16160 14758
rect 16224 14550 16252 14962
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16224 14074 16252 14486
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16040 12714 16068 13194
rect 16224 12986 16252 14010
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16316 12918 16344 19654
rect 16408 19514 16436 20402
rect 16500 20233 16528 21286
rect 16486 20224 16542 20233
rect 16486 20159 16542 20168
rect 16592 19802 16620 21422
rect 16684 21010 16712 21966
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16670 20904 16726 20913
rect 16670 20839 16672 20848
rect 16724 20839 16726 20848
rect 16672 20810 16724 20816
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16500 19786 16620 19802
rect 16488 19780 16620 19786
rect 16540 19774 16620 19780
rect 16488 19722 16540 19728
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16486 19544 16542 19553
rect 16396 19508 16448 19514
rect 16486 19479 16542 19488
rect 16396 19450 16448 19456
rect 16394 19408 16450 19417
rect 16500 19378 16528 19479
rect 16592 19417 16620 19654
rect 16684 19514 16712 20334
rect 16776 19922 16804 23854
rect 16960 23746 16988 23854
rect 17038 23800 17094 24600
rect 17682 23800 17738 24600
rect 18326 23800 18382 24600
rect 18432 23854 18920 23882
rect 17052 23746 17080 23800
rect 16960 23718 17080 23746
rect 17592 22092 17644 22098
rect 17696 22094 17724 23800
rect 18340 23746 18368 23800
rect 18432 23746 18460 23854
rect 18340 23718 18460 23746
rect 18234 22536 18290 22545
rect 18234 22471 18290 22480
rect 18328 22500 18380 22506
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 17696 22066 17908 22094
rect 17592 22034 17644 22040
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17316 21956 17368 21962
rect 17316 21898 17368 21904
rect 16856 21616 16908 21622
rect 17144 21593 17172 21898
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 16856 21558 16908 21564
rect 17130 21584 17186 21593
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16868 19802 16896 21558
rect 17040 21548 17092 21554
rect 17130 21519 17186 21528
rect 17040 21490 17092 21496
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16960 20505 16988 20810
rect 17052 20777 17080 21490
rect 17132 20800 17184 20806
rect 17038 20768 17094 20777
rect 17132 20742 17184 20748
rect 17038 20703 17094 20712
rect 16946 20496 17002 20505
rect 16946 20431 17002 20440
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16776 19774 16896 19802
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16578 19408 16634 19417
rect 16394 19343 16396 19352
rect 16448 19343 16450 19352
rect 16488 19372 16540 19378
rect 16396 19314 16448 19320
rect 16578 19343 16634 19352
rect 16488 19314 16540 19320
rect 16578 19272 16634 19281
rect 16500 19230 16578 19258
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16408 18222 16436 18702
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16408 18086 16436 18158
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16408 17678 16436 18022
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16408 17270 16436 17614
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 14260 16436 16934
rect 16500 16182 16528 19230
rect 16578 19207 16634 19216
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16592 17490 16620 17818
rect 16684 17610 16712 19450
rect 16776 19446 16804 19774
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16592 17462 16712 17490
rect 16684 16998 16712 17462
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16590 16712 16934
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16592 16114 16620 16458
rect 16776 16402 16804 19246
rect 16684 16374 16804 16402
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16486 16008 16542 16017
rect 16486 15943 16488 15952
rect 16540 15943 16542 15952
rect 16488 15914 16540 15920
rect 16684 15910 16712 16374
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16670 15464 16726 15473
rect 16500 14890 16528 15438
rect 16670 15399 16726 15408
rect 16684 15366 16712 15399
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16578 15192 16634 15201
rect 16578 15127 16634 15136
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16488 14272 16540 14278
rect 16408 14240 16488 14260
rect 16540 14240 16542 14249
rect 16408 14232 16486 14240
rect 16486 14175 16542 14184
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16500 12918 16528 13806
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 16040 12434 16068 12650
rect 15580 12406 15700 12434
rect 15764 12406 15884 12434
rect 15948 12406 16068 12434
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15384 10736 15436 10742
rect 15488 10713 15516 11222
rect 15384 10678 15436 10684
rect 15474 10704 15530 10713
rect 15396 10198 15424 10678
rect 15474 10639 15530 10648
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15488 9586 15516 10639
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15396 5166 15424 6122
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14384 3602 14412 5034
rect 14844 4214 14872 5102
rect 14945 4924 15253 4933
rect 14945 4922 14951 4924
rect 15007 4922 15031 4924
rect 15087 4922 15111 4924
rect 15167 4922 15191 4924
rect 15247 4922 15253 4924
rect 15007 4870 15009 4922
rect 15189 4870 15191 4922
rect 14945 4868 14951 4870
rect 15007 4868 15031 4870
rect 15087 4868 15111 4870
rect 15167 4868 15191 4870
rect 15247 4868 15253 4870
rect 14945 4859 15253 4868
rect 15488 4690 15516 6054
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14945 3836 15253 3845
rect 14945 3834 14951 3836
rect 15007 3834 15031 3836
rect 15087 3834 15111 3836
rect 15167 3834 15191 3836
rect 15247 3834 15253 3836
rect 15007 3782 15009 3834
rect 15189 3782 15191 3834
rect 14945 3780 14951 3782
rect 15007 3780 15031 3782
rect 15087 3780 15111 3782
rect 15167 3780 15191 3782
rect 15247 3780 15253 3782
rect 14945 3771 15253 3780
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 15488 3534 15516 4626
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 3749 2748 4057 2757
rect 3749 2746 3755 2748
rect 3811 2746 3835 2748
rect 3891 2746 3915 2748
rect 3971 2746 3995 2748
rect 4051 2746 4057 2748
rect 3811 2694 3813 2746
rect 3993 2694 3995 2746
rect 3749 2692 3755 2694
rect 3811 2692 3835 2694
rect 3891 2692 3915 2694
rect 3971 2692 3995 2694
rect 4051 2692 4057 2694
rect 3749 2683 4057 2692
rect 4540 2446 4568 2790
rect 9347 2748 9655 2757
rect 9347 2746 9353 2748
rect 9409 2746 9433 2748
rect 9489 2746 9513 2748
rect 9569 2746 9593 2748
rect 9649 2746 9655 2748
rect 9409 2694 9411 2746
rect 9591 2694 9593 2746
rect 9347 2692 9353 2694
rect 9409 2692 9433 2694
rect 9489 2692 9513 2694
rect 9569 2692 9593 2694
rect 9649 2692 9655 2694
rect 9347 2683 9655 2692
rect 10612 2446 10640 2790
rect 15580 2774 15608 12406
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15672 11218 15700 11834
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 10198 15700 10610
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15672 9722 15700 10134
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15764 5148 15792 12406
rect 15948 11830 15976 12406
rect 16500 12374 16528 12854
rect 16592 12442 16620 15127
rect 16776 15026 16804 16186
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16672 14272 16724 14278
rect 16724 14232 16804 14260
rect 16672 14214 16724 14220
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11898 16528 12106
rect 16684 11898 16712 12582
rect 16776 12288 16804 14232
rect 16868 13870 16896 19654
rect 16960 18766 16988 20334
rect 17052 18970 17080 20402
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 17052 18290 17080 18906
rect 17144 18358 17172 20742
rect 17236 19802 17264 21830
rect 17328 19922 17356 21898
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17420 21162 17448 21830
rect 17512 21690 17540 21830
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17420 21134 17540 21162
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17420 20398 17448 20878
rect 17512 20534 17540 21134
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17420 19854 17448 20198
rect 17500 19984 17552 19990
rect 17604 19972 17632 22034
rect 17880 22012 17908 22066
rect 18052 22024 18104 22030
rect 17880 21984 18052 22012
rect 18052 21966 18104 21972
rect 18156 21962 18184 22374
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 18248 21894 18276 22471
rect 18328 22442 18380 22448
rect 18236 21888 18288 21894
rect 18234 21856 18236 21865
rect 18288 21856 18290 21865
rect 17744 21788 18052 21797
rect 18234 21791 18290 21800
rect 17744 21786 17750 21788
rect 17806 21786 17830 21788
rect 17886 21786 17910 21788
rect 17966 21786 17990 21788
rect 18046 21786 18052 21788
rect 17806 21734 17808 21786
rect 17988 21734 17990 21786
rect 17744 21732 17750 21734
rect 17806 21732 17830 21734
rect 17886 21732 17910 21734
rect 17966 21732 17990 21734
rect 18046 21732 18052 21734
rect 17744 21723 18052 21732
rect 18142 21720 18198 21729
rect 18064 21664 18142 21672
rect 18340 21690 18368 22442
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 18064 21655 18198 21664
rect 18328 21684 18380 21690
rect 18064 21644 18184 21655
rect 18064 21486 18092 21644
rect 18328 21626 18380 21632
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17744 20700 18052 20709
rect 17744 20698 17750 20700
rect 17806 20698 17830 20700
rect 17886 20698 17910 20700
rect 17966 20698 17990 20700
rect 18046 20698 18052 20700
rect 17806 20646 17808 20698
rect 17988 20646 17990 20698
rect 17744 20644 17750 20646
rect 17806 20644 17830 20646
rect 17886 20644 17910 20646
rect 17966 20644 17990 20646
rect 18046 20644 18052 20646
rect 17744 20635 18052 20644
rect 18156 20602 18184 21490
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 17868 20528 17920 20534
rect 17682 20496 17738 20505
rect 17682 20431 17738 20440
rect 17866 20496 17868 20505
rect 17920 20496 17922 20505
rect 17866 20431 17922 20440
rect 17696 20058 17724 20431
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 17972 20233 18000 20334
rect 17958 20224 18014 20233
rect 17958 20159 18014 20168
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17552 19944 17632 19972
rect 17500 19926 17552 19932
rect 17408 19848 17460 19854
rect 17236 19774 17356 19802
rect 17408 19790 17460 19796
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17236 19417 17264 19654
rect 17222 19408 17278 19417
rect 17222 19343 17278 19352
rect 17328 18426 17356 19774
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16946 18184 17002 18193
rect 16946 18119 17002 18128
rect 16960 17134 16988 18119
rect 17132 17672 17184 17678
rect 17420 17626 17448 19654
rect 17604 19446 17632 19944
rect 17958 19816 18014 19825
rect 17958 19751 17960 19760
rect 18012 19751 18014 19760
rect 17960 19722 18012 19728
rect 17744 19612 18052 19621
rect 17744 19610 17750 19612
rect 17806 19610 17830 19612
rect 17886 19610 17910 19612
rect 17966 19610 17990 19612
rect 18046 19610 18052 19612
rect 17806 19558 17808 19610
rect 17988 19558 17990 19610
rect 17744 19556 17750 19558
rect 17806 19556 17830 19558
rect 17886 19556 17910 19558
rect 17966 19556 17990 19558
rect 18046 19556 18052 19558
rect 17744 19547 18052 19556
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 18156 18970 18184 20334
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18064 18850 18092 18906
rect 18248 18850 18276 21286
rect 18340 20806 18368 21626
rect 18432 21486 18460 22102
rect 18788 22092 18840 22098
rect 18788 22034 18840 22040
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18432 21010 18460 21286
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18524 20942 18552 21490
rect 18512 20936 18564 20942
rect 18418 20904 18474 20913
rect 18512 20878 18564 20884
rect 18418 20839 18474 20848
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18326 20632 18382 20641
rect 18326 20567 18382 20576
rect 18340 20369 18368 20567
rect 18326 20360 18382 20369
rect 18326 20295 18382 20304
rect 18340 19553 18368 20295
rect 18326 19544 18382 19553
rect 18326 19479 18328 19488
rect 18380 19479 18382 19488
rect 18328 19450 18380 19456
rect 18064 18822 18184 18850
rect 18248 18822 18368 18850
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17132 17614 17184 17620
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16960 14618 16988 15370
rect 17052 15366 17080 16118
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16960 13870 16988 14554
rect 17052 14074 17080 15302
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 16856 12300 16908 12306
rect 16776 12260 16856 12288
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16132 10198 16160 10610
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16224 9178 16252 11698
rect 16684 11082 16712 11834
rect 16776 11558 16804 12260
rect 16856 12242 16908 12248
rect 17052 12102 17080 13126
rect 17144 12646 17172 17614
rect 17328 17598 17448 17626
rect 17328 17270 17356 17598
rect 17408 17536 17460 17542
rect 17406 17504 17408 17513
rect 17460 17504 17462 17513
rect 17406 17439 17462 17448
rect 17512 17338 17540 18634
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17604 18426 17632 18566
rect 17744 18524 18052 18533
rect 17744 18522 17750 18524
rect 17806 18522 17830 18524
rect 17886 18522 17910 18524
rect 17966 18522 17990 18524
rect 18046 18522 18052 18524
rect 17806 18470 17808 18522
rect 17988 18470 17990 18522
rect 17744 18468 17750 18470
rect 17806 18468 17830 18470
rect 17886 18468 17910 18470
rect 17966 18468 17990 18470
rect 18046 18468 18052 18470
rect 17744 18459 18052 18468
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17604 16590 17632 18022
rect 18064 17610 18092 18294
rect 18156 18086 18184 18822
rect 18340 18766 18368 18822
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 17744 17436 18052 17445
rect 17744 17434 17750 17436
rect 17806 17434 17830 17436
rect 17886 17434 17910 17436
rect 17966 17434 17990 17436
rect 18046 17434 18052 17436
rect 17806 17382 17808 17434
rect 17988 17382 17990 17434
rect 17744 17380 17750 17382
rect 17806 17380 17830 17382
rect 17886 17380 17910 17382
rect 17966 17380 17990 17382
rect 18046 17380 18052 17382
rect 17744 17371 18052 17380
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17788 16794 17816 17206
rect 18156 17202 18184 17546
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17744 16348 18052 16357
rect 17744 16346 17750 16348
rect 17806 16346 17830 16348
rect 17886 16346 17910 16348
rect 17966 16346 17990 16348
rect 18046 16346 18052 16348
rect 17806 16294 17808 16346
rect 17988 16294 17990 16346
rect 17744 16292 17750 16294
rect 17806 16292 17830 16294
rect 17886 16292 17910 16294
rect 17966 16292 17990 16294
rect 18046 16292 18052 16294
rect 17744 16283 18052 16292
rect 18248 16250 18276 18158
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18340 17338 18368 18090
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18340 17066 18368 17138
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18432 16946 18460 20839
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18524 19174 18552 20538
rect 18616 19718 18644 21830
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18524 17066 18552 19110
rect 18708 18970 18736 21830
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18604 18692 18656 18698
rect 18604 18634 18656 18640
rect 18616 18358 18644 18634
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18800 18086 18828 22034
rect 18892 20602 18920 23854
rect 18970 23800 19026 24600
rect 19614 23800 19670 24600
rect 20258 23800 20314 24600
rect 20902 23800 20958 24600
rect 21546 23800 21602 24600
rect 22190 23800 22246 24600
rect 22834 23800 22890 24600
rect 23478 23800 23534 24600
rect 24122 23800 24178 24600
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18878 20224 18934 20233
rect 18878 20159 18934 20168
rect 18892 18766 18920 20159
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18984 17882 19012 23800
rect 19628 22642 19656 23800
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 20168 22092 20220 22098
rect 20272 22094 20300 23800
rect 20543 22332 20851 22341
rect 20543 22330 20549 22332
rect 20605 22330 20629 22332
rect 20685 22330 20709 22332
rect 20765 22330 20789 22332
rect 20845 22330 20851 22332
rect 20605 22278 20607 22330
rect 20787 22278 20789 22330
rect 20543 22276 20549 22278
rect 20605 22276 20629 22278
rect 20685 22276 20709 22278
rect 20765 22276 20789 22278
rect 20845 22276 20851 22278
rect 20543 22267 20851 22276
rect 20812 22160 20864 22166
rect 20810 22128 20812 22137
rect 20864 22128 20866 22137
rect 20272 22066 20576 22094
rect 20168 22034 20220 22040
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 19076 21690 19104 21830
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 19168 21570 19196 22034
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19246 21720 19302 21729
rect 19246 21655 19302 21664
rect 19076 21542 19196 21570
rect 19260 21554 19288 21655
rect 19352 21554 19380 21898
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19430 21584 19486 21593
rect 19248 21548 19300 21554
rect 19076 20641 19104 21542
rect 19248 21490 19300 21496
rect 19340 21548 19392 21554
rect 19430 21519 19486 21528
rect 19340 21490 19392 21496
rect 19246 21312 19302 21321
rect 19246 21247 19302 21256
rect 19156 21004 19208 21010
rect 19156 20946 19208 20952
rect 19062 20632 19118 20641
rect 19168 20602 19196 20946
rect 19260 20913 19288 21247
rect 19246 20904 19302 20913
rect 19246 20839 19302 20848
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19062 20567 19118 20576
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19260 20534 19288 20742
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19076 20058 19104 20402
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19352 19854 19380 20198
rect 19340 19848 19392 19854
rect 19246 19816 19302 19825
rect 19340 19790 19392 19796
rect 19246 19751 19302 19760
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 19260 17814 19288 19751
rect 19444 19689 19472 21519
rect 19628 20641 19656 21830
rect 19720 21146 19748 21830
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19614 20632 19670 20641
rect 19614 20567 19670 20576
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19430 19680 19486 19689
rect 19430 19615 19486 19624
rect 19430 19544 19486 19553
rect 19628 19514 19656 19722
rect 19430 19479 19486 19488
rect 19616 19508 19668 19514
rect 19444 19378 19472 19479
rect 19616 19450 19668 19456
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19628 18970 19656 19450
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18358 19380 18702
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19706 18592 19762 18601
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19352 17678 19380 18294
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19340 17672 19392 17678
rect 18786 17640 18842 17649
rect 18604 17604 18656 17610
rect 19340 17614 19392 17620
rect 18786 17575 18842 17584
rect 18604 17546 18656 17552
rect 18616 17338 18644 17546
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18800 17270 18828 17575
rect 19444 17338 19472 18226
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 19064 17128 19116 17134
rect 19116 17076 19380 17082
rect 19064 17070 19380 17076
rect 18512 17060 18564 17066
rect 19076 17054 19380 17070
rect 18512 17002 18564 17008
rect 18340 16918 18460 16946
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15688 17356 15846
rect 17408 15700 17460 15706
rect 17328 15660 17408 15688
rect 17222 15600 17278 15609
rect 17222 15535 17278 15544
rect 17236 15162 17264 15535
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17328 14414 17356 15660
rect 17408 15642 17460 15648
rect 17590 15600 17646 15609
rect 18248 15570 18276 16186
rect 18340 15706 18368 16918
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 17590 15535 17646 15544
rect 18236 15564 18288 15570
rect 17604 14618 17632 15535
rect 18236 15506 18288 15512
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 17744 15260 18052 15269
rect 17744 15258 17750 15260
rect 17806 15258 17830 15260
rect 17886 15258 17910 15260
rect 17966 15258 17990 15260
rect 18046 15258 18052 15260
rect 17806 15206 17808 15258
rect 17988 15206 17990 15258
rect 17744 15204 17750 15206
rect 17806 15204 17830 15206
rect 17886 15204 17910 15206
rect 17966 15204 17990 15206
rect 18046 15204 18052 15206
rect 17744 15195 18052 15204
rect 18156 15026 18184 15438
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18156 14618 18184 14962
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17236 13530 17264 14282
rect 17328 13870 17356 14350
rect 17744 14172 18052 14181
rect 17744 14170 17750 14172
rect 17806 14170 17830 14172
rect 17886 14170 17910 14172
rect 17966 14170 17990 14172
rect 18046 14170 18052 14172
rect 17806 14118 17808 14170
rect 17988 14118 17990 14170
rect 17744 14116 17750 14118
rect 17806 14116 17830 14118
rect 17886 14116 17910 14118
rect 17966 14116 17990 14118
rect 18046 14116 18052 14118
rect 17744 14107 18052 14116
rect 18156 14006 18184 14554
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18524 13938 18552 16186
rect 18616 15434 18644 16730
rect 19352 16697 19380 17054
rect 19338 16688 19394 16697
rect 19338 16623 19394 16632
rect 19536 16590 19564 17818
rect 19628 17610 19656 18566
rect 19706 18527 19762 18536
rect 19616 17604 19668 17610
rect 19616 17546 19668 17552
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 18694 16280 18750 16289
rect 18694 16215 18750 16224
rect 18708 15978 18736 16215
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 19076 15434 19104 15982
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18786 15192 18842 15201
rect 18786 15127 18842 15136
rect 18800 14618 18828 15127
rect 19168 14958 19196 15846
rect 19260 15570 19288 16526
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19352 15162 19380 15846
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19338 15056 19394 15065
rect 19338 14991 19394 15000
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19352 14822 19380 14991
rect 19536 14890 19564 15642
rect 19720 15609 19748 18527
rect 19812 17338 19840 21626
rect 20074 21584 20130 21593
rect 20074 21519 20130 21528
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19904 20806 19932 21422
rect 19892 20800 19944 20806
rect 19892 20742 19944 20748
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19904 18290 19932 20334
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19996 17882 20024 21422
rect 20088 21185 20116 21519
rect 20074 21176 20130 21185
rect 20074 21111 20130 21120
rect 20180 18358 20208 22034
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 20364 21026 20392 21830
rect 20456 21690 20484 21830
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20548 21434 20576 22066
rect 20810 22063 20866 22072
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20640 21536 20668 21898
rect 20824 21842 20852 22063
rect 20916 21962 20944 23800
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 21272 21888 21324 21894
rect 20824 21814 21036 21842
rect 21272 21830 21324 21836
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 20812 21684 20864 21690
rect 20864 21644 20944 21672
rect 20812 21626 20864 21632
rect 20640 21508 20852 21536
rect 20548 21418 20760 21434
rect 20548 21412 20772 21418
rect 20548 21406 20720 21412
rect 20720 21354 20772 21360
rect 20824 21350 20852 21508
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20543 21244 20851 21253
rect 20543 21242 20549 21244
rect 20605 21242 20629 21244
rect 20685 21242 20709 21244
rect 20765 21242 20789 21244
rect 20845 21242 20851 21244
rect 20605 21190 20607 21242
rect 20787 21190 20789 21242
rect 20543 21188 20549 21190
rect 20605 21188 20629 21190
rect 20685 21188 20709 21190
rect 20765 21188 20789 21190
rect 20845 21188 20851 21190
rect 20543 21179 20851 21188
rect 20364 20998 20668 21026
rect 20916 21010 20944 21644
rect 21008 21146 21036 21814
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21100 21049 21128 21422
rect 21086 21040 21142 21049
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20272 19786 20300 20810
rect 20548 20346 20576 20878
rect 20456 20318 20576 20346
rect 20640 20330 20668 20998
rect 20904 21004 20956 21010
rect 21086 20975 21142 20984
rect 20904 20946 20956 20952
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20628 20324 20680 20330
rect 20456 19854 20484 20318
rect 20628 20266 20680 20272
rect 20543 20156 20851 20165
rect 20543 20154 20549 20156
rect 20605 20154 20629 20156
rect 20685 20154 20709 20156
rect 20765 20154 20789 20156
rect 20845 20154 20851 20156
rect 20605 20102 20607 20154
rect 20787 20102 20789 20154
rect 20543 20100 20549 20102
rect 20605 20100 20629 20102
rect 20685 20100 20709 20102
rect 20765 20100 20789 20102
rect 20845 20100 20851 20102
rect 20543 20091 20851 20100
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20444 19848 20496 19854
rect 20720 19848 20772 19854
rect 20444 19790 20496 19796
rect 20718 19816 20720 19825
rect 20772 19816 20774 19825
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 18698 20392 19654
rect 20456 19446 20484 19790
rect 20718 19751 20774 19760
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20456 18748 20484 19382
rect 20824 19258 20852 19994
rect 20916 19378 20944 20334
rect 21008 19553 21036 20878
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19990 21128 20198
rect 21088 19984 21140 19990
rect 21088 19926 21140 19932
rect 21086 19680 21142 19689
rect 21086 19615 21142 19624
rect 20994 19544 21050 19553
rect 21100 19514 21128 19615
rect 20994 19479 21050 19488
rect 21088 19508 21140 19514
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20824 19230 20944 19258
rect 20543 19068 20851 19077
rect 20543 19066 20549 19068
rect 20605 19066 20629 19068
rect 20685 19066 20709 19068
rect 20765 19066 20789 19068
rect 20845 19066 20851 19068
rect 20605 19014 20607 19066
rect 20787 19014 20789 19066
rect 20543 19012 20549 19014
rect 20605 19012 20629 19014
rect 20685 19012 20709 19014
rect 20765 19012 20789 19014
rect 20845 19012 20851 19014
rect 20543 19003 20851 19012
rect 20536 18760 20588 18766
rect 20456 18720 20536 18748
rect 20720 18760 20772 18766
rect 20536 18702 20588 18708
rect 20640 18708 20720 18714
rect 20640 18702 20772 18708
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20640 18686 20760 18702
rect 20640 18358 20668 18686
rect 20916 18442 20944 19230
rect 21008 18902 21036 19479
rect 21088 19450 21140 19456
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 20824 18414 20944 18442
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 20088 17270 20116 18158
rect 20180 18154 20208 18294
rect 20824 18193 20852 18414
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 20810 18184 20866 18193
rect 20168 18148 20220 18154
rect 20810 18119 20866 18128
rect 20168 18090 20220 18096
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 17338 20208 17546
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19812 16590 19840 17138
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19996 16250 20024 17138
rect 20088 17134 20116 17206
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 20088 16046 20116 17070
rect 20180 16182 20208 17274
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19706 15600 19762 15609
rect 19706 15535 19762 15544
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14618 19472 14758
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17236 12238 17264 13466
rect 17744 13084 18052 13093
rect 17744 13082 17750 13084
rect 17806 13082 17830 13084
rect 17886 13082 17910 13084
rect 17966 13082 17990 13084
rect 18046 13082 18052 13084
rect 17806 13030 17808 13082
rect 17988 13030 17990 13082
rect 17744 13028 17750 13030
rect 17806 13028 17830 13030
rect 17886 13028 17910 13030
rect 17966 13028 17990 13030
rect 18046 13028 18052 13030
rect 17744 13019 18052 13028
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16960 11694 16988 12038
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 17052 11354 17080 11698
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16868 10130 16896 11290
rect 17328 11218 17356 12922
rect 18156 12850 18184 13806
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18326 13016 18382 13025
rect 18326 12951 18328 12960
rect 18380 12951 18382 12960
rect 18328 12922 18380 12928
rect 18432 12850 18460 13466
rect 18616 13394 18644 13670
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18616 12782 18644 13330
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 12209 18000 12242
rect 18328 12232 18380 12238
rect 17958 12200 18014 12209
rect 18328 12174 18380 12180
rect 17958 12135 18014 12144
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17420 11898 17448 12038
rect 17744 11996 18052 12005
rect 17744 11994 17750 11996
rect 17806 11994 17830 11996
rect 17886 11994 17910 11996
rect 17966 11994 17990 11996
rect 18046 11994 18052 11996
rect 17806 11942 17808 11994
rect 17988 11942 17990 11994
rect 17744 11940 17750 11942
rect 17806 11940 17830 11942
rect 17886 11940 17910 11942
rect 17966 11940 17990 11942
rect 18046 11940 18052 11942
rect 17744 11931 18052 11940
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11354 18000 11698
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 18064 11121 18092 11494
rect 18156 11257 18184 12038
rect 18248 11830 18276 12038
rect 18340 11898 18368 12174
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18326 11792 18382 11801
rect 18326 11727 18328 11736
rect 18380 11727 18382 11736
rect 18328 11698 18380 11704
rect 18142 11248 18198 11257
rect 18142 11183 18198 11192
rect 18050 11112 18106 11121
rect 17592 11076 17644 11082
rect 18050 11047 18106 11056
rect 17592 11018 17644 11024
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 17040 10056 17092 10062
rect 16946 10024 17002 10033
rect 17040 9998 17092 10004
rect 16946 9959 17002 9968
rect 16960 9926 16988 9959
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 17052 9738 17080 9998
rect 17236 9926 17264 10610
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 16960 9722 17080 9738
rect 16960 9716 17092 9722
rect 16960 9710 17040 9716
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8498 16160 8774
rect 16764 8628 16816 8634
rect 16960 8616 16988 9710
rect 17040 9658 17092 9664
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16816 8588 16988 8616
rect 16764 8570 16816 8576
rect 17052 8566 17080 9522
rect 17144 8945 17172 9862
rect 17236 9518 17264 9862
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17130 8936 17186 8945
rect 17130 8871 17186 8880
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 15934 8392 15990 8401
rect 15934 8327 15936 8336
rect 15988 8327 15990 8336
rect 15936 8298 15988 8304
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15844 6656 15896 6662
rect 15948 6644 15976 7346
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 15896 6616 15976 6644
rect 15844 6598 15896 6604
rect 15842 6352 15898 6361
rect 15842 6287 15898 6296
rect 15672 5120 15792 5148
rect 15672 4078 15700 5120
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15856 3942 15884 6287
rect 15948 5166 15976 6616
rect 16040 6361 16068 6666
rect 16026 6352 16082 6361
rect 16026 6287 16082 6296
rect 16132 5778 16160 8434
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16224 7206 16252 7822
rect 16776 7750 16804 8434
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 7002 16252 7142
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16224 6798 16252 6938
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16316 5817 16344 6598
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16302 5808 16358 5817
rect 16120 5772 16172 5778
rect 16358 5766 16436 5794
rect 16302 5743 16358 5752
rect 16120 5714 16172 5720
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16224 5370 16252 5578
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15948 3602 15976 4218
rect 16040 4214 16068 5170
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4208 16080 4214
rect 16028 4150 16080 4156
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16040 3534 16068 4150
rect 16132 4010 16160 4966
rect 16224 4486 16252 5306
rect 16316 4690 16344 5510
rect 16408 5302 16436 5766
rect 16592 5710 16620 6394
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16592 4486 16620 5646
rect 16684 5370 16712 6326
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16132 3602 16160 3946
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16224 3398 16252 4422
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 4010 16344 4082
rect 16396 4072 16448 4078
rect 16672 4072 16724 4078
rect 16396 4014 16448 4020
rect 16670 4040 16672 4049
rect 16724 4040 16726 4049
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16408 2922 16436 4014
rect 16670 3975 16726 3984
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16500 3602 16528 3878
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16776 2990 16804 7686
rect 16960 6730 16988 7686
rect 17052 7478 17080 7686
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 17144 7290 17172 8871
rect 17328 8401 17356 9318
rect 17314 8392 17370 8401
rect 17314 8327 17370 8336
rect 17052 7262 17172 7290
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16960 5914 16988 6666
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16868 4128 16896 5510
rect 16948 4140 17000 4146
rect 16868 4100 16948 4128
rect 16948 4082 17000 4088
rect 17052 4078 17080 7262
rect 17512 6662 17540 9522
rect 17604 9489 17632 11018
rect 17744 10908 18052 10917
rect 17744 10906 17750 10908
rect 17806 10906 17830 10908
rect 17886 10906 17910 10908
rect 17966 10906 17990 10908
rect 18046 10906 18052 10908
rect 17806 10854 17808 10906
rect 17988 10854 17990 10906
rect 17744 10852 17750 10854
rect 17806 10852 17830 10854
rect 17886 10852 17910 10854
rect 17966 10852 17990 10854
rect 18046 10852 18052 10854
rect 17744 10843 18052 10852
rect 18432 10198 18460 12582
rect 18512 12436 18564 12442
rect 18616 12434 18644 12718
rect 18616 12406 18736 12434
rect 18512 12378 18564 12384
rect 18524 11642 18552 12378
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18616 11898 18644 12174
rect 18708 12170 18736 12406
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18708 11762 18736 12106
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18800 11830 18828 12038
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18524 11614 18736 11642
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 17744 9820 18052 9829
rect 17744 9818 17750 9820
rect 17806 9818 17830 9820
rect 17886 9818 17910 9820
rect 17966 9818 17990 9820
rect 18046 9818 18052 9820
rect 17806 9766 17808 9818
rect 17988 9766 17990 9818
rect 17744 9764 17750 9766
rect 17806 9764 17830 9766
rect 17886 9764 17910 9766
rect 17966 9764 17990 9766
rect 18046 9764 18052 9766
rect 17744 9755 18052 9764
rect 18340 9761 18368 9930
rect 18326 9752 18382 9761
rect 18326 9687 18382 9696
rect 17774 9616 17830 9625
rect 17774 9551 17776 9560
rect 17828 9551 17830 9560
rect 17776 9522 17828 9528
rect 17590 9480 17646 9489
rect 17590 9415 17646 9424
rect 17776 9376 17828 9382
rect 17828 9324 18000 9330
rect 17776 9318 18000 9324
rect 17788 9302 18000 9318
rect 17972 8906 18000 9302
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17744 8732 18052 8741
rect 17744 8730 17750 8732
rect 17806 8730 17830 8732
rect 17886 8730 17910 8732
rect 17966 8730 17990 8732
rect 18046 8730 18052 8732
rect 17806 8678 17808 8730
rect 17988 8678 17990 8730
rect 17744 8676 17750 8678
rect 17806 8676 17830 8678
rect 17886 8676 17910 8678
rect 17966 8676 17990 8678
rect 18046 8676 18052 8678
rect 17744 8667 18052 8676
rect 18156 8430 18184 8910
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18052 7744 18104 7750
rect 18104 7704 18184 7732
rect 18052 7686 18104 7692
rect 17744 7644 18052 7653
rect 17744 7642 17750 7644
rect 17806 7642 17830 7644
rect 17886 7642 17910 7644
rect 17966 7642 17990 7644
rect 18046 7642 18052 7644
rect 17806 7590 17808 7642
rect 17988 7590 17990 7642
rect 17744 7588 17750 7590
rect 17806 7588 17830 7590
rect 17886 7588 17910 7590
rect 17966 7588 17990 7590
rect 18046 7588 18052 7590
rect 17744 7579 18052 7588
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17972 7154 18000 7482
rect 18156 7313 18184 7704
rect 18248 7546 18276 8774
rect 18340 7993 18368 8842
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18326 7984 18382 7993
rect 18326 7919 18382 7928
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18142 7304 18198 7313
rect 18142 7239 18144 7248
rect 18196 7239 18198 7248
rect 18144 7210 18196 7216
rect 17604 6798 17632 7142
rect 17972 7126 18184 7154
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17144 6118 17172 6326
rect 17604 6322 17632 6734
rect 18156 6633 18184 7126
rect 18142 6624 18198 6633
rect 17744 6556 18052 6565
rect 18142 6559 18198 6568
rect 17744 6554 17750 6556
rect 17806 6554 17830 6556
rect 17886 6554 17910 6556
rect 17966 6554 17990 6556
rect 18046 6554 18052 6556
rect 17806 6502 17808 6554
rect 17988 6502 17990 6554
rect 17744 6500 17750 6502
rect 17806 6500 17830 6502
rect 17886 6500 17910 6502
rect 17966 6500 17990 6502
rect 18046 6500 18052 6502
rect 17744 6491 18052 6500
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17144 5710 17172 6054
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17236 4146 17264 5782
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17328 4214 17356 5170
rect 17420 4622 17448 6190
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 5370 17540 5714
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17604 4826 17632 5646
rect 17744 5468 18052 5477
rect 17744 5466 17750 5468
rect 17806 5466 17830 5468
rect 17886 5466 17910 5468
rect 17966 5466 17990 5468
rect 18046 5466 18052 5468
rect 17806 5414 17808 5466
rect 17988 5414 17990 5466
rect 17744 5412 17750 5414
rect 17806 5412 17830 5414
rect 17886 5412 17910 5414
rect 17966 5412 17990 5414
rect 18046 5412 18052 5414
rect 17744 5403 18052 5412
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17744 4380 18052 4389
rect 17744 4378 17750 4380
rect 17806 4378 17830 4380
rect 17886 4378 17910 4380
rect 17966 4378 17990 4380
rect 18046 4378 18052 4380
rect 17806 4326 17808 4378
rect 17988 4326 17990 4378
rect 17744 4324 17750 4326
rect 17806 4324 17830 4326
rect 17886 4324 17910 4326
rect 17966 4324 17990 4326
rect 18046 4324 18052 4326
rect 17744 4315 18052 4324
rect 17316 4208 17368 4214
rect 17316 4150 17368 4156
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 17236 3738 17264 4082
rect 17328 4026 17356 4150
rect 17328 3998 17448 4026
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 3194 17356 3334
rect 17420 3194 17448 3998
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3602 18092 3878
rect 18156 3602 18184 6394
rect 18248 4690 18276 7482
rect 18340 6866 18368 7686
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18236 4548 18288 4554
rect 18340 4536 18368 6598
rect 18288 4508 18368 4536
rect 18236 4490 18288 4496
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18340 3534 18368 4508
rect 18432 4078 18460 8570
rect 18524 7585 18552 10950
rect 18616 9178 18644 11494
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18708 7750 18736 11614
rect 18892 7886 18920 14486
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19168 13258 19196 14350
rect 19444 14226 19472 14554
rect 19536 14414 19564 14826
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19444 14198 19564 14226
rect 19338 13424 19394 13433
rect 19338 13359 19394 13368
rect 19352 13326 19380 13359
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19064 13184 19116 13190
rect 19444 13161 19472 13194
rect 19064 13126 19116 13132
rect 19430 13152 19486 13161
rect 19076 12889 19104 13126
rect 19430 13087 19486 13096
rect 19062 12880 19118 12889
rect 19062 12815 19118 12824
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19062 12744 19118 12753
rect 19062 12679 19118 12688
rect 19076 12646 19104 12679
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19352 12345 19380 12786
rect 19338 12336 19394 12345
rect 19338 12271 19394 12280
rect 19340 12232 19392 12238
rect 19392 12192 19472 12220
rect 19340 12174 19392 12180
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11354 19288 11698
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19064 11280 19116 11286
rect 19340 11280 19392 11286
rect 19064 11222 19116 11228
rect 19338 11248 19340 11257
rect 19392 11248 19394 11257
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18984 9654 19012 10950
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 9382 19012 9454
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18510 7576 18566 7585
rect 18510 7511 18566 7520
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18524 6254 18552 6802
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18616 5710 18644 6666
rect 18708 6458 18736 6938
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18708 5030 18736 6258
rect 18800 6118 18828 7414
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18800 5302 18828 6054
rect 18788 5296 18840 5302
rect 18788 5238 18840 5244
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18708 4622 18736 4966
rect 18892 4690 18920 7346
rect 18984 6304 19012 9318
rect 19076 9110 19104 11222
rect 19338 11183 19394 11192
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19168 10674 19196 10950
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19260 10169 19288 11018
rect 19352 10849 19380 11086
rect 19338 10840 19394 10849
rect 19338 10775 19394 10784
rect 19444 10742 19472 12192
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19246 10160 19302 10169
rect 19246 10095 19302 10104
rect 19340 10056 19392 10062
rect 19444 10044 19472 10678
rect 19536 10062 19564 14198
rect 19628 14074 19656 14962
rect 19798 14920 19854 14929
rect 19798 14855 19854 14864
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19812 14006 19840 14855
rect 20088 14822 20116 15982
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19800 14000 19852 14006
rect 19706 13968 19762 13977
rect 19800 13942 19852 13948
rect 19706 13903 19762 13912
rect 19720 13190 19748 13903
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19628 12170 19656 13126
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11937 19840 12038
rect 19798 11928 19854 11937
rect 19798 11863 19854 11872
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19812 10062 19840 10406
rect 19392 10016 19472 10044
rect 19524 10056 19576 10062
rect 19340 9998 19392 10004
rect 19524 9998 19576 10004
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19338 9888 19394 9897
rect 19338 9823 19394 9832
rect 19352 9722 19380 9823
rect 19706 9752 19762 9761
rect 19340 9716 19392 9722
rect 19706 9687 19762 9696
rect 19340 9658 19392 9664
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 19168 8809 19196 9590
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 9081 19380 9318
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19154 8800 19210 8809
rect 19154 8735 19210 8744
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19168 8430 19196 8570
rect 19338 8528 19394 8537
rect 19248 8492 19300 8498
rect 19338 8463 19394 8472
rect 19248 8434 19300 8440
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19260 7750 19288 8434
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19156 7200 19208 7206
rect 19062 7168 19118 7177
rect 19156 7142 19208 7148
rect 19062 7103 19118 7112
rect 19076 6644 19104 7103
rect 19168 7041 19196 7142
rect 19154 7032 19210 7041
rect 19260 7002 19288 7686
rect 19352 7177 19380 8463
rect 19444 7478 19472 8978
rect 19522 8664 19578 8673
rect 19522 8599 19524 8608
rect 19576 8599 19578 8608
rect 19524 8570 19576 8576
rect 19628 8430 19656 9590
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19628 8294 19656 8366
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19338 7168 19394 7177
rect 19338 7103 19394 7112
rect 19154 6967 19210 6976
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19156 6792 19208 6798
rect 19248 6792 19300 6798
rect 19208 6752 19248 6780
rect 19156 6734 19208 6740
rect 19248 6734 19300 6740
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19156 6656 19208 6662
rect 19076 6616 19156 6644
rect 19156 6598 19208 6604
rect 19248 6316 19300 6322
rect 18984 6276 19248 6304
rect 19248 6258 19300 6264
rect 18972 6112 19024 6118
rect 18970 6080 18972 6089
rect 19024 6080 19026 6089
rect 18970 6015 19026 6024
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18984 4486 19012 6015
rect 19062 5944 19118 5953
rect 19062 5879 19118 5888
rect 19076 5846 19104 5879
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19168 5370 19196 5510
rect 19352 5409 19380 6666
rect 19430 6488 19486 6497
rect 19430 6423 19486 6432
rect 19338 5400 19394 5409
rect 19156 5364 19208 5370
rect 19338 5335 19394 5344
rect 19156 5306 19208 5312
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18708 4282 18736 4422
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 19246 4176 19302 4185
rect 19246 4111 19302 4120
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 19168 3398 19196 3538
rect 18512 3392 18564 3398
rect 18510 3360 18512 3369
rect 19156 3392 19208 3398
rect 18564 3360 18566 3369
rect 19156 3334 19208 3340
rect 17744 3292 18052 3301
rect 18510 3295 18566 3304
rect 17744 3290 17750 3292
rect 17806 3290 17830 3292
rect 17886 3290 17910 3292
rect 17966 3290 17990 3292
rect 18046 3290 18052 3292
rect 17806 3238 17808 3290
rect 17988 3238 17990 3290
rect 17744 3236 17750 3238
rect 17806 3236 17830 3238
rect 17886 3236 17910 3238
rect 17966 3236 17990 3238
rect 18046 3236 18052 3238
rect 17744 3227 18052 3236
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 14945 2748 15253 2757
rect 14945 2746 14951 2748
rect 15007 2746 15031 2748
rect 15087 2746 15111 2748
rect 15167 2746 15191 2748
rect 15247 2746 15253 2748
rect 15007 2694 15009 2746
rect 15189 2694 15191 2746
rect 14945 2692 14951 2694
rect 15007 2692 15031 2694
rect 15087 2692 15111 2694
rect 15167 2692 15191 2694
rect 15247 2692 15253 2694
rect 14945 2683 15253 2692
rect 15488 2746 15608 2774
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 800 2176 2246
rect 6196 800 6224 2382
rect 15488 2310 15516 2746
rect 19260 2582 19288 4111
rect 19352 3738 19380 4490
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19352 2990 19380 3470
rect 19444 3126 19472 6423
rect 19536 4978 19564 7958
rect 19628 7750 19656 8230
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19720 7698 19748 9687
rect 19904 8838 19932 14282
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19996 12714 20024 13874
rect 20088 13734 20116 14758
rect 20272 14521 20300 18022
rect 20543 17980 20851 17989
rect 20543 17978 20549 17980
rect 20605 17978 20629 17980
rect 20685 17978 20709 17980
rect 20765 17978 20789 17980
rect 20845 17978 20851 17980
rect 20605 17926 20607 17978
rect 20787 17926 20789 17978
rect 20543 17924 20549 17926
rect 20605 17924 20629 17926
rect 20685 17924 20709 17926
rect 20765 17924 20789 17926
rect 20845 17924 20851 17926
rect 20543 17915 20851 17924
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20364 16250 20392 17546
rect 20456 16794 20484 17818
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17270 20760 17614
rect 21008 17338 21036 18226
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20543 16892 20851 16901
rect 20543 16890 20549 16892
rect 20605 16890 20629 16892
rect 20685 16890 20709 16892
rect 20765 16890 20789 16892
rect 20845 16890 20851 16892
rect 20605 16838 20607 16890
rect 20787 16838 20789 16890
rect 20543 16836 20549 16838
rect 20605 16836 20629 16838
rect 20685 16836 20709 16838
rect 20765 16836 20789 16838
rect 20845 16836 20851 16838
rect 20543 16827 20851 16836
rect 20916 16794 20944 17002
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20640 16425 20668 16458
rect 21008 16454 21036 17138
rect 21100 16998 21128 17478
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21086 16552 21142 16561
rect 21086 16487 21142 16496
rect 20996 16448 21048 16454
rect 20626 16416 20682 16425
rect 20996 16390 21048 16396
rect 20626 16351 20682 16360
rect 21100 16250 21128 16487
rect 21192 16289 21220 20742
rect 21284 20058 21312 21830
rect 21376 21690 21404 21830
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21468 21554 21496 22442
rect 21560 21690 21588 23800
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 22020 22234 22048 22578
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 21548 21684 21600 21690
rect 21548 21626 21600 21632
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21376 21457 21404 21490
rect 21362 21448 21418 21457
rect 21362 21383 21418 21392
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21362 20496 21418 20505
rect 21362 20431 21364 20440
rect 21416 20431 21418 20440
rect 21364 20402 21416 20408
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21376 19514 21404 20198
rect 21468 19854 21496 21082
rect 21546 20632 21602 20641
rect 21546 20567 21548 20576
rect 21600 20567 21602 20576
rect 21548 20538 21600 20544
rect 21456 19848 21508 19854
rect 21508 19808 21588 19836
rect 21456 19790 21508 19796
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 19514 21496 19654
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21270 19408 21326 19417
rect 21560 19394 21588 19808
rect 21270 19343 21272 19352
rect 21324 19343 21326 19352
rect 21468 19366 21588 19394
rect 21272 19314 21324 19320
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18154 21312 19110
rect 21272 18148 21324 18154
rect 21272 18090 21324 18096
rect 21468 17954 21496 19366
rect 21652 19174 21680 22170
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21744 19310 21772 22102
rect 22204 22094 22232 23800
rect 22374 22128 22430 22137
rect 22284 22094 22336 22098
rect 22204 22092 22336 22094
rect 22204 22066 22284 22092
rect 22374 22063 22430 22072
rect 22284 22034 22336 22040
rect 21824 22024 21876 22030
rect 21822 21992 21824 22001
rect 22100 22024 22152 22030
rect 21876 21992 21878 22001
rect 22296 22003 22324 22034
rect 22100 21966 22152 21972
rect 21822 21927 21878 21936
rect 21916 21616 21968 21622
rect 21968 21576 22048 21604
rect 21916 21558 21968 21564
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21836 19334 21864 21014
rect 22020 20806 22048 21576
rect 22112 20913 22140 21966
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22098 20904 22154 20913
rect 22204 20874 22232 21490
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22098 20839 22154 20848
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22296 20584 22324 20878
rect 22388 20602 22416 22063
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22572 21865 22600 21966
rect 22558 21856 22614 21865
rect 22558 21791 22614 21800
rect 22848 21690 22876 23800
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22466 21584 22522 21593
rect 22466 21519 22468 21528
rect 22520 21519 22522 21528
rect 22650 21584 22706 21593
rect 22650 21519 22706 21528
rect 22744 21548 22796 21554
rect 22468 21490 22520 21496
rect 22664 21146 22692 21519
rect 22744 21490 22796 21496
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22020 20556 22324 20584
rect 22376 20596 22428 20602
rect 21732 19304 21784 19310
rect 21836 19306 21956 19334
rect 21732 19246 21784 19252
rect 21833 19236 21885 19242
rect 21833 19178 21885 19184
rect 21640 19168 21692 19174
rect 21560 19128 21640 19156
rect 21560 18086 21588 19128
rect 21640 19110 21692 19116
rect 21732 19168 21784 19174
rect 21845 19122 21873 19178
rect 21732 19110 21784 19116
rect 21744 18442 21772 19110
rect 21652 18414 21772 18442
rect 21836 19094 21873 19122
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21468 17926 21588 17954
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21376 17746 21404 17818
rect 21560 17762 21588 17926
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21468 17734 21588 17762
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 16590 21312 17478
rect 21376 17270 21404 17682
rect 21364 17264 21416 17270
rect 21364 17206 21416 17212
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21376 16998 21404 17070
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21376 16289 21404 16594
rect 21178 16280 21234 16289
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 21088 16244 21140 16250
rect 21178 16215 21234 16224
rect 21362 16280 21418 16289
rect 21362 16215 21418 16224
rect 21088 16186 21140 16192
rect 20364 15706 20392 16186
rect 21086 16144 21142 16153
rect 20904 16108 20956 16114
rect 21086 16079 21142 16088
rect 21270 16144 21326 16153
rect 21270 16079 21272 16088
rect 20904 16050 20956 16056
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20456 15434 20484 15982
rect 20543 15804 20851 15813
rect 20543 15802 20549 15804
rect 20605 15802 20629 15804
rect 20685 15802 20709 15804
rect 20765 15802 20789 15804
rect 20845 15802 20851 15804
rect 20605 15750 20607 15802
rect 20787 15750 20789 15802
rect 20543 15748 20549 15750
rect 20605 15748 20629 15750
rect 20685 15748 20709 15750
rect 20765 15748 20789 15750
rect 20845 15748 20851 15750
rect 20543 15739 20851 15748
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20548 15434 20576 15574
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20456 14618 20484 15370
rect 20916 15366 20944 16050
rect 21100 15366 21128 16079
rect 21324 16079 21326 16088
rect 21272 16050 21324 16056
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 20543 14716 20851 14725
rect 20543 14714 20549 14716
rect 20605 14714 20629 14716
rect 20685 14714 20709 14716
rect 20765 14714 20789 14716
rect 20845 14714 20851 14716
rect 20605 14662 20607 14714
rect 20787 14662 20789 14714
rect 20543 14660 20549 14662
rect 20605 14660 20629 14662
rect 20685 14660 20709 14662
rect 20765 14660 20789 14662
rect 20845 14660 20851 14662
rect 20543 14651 20851 14660
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 21100 14550 21128 14894
rect 21088 14544 21140 14550
rect 20258 14512 20314 14521
rect 21088 14486 21140 14492
rect 20258 14447 20314 14456
rect 21192 14278 21220 15302
rect 21284 14482 21312 15506
rect 21468 14498 21496 17734
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21560 16561 21588 17614
rect 21652 17066 21680 18414
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 21744 17882 21772 18294
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21836 17785 21864 19094
rect 21928 18630 21956 19306
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21928 18086 21956 18566
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21822 17776 21878 17785
rect 21822 17711 21878 17720
rect 22020 17592 22048 20556
rect 22376 20538 22428 20544
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22112 17746 22140 19858
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 21744 17564 22048 17592
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21546 16552 21602 16561
rect 21744 16538 21772 17564
rect 21822 17504 21878 17513
rect 21822 17439 21878 17448
rect 21546 16487 21602 16496
rect 21652 16510 21772 16538
rect 21652 15586 21680 16510
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21744 16046 21772 16390
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21836 15706 21864 17439
rect 22112 17270 22140 17682
rect 22204 17649 22232 20402
rect 22756 20074 22784 21490
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 23032 21049 23060 21286
rect 23018 21040 23074 21049
rect 23018 20975 23074 20984
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 23032 20505 23060 20742
rect 23018 20496 23074 20505
rect 22928 20460 22980 20466
rect 23018 20431 23074 20440
rect 22928 20402 22980 20408
rect 22664 20046 22784 20074
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22296 18737 22324 19654
rect 22282 18728 22338 18737
rect 22282 18663 22338 18672
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22296 18426 22324 18566
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22388 18329 22416 19654
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22374 18320 22430 18329
rect 22374 18255 22430 18264
rect 22480 18222 22508 19246
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22480 17882 22508 18158
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22190 17640 22246 17649
rect 22190 17575 22246 17584
rect 22284 17604 22336 17610
rect 22284 17546 22336 17552
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16658 22048 16934
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 21928 16114 21956 16458
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21916 15972 21968 15978
rect 22020 15960 22048 16594
rect 21968 15932 22048 15960
rect 21916 15914 21968 15920
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21560 15558 21680 15586
rect 21836 15570 21864 15642
rect 22020 15638 22048 15932
rect 22112 15638 22140 17070
rect 22204 16794 22232 17478
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22296 16250 22324 17546
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 17270 22508 17478
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22376 16448 22428 16454
rect 22374 16416 22376 16425
rect 22428 16416 22430 16425
rect 22374 16351 22430 16360
rect 22374 16280 22430 16289
rect 22284 16244 22336 16250
rect 22374 16215 22430 16224
rect 22284 16186 22336 16192
rect 22388 16182 22416 16215
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22480 16114 22508 17206
rect 22572 17202 22600 19654
rect 22664 17241 22692 20046
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 22834 19952 22890 19961
rect 22756 18834 22784 19926
rect 22834 19887 22890 19896
rect 22848 19854 22876 19887
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22756 18426 22784 18770
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22742 17640 22798 17649
rect 22742 17575 22798 17584
rect 22650 17232 22706 17241
rect 22560 17196 22612 17202
rect 22650 17167 22706 17176
rect 22560 17138 22612 17144
rect 22572 16726 22600 17138
rect 22756 17105 22784 17575
rect 22742 17096 22798 17105
rect 22742 17031 22798 17040
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22572 16250 22600 16526
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22388 15706 22416 15982
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 21824 15564 21876 15570
rect 21560 15201 21588 15558
rect 21824 15506 21876 15512
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21546 15192 21602 15201
rect 21652 15162 21680 15438
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21546 15127 21602 15136
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21730 15056 21786 15065
rect 21730 14991 21732 15000
rect 21784 14991 21786 15000
rect 21732 14962 21784 14968
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21376 14470 21496 14498
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20088 13326 20116 13670
rect 20543 13628 20851 13637
rect 20543 13626 20549 13628
rect 20605 13626 20629 13628
rect 20685 13626 20709 13628
rect 20765 13626 20789 13628
rect 20845 13626 20851 13628
rect 20605 13574 20607 13626
rect 20787 13574 20789 13626
rect 20543 13572 20549 13574
rect 20605 13572 20629 13574
rect 20685 13572 20709 13574
rect 20765 13572 20789 13574
rect 20845 13572 20851 13574
rect 20543 13563 20851 13572
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19984 12232 20036 12238
rect 20088 12220 20116 13262
rect 20916 13258 20944 14010
rect 21284 14006 21312 14418
rect 21376 14385 21404 14470
rect 21456 14408 21508 14414
rect 21362 14376 21418 14385
rect 21456 14350 21508 14356
rect 21362 14311 21418 14320
rect 21272 14000 21324 14006
rect 21272 13942 21324 13948
rect 21284 13818 21312 13942
rect 21468 13938 21496 14350
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21284 13790 21404 13818
rect 21086 13288 21142 13297
rect 20904 13252 20956 13258
rect 21086 13223 21088 13232
rect 20904 13194 20956 13200
rect 21140 13223 21142 13232
rect 21088 13194 21140 13200
rect 21086 13016 21142 13025
rect 21086 12951 21142 12960
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20036 12192 20116 12220
rect 19984 12174 20036 12180
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19996 11665 20024 11834
rect 19982 11656 20038 11665
rect 19982 11591 20038 11600
rect 20272 10656 20300 12038
rect 20364 11898 20392 12786
rect 20543 12540 20851 12549
rect 20543 12538 20549 12540
rect 20605 12538 20629 12540
rect 20685 12538 20709 12540
rect 20765 12538 20789 12540
rect 20845 12538 20851 12540
rect 20605 12486 20607 12538
rect 20787 12486 20789 12538
rect 20543 12484 20549 12486
rect 20605 12484 20629 12486
rect 20685 12484 20709 12486
rect 20765 12484 20789 12486
rect 20845 12484 20851 12486
rect 20543 12475 20851 12484
rect 20994 12064 21050 12073
rect 20994 11999 21050 12008
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 21008 11830 21036 11999
rect 21100 11898 21128 12951
rect 21178 12880 21234 12889
rect 21178 12815 21234 12824
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20364 11150 20392 11494
rect 20543 11452 20851 11461
rect 20543 11450 20549 11452
rect 20605 11450 20629 11452
rect 20685 11450 20709 11452
rect 20765 11450 20789 11452
rect 20845 11450 20851 11452
rect 20605 11398 20607 11450
rect 20787 11398 20789 11450
rect 20543 11396 20549 11398
rect 20605 11396 20629 11398
rect 20685 11396 20709 11398
rect 20765 11396 20789 11398
rect 20845 11396 20851 11398
rect 20543 11387 20851 11396
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20902 11112 20958 11121
rect 20640 10742 20668 11086
rect 20902 11047 20958 11056
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20352 10668 20404 10674
rect 20272 10628 20352 10656
rect 20352 10610 20404 10616
rect 20543 10364 20851 10373
rect 20543 10362 20549 10364
rect 20605 10362 20629 10364
rect 20685 10362 20709 10364
rect 20765 10362 20789 10364
rect 20845 10362 20851 10364
rect 20605 10310 20607 10362
rect 20787 10310 20789 10362
rect 20543 10308 20549 10310
rect 20605 10308 20629 10310
rect 20685 10308 20709 10310
rect 20765 10308 20789 10310
rect 20845 10308 20851 10310
rect 20543 10299 20851 10308
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20364 9586 20392 10202
rect 20720 10192 20772 10198
rect 20718 10160 20720 10169
rect 20772 10160 20774 10169
rect 20718 10095 20774 10104
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19812 8650 19840 8774
rect 19996 8650 20024 9522
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 9178 20300 9318
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 19812 8622 20024 8650
rect 19890 7712 19946 7721
rect 19628 7528 19656 7686
rect 19720 7670 19890 7698
rect 19890 7647 19946 7656
rect 19628 7500 19840 7528
rect 19628 7342 19656 7500
rect 19706 7440 19762 7449
rect 19706 7375 19762 7384
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19614 7168 19670 7177
rect 19614 7103 19670 7112
rect 19628 6730 19656 7103
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19720 5681 19748 7375
rect 19812 6798 19840 7500
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19706 5672 19762 5681
rect 19706 5607 19762 5616
rect 19708 5024 19760 5030
rect 19536 4972 19708 4978
rect 19536 4966 19760 4972
rect 19536 4950 19748 4966
rect 19536 4078 19564 4950
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19522 3632 19578 3641
rect 19720 3602 19748 4422
rect 19812 4282 19840 4422
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19522 3567 19578 3576
rect 19708 3596 19760 3602
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19536 3058 19564 3567
rect 19708 3538 19760 3544
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19522 2952 19578 2961
rect 19432 2916 19484 2922
rect 19522 2887 19524 2896
rect 19432 2858 19484 2864
rect 19576 2887 19578 2896
rect 19524 2858 19576 2864
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19352 2650 19380 2790
rect 19444 2774 19472 2858
rect 19444 2746 19564 2774
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19536 2514 19564 2746
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 19812 2446 19840 3062
rect 19904 2922 19932 7647
rect 19996 6225 20024 8622
rect 20166 8528 20222 8537
rect 20166 8463 20222 8472
rect 20074 7848 20130 7857
rect 20074 7783 20130 7792
rect 19982 6216 20038 6225
rect 19982 6151 20038 6160
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19996 5914 20024 6054
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 20088 5710 20116 7783
rect 20180 6882 20208 8463
rect 20272 8294 20300 8842
rect 20364 8634 20392 9522
rect 20456 8906 20484 9862
rect 20543 9276 20851 9285
rect 20543 9274 20549 9276
rect 20605 9274 20629 9276
rect 20685 9274 20709 9276
rect 20765 9274 20789 9276
rect 20845 9274 20851 9276
rect 20605 9222 20607 9274
rect 20787 9222 20789 9274
rect 20543 9220 20549 9222
rect 20605 9220 20629 9222
rect 20685 9220 20709 9222
rect 20765 9220 20789 9222
rect 20845 9220 20851 9222
rect 20543 9211 20851 9220
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20272 7818 20300 8230
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20180 6854 20300 6882
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20180 6118 20208 6666
rect 20272 6361 20300 6854
rect 20258 6352 20314 6361
rect 20258 6287 20314 6296
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20180 5642 20208 6054
rect 20168 5636 20220 5642
rect 20168 5578 20220 5584
rect 20076 5568 20128 5574
rect 20074 5536 20076 5545
rect 20128 5536 20130 5545
rect 20074 5471 20130 5480
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20088 5273 20116 5306
rect 20074 5264 20130 5273
rect 19984 5228 20036 5234
rect 20074 5199 20130 5208
rect 19984 5170 20036 5176
rect 19996 4826 20024 5170
rect 20180 5166 20208 5578
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5370 20300 5510
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20168 5160 20220 5166
rect 20168 5102 20220 5108
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19996 3058 20024 3878
rect 20088 3738 20116 4558
rect 20180 4554 20208 5102
rect 20258 4584 20314 4593
rect 20168 4548 20220 4554
rect 20258 4519 20260 4528
rect 20168 4490 20220 4496
rect 20312 4519 20314 4528
rect 20260 4490 20312 4496
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20180 3534 20208 4490
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 3670 20300 3878
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 20180 2990 20208 3470
rect 20364 3194 20392 8570
rect 20548 8537 20576 8842
rect 20640 8838 20668 9114
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20534 8528 20590 8537
rect 20534 8463 20590 8472
rect 20456 8350 20668 8378
rect 20456 7721 20484 8350
rect 20640 8294 20668 8350
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20543 8188 20851 8197
rect 20543 8186 20549 8188
rect 20605 8186 20629 8188
rect 20685 8186 20709 8188
rect 20765 8186 20789 8188
rect 20845 8186 20851 8188
rect 20605 8134 20607 8186
rect 20787 8134 20789 8186
rect 20543 8132 20549 8134
rect 20605 8132 20629 8134
rect 20685 8132 20709 8134
rect 20765 8132 20789 8134
rect 20845 8132 20851 8134
rect 20543 8123 20851 8132
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20824 7721 20852 7754
rect 20442 7712 20498 7721
rect 20442 7647 20498 7656
rect 20810 7712 20866 7721
rect 20810 7647 20866 7656
rect 20543 7100 20851 7109
rect 20543 7098 20549 7100
rect 20605 7098 20629 7100
rect 20685 7098 20709 7100
rect 20765 7098 20789 7100
rect 20845 7098 20851 7100
rect 20605 7046 20607 7098
rect 20787 7046 20789 7098
rect 20543 7044 20549 7046
rect 20605 7044 20629 7046
rect 20685 7044 20709 7046
rect 20765 7044 20789 7046
rect 20845 7044 20851 7046
rect 20543 7035 20851 7044
rect 20536 6928 20588 6934
rect 20916 6882 20944 11047
rect 20994 9616 21050 9625
rect 20994 9551 21050 9560
rect 21008 9353 21036 9551
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20994 9344 21050 9353
rect 20994 9279 21050 9288
rect 21100 8974 21128 9454
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 21192 8498 21220 12815
rect 21270 12744 21326 12753
rect 21270 12679 21326 12688
rect 21284 11880 21312 12679
rect 21376 12306 21404 13790
rect 21468 13394 21496 13874
rect 21560 13802 21588 14758
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21560 13274 21588 13738
rect 21652 13530 21680 14350
rect 21744 13977 21772 14962
rect 21730 13968 21786 13977
rect 21730 13903 21786 13912
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21836 13394 21864 15302
rect 21928 15094 21956 15302
rect 22480 15162 22508 15846
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22020 14006 22048 14758
rect 22480 14482 22508 14758
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 21928 13870 21956 13942
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21560 13246 21680 13274
rect 21548 13184 21600 13190
rect 21468 13144 21548 13172
rect 21468 12442 21496 13144
rect 21548 13126 21600 13132
rect 21652 12850 21680 13246
rect 22020 12850 22048 13670
rect 21640 12844 21692 12850
rect 22008 12844 22060 12850
rect 21640 12786 21692 12792
rect 21928 12804 22008 12832
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21652 12322 21680 12786
rect 21928 12442 21956 12804
rect 22008 12786 22060 12792
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21560 12294 21680 12322
rect 21284 11852 21404 11880
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21284 11082 21312 11698
rect 21376 11150 21404 11852
rect 21560 11762 21588 12294
rect 22020 12238 22048 12582
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21652 11830 21680 12106
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21284 10470 21312 11018
rect 21560 10742 21588 11698
rect 21638 11656 21694 11665
rect 21638 11591 21694 11600
rect 21652 11558 21680 11591
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21744 11218 21772 12174
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 22020 11354 22048 12038
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22112 11234 22140 14350
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22204 12306 22232 13262
rect 22388 12986 22416 14214
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22296 11286 22324 11766
rect 22388 11694 22416 12242
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 22020 11206 22140 11234
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 21560 10470 21588 10678
rect 21744 10606 21772 11154
rect 21732 10600 21784 10606
rect 21732 10542 21784 10548
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21468 10062 21496 10406
rect 21914 10160 21970 10169
rect 21914 10095 21970 10104
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21284 9625 21312 9658
rect 21270 9616 21326 9625
rect 21270 9551 21326 9560
rect 21928 9518 21956 10095
rect 22020 9926 22048 11206
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22100 10736 22152 10742
rect 22098 10704 22100 10713
rect 22152 10704 22154 10713
rect 22098 10639 22154 10648
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 10062 22140 10406
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22296 9994 22324 10610
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 22388 9926 22416 10950
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22112 9654 22140 9862
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 21916 9512 21968 9518
rect 22284 9512 22336 9518
rect 21916 9454 21968 9460
rect 22204 9472 22284 9500
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21822 8936 21878 8945
rect 21822 8871 21824 8880
rect 21876 8871 21878 8880
rect 21824 8842 21876 8848
rect 21652 8622 22048 8650
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20536 6870 20588 6876
rect 20442 6488 20498 6497
rect 20442 6423 20498 6432
rect 20456 5846 20484 6423
rect 20548 6390 20576 6870
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20824 6854 20944 6882
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6497 20668 6598
rect 20626 6488 20682 6497
rect 20732 6458 20760 6802
rect 20824 6730 20852 6854
rect 20904 6792 20956 6798
rect 20902 6760 20904 6769
rect 20956 6760 20958 6769
rect 20812 6724 20864 6730
rect 20902 6695 20958 6704
rect 20812 6666 20864 6672
rect 20902 6624 20958 6633
rect 20902 6559 20958 6568
rect 20916 6458 20944 6559
rect 20626 6423 20682 6432
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20543 6012 20851 6021
rect 20543 6010 20549 6012
rect 20605 6010 20629 6012
rect 20685 6010 20709 6012
rect 20765 6010 20789 6012
rect 20845 6010 20851 6012
rect 20605 5958 20607 6010
rect 20787 5958 20789 6010
rect 20543 5956 20549 5958
rect 20605 5956 20629 5958
rect 20685 5956 20709 5958
rect 20765 5956 20789 5958
rect 20845 5956 20851 5958
rect 20543 5947 20851 5956
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20534 5400 20590 5409
rect 20534 5335 20590 5344
rect 20548 5302 20576 5335
rect 20536 5296 20588 5302
rect 20536 5238 20588 5244
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20456 4282 20484 4966
rect 20543 4924 20851 4933
rect 20543 4922 20549 4924
rect 20605 4922 20629 4924
rect 20685 4922 20709 4924
rect 20765 4922 20789 4924
rect 20845 4922 20851 4924
rect 20605 4870 20607 4922
rect 20787 4870 20789 4922
rect 20543 4868 20549 4870
rect 20605 4868 20629 4870
rect 20685 4868 20709 4870
rect 20765 4868 20789 4870
rect 20845 4868 20851 4870
rect 20543 4859 20851 4868
rect 20810 4720 20866 4729
rect 20810 4655 20866 4664
rect 20824 4622 20852 4655
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20548 4146 20576 4490
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20456 3720 20484 4014
rect 20543 3836 20851 3845
rect 20543 3834 20549 3836
rect 20605 3834 20629 3836
rect 20685 3834 20709 3836
rect 20765 3834 20789 3836
rect 20845 3834 20851 3836
rect 20605 3782 20607 3834
rect 20787 3782 20789 3834
rect 20543 3780 20549 3782
rect 20605 3780 20629 3782
rect 20685 3780 20709 3782
rect 20765 3780 20789 3782
rect 20845 3780 20851 3782
rect 20543 3771 20851 3780
rect 20456 3692 20576 3720
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20456 3194 20484 3334
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20364 3074 20392 3130
rect 20364 3046 20484 3074
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19996 2650 20024 2790
rect 20180 2650 20208 2926
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 20364 2378 20392 2790
rect 20456 2650 20484 3046
rect 20548 2922 20576 3692
rect 20916 3534 20944 5850
rect 21008 5370 21036 8026
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21100 6866 21128 7958
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 21100 3602 21128 6598
rect 21192 6458 21220 7890
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21180 5720 21232 5726
rect 21180 5662 21232 5668
rect 21192 5409 21220 5662
rect 21178 5400 21234 5409
rect 21178 5335 21234 5344
rect 21178 5128 21234 5137
rect 21178 5063 21234 5072
rect 21192 4622 21220 5063
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 20543 2748 20851 2757
rect 20543 2746 20549 2748
rect 20605 2746 20629 2748
rect 20685 2746 20709 2748
rect 20765 2746 20789 2748
rect 20845 2746 20851 2748
rect 20605 2694 20607 2746
rect 20787 2694 20789 2746
rect 20543 2692 20549 2694
rect 20605 2692 20629 2694
rect 20685 2692 20709 2694
rect 20765 2692 20789 2694
rect 20845 2692 20851 2694
rect 20543 2683 20851 2692
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20916 2446 20944 2994
rect 21100 2854 21128 3402
rect 21192 3058 21220 4558
rect 21284 4146 21312 8298
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21376 7018 21404 7822
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21468 7449 21496 7482
rect 21454 7440 21510 7449
rect 21454 7375 21510 7384
rect 21456 7200 21508 7206
rect 21454 7168 21456 7177
rect 21560 7188 21588 8434
rect 21652 7546 21680 8622
rect 22020 8498 22048 8622
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22112 8378 22140 9114
rect 21836 8362 22140 8378
rect 21824 8356 22140 8362
rect 21876 8350 22140 8356
rect 21824 8298 21876 8304
rect 22112 8294 22140 8350
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 21822 7984 21878 7993
rect 21732 7948 21784 7954
rect 21822 7919 21878 7928
rect 22006 7984 22062 7993
rect 22006 7919 22062 7928
rect 21732 7890 21784 7896
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21508 7168 21588 7188
rect 21510 7160 21588 7168
rect 21454 7103 21510 7112
rect 21376 6990 21496 7018
rect 21468 6644 21496 6990
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21548 6656 21600 6662
rect 21468 6616 21548 6644
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21376 5370 21404 6190
rect 21468 5574 21496 6616
rect 21548 6598 21600 6604
rect 21546 6352 21602 6361
rect 21546 6287 21602 6296
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21560 5234 21588 6287
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21652 4826 21680 6802
rect 21744 6186 21772 7890
rect 21836 7342 21864 7919
rect 22020 7750 22048 7919
rect 22098 7848 22154 7857
rect 22098 7783 22154 7792
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21822 6624 21878 6633
rect 21822 6559 21878 6568
rect 21836 6254 21864 6559
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21744 5914 21772 6122
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21730 5808 21786 5817
rect 21730 5743 21786 5752
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21270 4040 21326 4049
rect 21376 4010 21404 4082
rect 21270 3975 21326 3984
rect 21364 4004 21416 4010
rect 21284 3398 21312 3975
rect 21364 3946 21416 3952
rect 21376 3738 21404 3946
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 21560 3641 21588 3878
rect 21546 3632 21602 3641
rect 21546 3567 21602 3576
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 21744 2961 21772 5743
rect 21836 4690 21864 6054
rect 21914 5944 21970 5953
rect 21914 5879 21970 5888
rect 21928 5778 21956 5879
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21730 2952 21786 2961
rect 21730 2887 21786 2896
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 22020 2446 22048 7686
rect 22112 7546 22140 7783
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22112 6089 22140 7210
rect 22204 6633 22232 9472
rect 22284 9454 22336 9460
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22296 7546 22324 8366
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22296 7041 22324 7346
rect 22388 7206 22416 7822
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22282 7032 22338 7041
rect 22282 6967 22338 6976
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22190 6624 22246 6633
rect 22190 6559 22246 6568
rect 22296 6474 22324 6802
rect 22204 6446 22324 6474
rect 22204 6390 22232 6446
rect 22192 6384 22244 6390
rect 22284 6384 22336 6390
rect 22192 6326 22244 6332
rect 22282 6352 22284 6361
rect 22336 6352 22338 6361
rect 22282 6287 22338 6296
rect 22190 6216 22246 6225
rect 22190 6151 22246 6160
rect 22098 6080 22154 6089
rect 22098 6015 22154 6024
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22112 4690 22140 5850
rect 22204 5302 22232 6151
rect 22296 5370 22324 6287
rect 22388 6254 22416 6938
rect 22480 6361 22508 14282
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22572 13394 22600 13670
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22664 12374 22692 16390
rect 22756 15502 22784 16934
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22756 15162 22784 15302
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 22756 12238 22784 14486
rect 22848 14074 22876 19314
rect 22940 17066 22968 20402
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23124 19961 23152 20266
rect 23110 19952 23166 19961
rect 23110 19887 23166 19896
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 18873 23060 19654
rect 23112 19304 23164 19310
rect 23110 19272 23112 19281
rect 23164 19272 23166 19281
rect 23110 19207 23166 19216
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23018 18864 23074 18873
rect 23018 18799 23074 18808
rect 23020 18760 23072 18766
rect 23020 18702 23072 18708
rect 23032 17338 23060 18702
rect 23124 18329 23152 19110
rect 23216 18601 23244 21966
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23308 19417 23336 20198
rect 23294 19408 23350 19417
rect 23294 19343 23350 19352
rect 23202 18592 23258 18601
rect 23202 18527 23258 18536
rect 23110 18320 23166 18329
rect 23110 18255 23166 18264
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 22928 17060 22980 17066
rect 22928 17002 22980 17008
rect 23032 16794 23060 17274
rect 23124 17241 23152 17478
rect 23110 17232 23166 17241
rect 23110 17167 23166 17176
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23216 16182 23244 17818
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22940 15978 22968 16050
rect 22928 15972 22980 15978
rect 22928 15914 22980 15920
rect 22940 15065 22968 15914
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22926 15056 22982 15065
rect 22926 14991 22982 15000
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23032 14414 23060 14758
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22940 13394 22968 14214
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 23124 12850 23152 15846
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23216 14521 23244 14962
rect 23202 14512 23258 14521
rect 23202 14447 23258 14456
rect 23308 14396 23336 17138
rect 23216 14368 23336 14396
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22940 12434 22968 12582
rect 23216 12434 23244 14368
rect 22940 12406 23060 12434
rect 23216 12406 23336 12434
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22744 12232 22796 12238
rect 22650 12200 22706 12209
rect 22744 12174 22796 12180
rect 22650 12135 22706 12144
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22572 11642 22600 12038
rect 22664 11830 22692 12135
rect 22744 12096 22796 12102
rect 22742 12064 22744 12073
rect 22796 12064 22798 12073
rect 22742 11999 22798 12008
rect 22834 11928 22890 11937
rect 22834 11863 22890 11872
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 22572 11614 22692 11642
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22572 10810 22600 11494
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22664 10062 22692 11614
rect 22848 11218 22876 11863
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22834 10024 22890 10033
rect 22834 9959 22890 9968
rect 22848 9654 22876 9959
rect 22836 9648 22888 9654
rect 22742 9616 22798 9625
rect 22836 9590 22888 9596
rect 22742 9551 22798 9560
rect 22558 9480 22614 9489
rect 22558 9415 22614 9424
rect 22572 8906 22600 9415
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22664 9042 22692 9318
rect 22756 9042 22784 9551
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22834 7576 22890 7585
rect 22834 7511 22890 7520
rect 22848 7478 22876 7511
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 22940 7410 22968 12310
rect 23032 12306 23060 12406
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 11218 23060 12242
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 23308 10146 23336 12406
rect 23400 10742 23428 21830
rect 23492 20058 23520 23800
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23584 15473 23612 20334
rect 23676 16017 23704 20878
rect 24136 19446 24164 23800
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 23662 16008 23718 16017
rect 23662 15943 23718 15952
rect 23570 15464 23626 15473
rect 23570 15399 23626 15408
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23308 10118 23796 10146
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23032 8974 23060 9318
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23032 8838 23060 8910
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22742 7304 22798 7313
rect 22652 7268 22704 7274
rect 22742 7239 22798 7248
rect 22652 7210 22704 7216
rect 22664 6905 22692 7210
rect 22650 6896 22706 6905
rect 22650 6831 22706 6840
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22466 6352 22522 6361
rect 22466 6287 22522 6296
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 22374 6080 22430 6089
rect 22374 6015 22430 6024
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22112 4282 22140 4422
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22112 2514 22140 4082
rect 22296 3602 22324 4558
rect 22388 3738 22416 6015
rect 22468 5772 22520 5778
rect 22572 5760 22600 6734
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22520 5732 22600 5760
rect 22468 5714 22520 5720
rect 22558 5672 22614 5681
rect 22558 5607 22614 5616
rect 22572 5574 22600 5607
rect 22560 5568 22612 5574
rect 22466 5536 22522 5545
rect 22560 5510 22612 5516
rect 22466 5471 22522 5480
rect 22480 4026 22508 5471
rect 22664 5409 22692 6598
rect 22650 5400 22706 5409
rect 22650 5335 22652 5344
rect 22704 5335 22706 5344
rect 22652 5306 22704 5312
rect 22650 5264 22706 5273
rect 22560 5228 22612 5234
rect 22650 5199 22706 5208
rect 22560 5170 22612 5176
rect 22572 4185 22600 5170
rect 22664 4690 22692 5199
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22558 4176 22614 4185
rect 22558 4111 22614 4120
rect 22756 4078 22784 7239
rect 23032 7206 23060 8774
rect 23110 8528 23166 8537
rect 23110 8463 23112 8472
rect 23164 8463 23166 8472
rect 23112 8434 23164 8440
rect 23112 7744 23164 7750
rect 23112 7686 23164 7692
rect 22836 7200 22888 7206
rect 23020 7200 23072 7206
rect 22888 7148 22968 7154
rect 22836 7142 22968 7148
rect 23020 7142 23072 7148
rect 22848 7126 22968 7142
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 22848 5817 22876 6122
rect 22834 5808 22890 5817
rect 22834 5743 22890 5752
rect 22848 5710 22876 5743
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22940 5522 22968 7126
rect 23032 6458 23060 7142
rect 23124 7002 23152 7686
rect 23112 6996 23164 7002
rect 23112 6938 23164 6944
rect 23110 6896 23166 6905
rect 23110 6831 23166 6840
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23018 6352 23074 6361
rect 23018 6287 23074 6296
rect 23032 5914 23060 6287
rect 23124 6186 23152 6831
rect 23112 6180 23164 6186
rect 23112 6122 23164 6128
rect 23020 5908 23072 5914
rect 23216 5896 23244 9046
rect 23294 8664 23350 8673
rect 23294 8599 23350 8608
rect 23308 6322 23336 8599
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23020 5850 23072 5856
rect 23124 5868 23244 5896
rect 23124 5545 23152 5868
rect 23202 5808 23258 5817
rect 23202 5743 23258 5752
rect 22848 5494 22968 5522
rect 23110 5536 23166 5545
rect 22744 4072 22796 4078
rect 22480 3998 22600 4026
rect 22744 4014 22796 4020
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22480 3466 22508 3878
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22204 2446 22232 2926
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 22192 2304 22244 2310
rect 22296 2258 22324 3402
rect 22572 3398 22600 3998
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22560 3392 22612 3398
rect 22466 3360 22522 3369
rect 22560 3334 22612 3340
rect 22466 3295 22522 3304
rect 22480 2582 22508 3295
rect 22664 3058 22692 3878
rect 22742 3768 22798 3777
rect 22742 3703 22798 3712
rect 22756 3534 22784 3703
rect 22848 3670 22876 5494
rect 23110 5471 23166 5480
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22940 5273 22968 5306
rect 22926 5264 22982 5273
rect 22926 5199 22982 5208
rect 23018 4720 23074 4729
rect 23018 4655 23074 4664
rect 23032 3738 23060 4655
rect 23110 4176 23166 4185
rect 23110 4111 23166 4120
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 22836 3664 22888 3670
rect 22836 3606 22888 3612
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 23124 3194 23152 4111
rect 23216 4010 23244 5743
rect 23308 4758 23336 6258
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23400 4622 23428 6802
rect 23492 6390 23520 9862
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23662 8392 23718 8401
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23584 4146 23612 8366
rect 23662 8327 23718 8336
rect 23676 5778 23704 8327
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23768 4078 23796 10118
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23204 4004 23256 4010
rect 23204 3946 23256 3952
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23018 3088 23074 3097
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22744 3052 22796 3058
rect 23018 3023 23074 3032
rect 22744 2994 22796 3000
rect 22664 2650 22692 2994
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22468 2576 22520 2582
rect 22468 2518 22520 2524
rect 22650 2544 22706 2553
rect 22480 2446 22508 2518
rect 22756 2514 22784 2994
rect 23032 2650 23060 3023
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23860 2582 23888 13806
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 22650 2479 22706 2488
rect 22744 2508 22796 2514
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22664 2310 22692 2479
rect 22744 2450 22796 2456
rect 22244 2252 22324 2258
rect 22192 2246 22324 2252
rect 22376 2304 22428 2310
rect 22376 2246 22428 2252
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 6548 2204 6856 2213
rect 6548 2202 6554 2204
rect 6610 2202 6634 2204
rect 6690 2202 6714 2204
rect 6770 2202 6794 2204
rect 6850 2202 6856 2204
rect 6610 2150 6612 2202
rect 6792 2150 6794 2202
rect 6548 2148 6554 2150
rect 6610 2148 6634 2150
rect 6690 2148 6714 2150
rect 6770 2148 6794 2150
rect 6850 2148 6856 2150
rect 6548 2139 6856 2148
rect 10244 800 10272 2246
rect 22204 2230 22324 2246
rect 12146 2204 12454 2213
rect 12146 2202 12152 2204
rect 12208 2202 12232 2204
rect 12288 2202 12312 2204
rect 12368 2202 12392 2204
rect 12448 2202 12454 2204
rect 12208 2150 12210 2202
rect 12390 2150 12392 2202
rect 12146 2148 12152 2150
rect 12208 2148 12232 2150
rect 12288 2148 12312 2150
rect 12368 2148 12392 2150
rect 12448 2148 12454 2150
rect 12146 2139 12454 2148
rect 17744 2204 18052 2213
rect 17744 2202 17750 2204
rect 17806 2202 17830 2204
rect 17886 2202 17910 2204
rect 17966 2202 17990 2204
rect 18046 2202 18052 2204
rect 17806 2150 17808 2202
rect 17988 2150 17990 2202
rect 17744 2148 17750 2150
rect 17806 2148 17830 2150
rect 17886 2148 17910 2150
rect 17966 2148 17990 2150
rect 18046 2148 18052 2150
rect 17744 2139 18052 2148
rect 22388 800 22416 2246
rect 2134 0 2190 800
rect 6182 0 6238 800
rect 10230 0 10286 800
rect 14278 0 14334 800
rect 18326 0 18382 800
rect 22374 0 22430 800
<< via2 >>
rect 2318 21664 2374 21720
rect 2042 20884 2044 20904
rect 2044 20884 2096 20904
rect 2096 20884 2098 20904
rect 2042 20848 2098 20884
rect 3330 22480 3386 22536
rect 2962 22072 3018 22128
rect 2778 21800 2834 21856
rect 2686 20848 2742 20904
rect 3054 21664 3110 21720
rect 3755 22330 3811 22332
rect 3835 22330 3891 22332
rect 3915 22330 3971 22332
rect 3995 22330 4051 22332
rect 3755 22278 3801 22330
rect 3801 22278 3811 22330
rect 3835 22278 3865 22330
rect 3865 22278 3877 22330
rect 3877 22278 3891 22330
rect 3915 22278 3929 22330
rect 3929 22278 3941 22330
rect 3941 22278 3971 22330
rect 3995 22278 4005 22330
rect 4005 22278 4051 22330
rect 3755 22276 3811 22278
rect 3835 22276 3891 22278
rect 3915 22276 3971 22278
rect 3995 22276 4051 22278
rect 3606 21972 3608 21992
rect 3608 21972 3660 21992
rect 3660 21972 3662 21992
rect 3606 21936 3662 21972
rect 3790 22072 3846 22128
rect 4434 22208 4490 22264
rect 3422 21392 3478 21448
rect 3422 20984 3478 21040
rect 3146 20576 3202 20632
rect 3238 20440 3294 20496
rect 2778 18264 2834 18320
rect 3755 21242 3811 21244
rect 3835 21242 3891 21244
rect 3915 21242 3971 21244
rect 3995 21242 4051 21244
rect 3755 21190 3801 21242
rect 3801 21190 3811 21242
rect 3835 21190 3865 21242
rect 3865 21190 3877 21242
rect 3877 21190 3891 21242
rect 3915 21190 3929 21242
rect 3929 21190 3941 21242
rect 3941 21190 3971 21242
rect 3995 21190 4005 21242
rect 4005 21190 4051 21242
rect 3755 21188 3811 21190
rect 3835 21188 3891 21190
rect 3915 21188 3971 21190
rect 3995 21188 4051 21190
rect 4526 21800 4582 21856
rect 4526 21256 4582 21312
rect 4250 20848 4306 20904
rect 3755 20154 3811 20156
rect 3835 20154 3891 20156
rect 3915 20154 3971 20156
rect 3995 20154 4051 20156
rect 3755 20102 3801 20154
rect 3801 20102 3811 20154
rect 3835 20102 3865 20154
rect 3865 20102 3877 20154
rect 3877 20102 3891 20154
rect 3915 20102 3929 20154
rect 3929 20102 3941 20154
rect 3941 20102 3971 20154
rect 3995 20102 4005 20154
rect 4005 20102 4051 20154
rect 3755 20100 3811 20102
rect 3835 20100 3891 20102
rect 3915 20100 3971 20102
rect 3995 20100 4051 20102
rect 3755 19066 3811 19068
rect 3835 19066 3891 19068
rect 3915 19066 3971 19068
rect 3995 19066 4051 19068
rect 3755 19014 3801 19066
rect 3801 19014 3811 19066
rect 3835 19014 3865 19066
rect 3865 19014 3877 19066
rect 3877 19014 3891 19066
rect 3915 19014 3929 19066
rect 3929 19014 3941 19066
rect 3941 19014 3971 19066
rect 3995 19014 4005 19066
rect 4005 19014 4051 19066
rect 3755 19012 3811 19014
rect 3835 19012 3891 19014
rect 3915 19012 3971 19014
rect 3995 19012 4051 19014
rect 3514 18672 3570 18728
rect 3882 18536 3938 18592
rect 3422 18400 3478 18456
rect 1490 15308 1492 15328
rect 1492 15308 1544 15328
rect 1544 15308 1546 15328
rect 1490 15272 1546 15308
rect 1398 9152 1454 9208
rect 4158 17992 4214 18048
rect 3755 17978 3811 17980
rect 3835 17978 3891 17980
rect 3915 17978 3971 17980
rect 3995 17978 4051 17980
rect 3755 17926 3801 17978
rect 3801 17926 3811 17978
rect 3835 17926 3865 17978
rect 3865 17926 3877 17978
rect 3877 17926 3891 17978
rect 3915 17926 3929 17978
rect 3929 17926 3941 17978
rect 3941 17926 3971 17978
rect 3995 17926 4005 17978
rect 4005 17926 4051 17978
rect 3755 17924 3811 17926
rect 3835 17924 3891 17926
rect 3915 17924 3971 17926
rect 3995 17924 4051 17926
rect 4066 17584 4122 17640
rect 3755 16890 3811 16892
rect 3835 16890 3891 16892
rect 3915 16890 3971 16892
rect 3995 16890 4051 16892
rect 3755 16838 3801 16890
rect 3801 16838 3811 16890
rect 3835 16838 3865 16890
rect 3865 16838 3877 16890
rect 3877 16838 3891 16890
rect 3915 16838 3929 16890
rect 3929 16838 3941 16890
rect 3941 16838 3971 16890
rect 3995 16838 4005 16890
rect 4005 16838 4051 16890
rect 3755 16836 3811 16838
rect 3835 16836 3891 16838
rect 3915 16836 3971 16838
rect 3995 16836 4051 16838
rect 3755 15802 3811 15804
rect 3835 15802 3891 15804
rect 3915 15802 3971 15804
rect 3995 15802 4051 15804
rect 3755 15750 3801 15802
rect 3801 15750 3811 15802
rect 3835 15750 3865 15802
rect 3865 15750 3877 15802
rect 3877 15750 3891 15802
rect 3915 15750 3929 15802
rect 3929 15750 3941 15802
rect 3941 15750 3971 15802
rect 3995 15750 4005 15802
rect 4005 15750 4051 15802
rect 3755 15748 3811 15750
rect 3835 15748 3891 15750
rect 3915 15748 3971 15750
rect 3995 15748 4051 15750
rect 5354 22344 5410 22400
rect 4802 20576 4858 20632
rect 4986 20576 5042 20632
rect 4986 18128 5042 18184
rect 5170 18536 5226 18592
rect 7194 22208 7250 22264
rect 6182 21836 6184 21856
rect 6184 21836 6236 21856
rect 6236 21836 6238 21856
rect 6182 21800 6238 21836
rect 6550 21936 6606 21992
rect 6734 21972 6736 21992
rect 6736 21972 6788 21992
rect 6788 21972 6790 21992
rect 6734 21936 6790 21972
rect 6366 21664 6422 21720
rect 6090 21120 6146 21176
rect 5446 18808 5502 18864
rect 5722 19896 5778 19952
rect 5630 18808 5686 18864
rect 5262 18400 5318 18456
rect 5170 17992 5226 18048
rect 4250 15272 4306 15328
rect 3755 14714 3811 14716
rect 3835 14714 3891 14716
rect 3915 14714 3971 14716
rect 3995 14714 4051 14716
rect 3755 14662 3801 14714
rect 3801 14662 3811 14714
rect 3835 14662 3865 14714
rect 3865 14662 3877 14714
rect 3877 14662 3891 14714
rect 3915 14662 3929 14714
rect 3929 14662 3941 14714
rect 3941 14662 3971 14714
rect 3995 14662 4005 14714
rect 4005 14662 4051 14714
rect 3755 14660 3811 14662
rect 3835 14660 3891 14662
rect 3915 14660 3971 14662
rect 3995 14660 4051 14662
rect 3755 13626 3811 13628
rect 3835 13626 3891 13628
rect 3915 13626 3971 13628
rect 3995 13626 4051 13628
rect 3755 13574 3801 13626
rect 3801 13574 3811 13626
rect 3835 13574 3865 13626
rect 3865 13574 3877 13626
rect 3877 13574 3891 13626
rect 3915 13574 3929 13626
rect 3929 13574 3941 13626
rect 3941 13574 3971 13626
rect 3995 13574 4005 13626
rect 4005 13574 4051 13626
rect 3755 13572 3811 13574
rect 3835 13572 3891 13574
rect 3915 13572 3971 13574
rect 3995 13572 4051 13574
rect 4158 12824 4214 12880
rect 3755 12538 3811 12540
rect 3835 12538 3891 12540
rect 3915 12538 3971 12540
rect 3995 12538 4051 12540
rect 3755 12486 3801 12538
rect 3801 12486 3811 12538
rect 3835 12486 3865 12538
rect 3865 12486 3877 12538
rect 3877 12486 3891 12538
rect 3915 12486 3929 12538
rect 3929 12486 3941 12538
rect 3941 12486 3971 12538
rect 3995 12486 4005 12538
rect 4005 12486 4051 12538
rect 3755 12484 3811 12486
rect 3835 12484 3891 12486
rect 3915 12484 3971 12486
rect 3995 12484 4051 12486
rect 3882 11736 3938 11792
rect 3755 11450 3811 11452
rect 3835 11450 3891 11452
rect 3915 11450 3971 11452
rect 3995 11450 4051 11452
rect 3755 11398 3801 11450
rect 3801 11398 3811 11450
rect 3835 11398 3865 11450
rect 3865 11398 3877 11450
rect 3877 11398 3891 11450
rect 3915 11398 3929 11450
rect 3929 11398 3941 11450
rect 3941 11398 3971 11450
rect 3995 11398 4005 11450
rect 4005 11398 4051 11450
rect 3755 11396 3811 11398
rect 3835 11396 3891 11398
rect 3915 11396 3971 11398
rect 3995 11396 4051 11398
rect 3755 10362 3811 10364
rect 3835 10362 3891 10364
rect 3915 10362 3971 10364
rect 3995 10362 4051 10364
rect 3755 10310 3801 10362
rect 3801 10310 3811 10362
rect 3835 10310 3865 10362
rect 3865 10310 3877 10362
rect 3877 10310 3891 10362
rect 3915 10310 3929 10362
rect 3929 10310 3941 10362
rect 3941 10310 3971 10362
rect 3995 10310 4005 10362
rect 4005 10310 4051 10362
rect 3755 10308 3811 10310
rect 3835 10308 3891 10310
rect 3915 10308 3971 10310
rect 3995 10308 4051 10310
rect 4894 15020 4950 15056
rect 4894 15000 4896 15020
rect 4896 15000 4948 15020
rect 4948 15000 4950 15020
rect 6090 20712 6146 20768
rect 7010 21800 7066 21856
rect 6554 21786 6610 21788
rect 6634 21786 6690 21788
rect 6714 21786 6770 21788
rect 6794 21786 6850 21788
rect 6554 21734 6600 21786
rect 6600 21734 6610 21786
rect 6634 21734 6664 21786
rect 6664 21734 6676 21786
rect 6676 21734 6690 21786
rect 6714 21734 6728 21786
rect 6728 21734 6740 21786
rect 6740 21734 6770 21786
rect 6794 21734 6804 21786
rect 6804 21734 6850 21786
rect 6554 21732 6610 21734
rect 6634 21732 6690 21734
rect 6714 21732 6770 21734
rect 6794 21732 6850 21734
rect 6274 20576 6330 20632
rect 7102 21664 7158 21720
rect 7102 21256 7158 21312
rect 6642 20848 6698 20904
rect 6826 20884 6828 20904
rect 6828 20884 6880 20904
rect 6880 20884 6882 20904
rect 6826 20848 6882 20884
rect 8758 22344 8814 22400
rect 9353 22330 9409 22332
rect 9433 22330 9489 22332
rect 9513 22330 9569 22332
rect 9593 22330 9649 22332
rect 9353 22278 9399 22330
rect 9399 22278 9409 22330
rect 9433 22278 9463 22330
rect 9463 22278 9475 22330
rect 9475 22278 9489 22330
rect 9513 22278 9527 22330
rect 9527 22278 9539 22330
rect 9539 22278 9569 22330
rect 9593 22278 9603 22330
rect 9603 22278 9649 22330
rect 9353 22276 9409 22278
rect 9433 22276 9489 22278
rect 9513 22276 9569 22278
rect 9593 22276 9649 22278
rect 8574 21836 8576 21856
rect 8576 21836 8628 21856
rect 8628 21836 8630 21856
rect 6554 20698 6610 20700
rect 6634 20698 6690 20700
rect 6714 20698 6770 20700
rect 6794 20698 6850 20700
rect 6554 20646 6600 20698
rect 6600 20646 6610 20698
rect 6634 20646 6664 20698
rect 6664 20646 6676 20698
rect 6676 20646 6690 20698
rect 6714 20646 6728 20698
rect 6728 20646 6740 20698
rect 6740 20646 6770 20698
rect 6794 20646 6804 20698
rect 6804 20646 6850 20698
rect 6554 20644 6610 20646
rect 6634 20644 6690 20646
rect 6714 20644 6770 20646
rect 6794 20644 6850 20646
rect 6554 19610 6610 19612
rect 6634 19610 6690 19612
rect 6714 19610 6770 19612
rect 6794 19610 6850 19612
rect 6554 19558 6600 19610
rect 6600 19558 6610 19610
rect 6634 19558 6664 19610
rect 6664 19558 6676 19610
rect 6676 19558 6690 19610
rect 6714 19558 6728 19610
rect 6728 19558 6740 19610
rect 6740 19558 6770 19610
rect 6794 19558 6804 19610
rect 6804 19558 6850 19610
rect 6554 19556 6610 19558
rect 6634 19556 6690 19558
rect 6714 19556 6770 19558
rect 6794 19556 6850 19558
rect 6090 18672 6146 18728
rect 6554 18522 6610 18524
rect 6634 18522 6690 18524
rect 6714 18522 6770 18524
rect 6794 18522 6850 18524
rect 6554 18470 6600 18522
rect 6600 18470 6610 18522
rect 6634 18470 6664 18522
rect 6664 18470 6676 18522
rect 6676 18470 6690 18522
rect 6714 18470 6728 18522
rect 6728 18470 6740 18522
rect 6740 18470 6770 18522
rect 6794 18470 6804 18522
rect 6804 18470 6850 18522
rect 6554 18468 6610 18470
rect 6634 18468 6690 18470
rect 6714 18468 6770 18470
rect 6794 18468 6850 18470
rect 6458 17992 6514 18048
rect 7286 20304 7342 20360
rect 6918 17720 6974 17776
rect 6554 17434 6610 17436
rect 6634 17434 6690 17436
rect 6714 17434 6770 17436
rect 6794 17434 6850 17436
rect 6554 17382 6600 17434
rect 6600 17382 6610 17434
rect 6634 17382 6664 17434
rect 6664 17382 6676 17434
rect 6676 17382 6690 17434
rect 6714 17382 6728 17434
rect 6728 17382 6740 17434
rect 6740 17382 6770 17434
rect 6794 17382 6804 17434
rect 6804 17382 6850 17434
rect 6554 17380 6610 17382
rect 6634 17380 6690 17382
rect 6714 17380 6770 17382
rect 6794 17380 6850 17382
rect 6554 16346 6610 16348
rect 6634 16346 6690 16348
rect 6714 16346 6770 16348
rect 6794 16346 6850 16348
rect 6554 16294 6600 16346
rect 6600 16294 6610 16346
rect 6634 16294 6664 16346
rect 6664 16294 6676 16346
rect 6676 16294 6690 16346
rect 6714 16294 6728 16346
rect 6728 16294 6740 16346
rect 6740 16294 6770 16346
rect 6794 16294 6804 16346
rect 6804 16294 6850 16346
rect 6554 16292 6610 16294
rect 6634 16292 6690 16294
rect 6714 16292 6770 16294
rect 6794 16292 6850 16294
rect 6554 15258 6610 15260
rect 6634 15258 6690 15260
rect 6714 15258 6770 15260
rect 6794 15258 6850 15260
rect 6554 15206 6600 15258
rect 6600 15206 6610 15258
rect 6634 15206 6664 15258
rect 6664 15206 6676 15258
rect 6676 15206 6690 15258
rect 6714 15206 6728 15258
rect 6728 15206 6740 15258
rect 6740 15206 6770 15258
rect 6794 15206 6804 15258
rect 6804 15206 6850 15258
rect 6554 15204 6610 15206
rect 6634 15204 6690 15206
rect 6714 15204 6770 15206
rect 6794 15204 6850 15206
rect 5354 13388 5410 13424
rect 5354 13368 5356 13388
rect 5356 13368 5408 13388
rect 5408 13368 5410 13388
rect 7194 18264 7250 18320
rect 7470 17584 7526 17640
rect 8574 21800 8630 21836
rect 8758 21800 8814 21856
rect 8758 21120 8814 21176
rect 10230 22208 10286 22264
rect 9862 21936 9918 21992
rect 10046 21936 10102 21992
rect 9402 21800 9458 21856
rect 9126 21392 9182 21448
rect 10046 21528 10102 21584
rect 9126 21120 9182 21176
rect 9353 21242 9409 21244
rect 9433 21242 9489 21244
rect 9513 21242 9569 21244
rect 9593 21242 9649 21244
rect 9353 21190 9399 21242
rect 9399 21190 9409 21242
rect 9433 21190 9463 21242
rect 9463 21190 9475 21242
rect 9475 21190 9489 21242
rect 9513 21190 9527 21242
rect 9527 21190 9539 21242
rect 9539 21190 9569 21242
rect 9593 21190 9603 21242
rect 9603 21190 9649 21242
rect 9353 21188 9409 21190
rect 9433 21188 9489 21190
rect 9513 21188 9569 21190
rect 9593 21188 9649 21190
rect 8666 18128 8722 18184
rect 9770 21256 9826 21312
rect 10138 20848 10194 20904
rect 9353 20154 9409 20156
rect 9433 20154 9489 20156
rect 9513 20154 9569 20156
rect 9593 20154 9649 20156
rect 9353 20102 9399 20154
rect 9399 20102 9409 20154
rect 9433 20102 9463 20154
rect 9463 20102 9475 20154
rect 9475 20102 9489 20154
rect 9513 20102 9527 20154
rect 9527 20102 9539 20154
rect 9539 20102 9569 20154
rect 9593 20102 9603 20154
rect 9603 20102 9649 20154
rect 9353 20100 9409 20102
rect 9433 20100 9489 20102
rect 9513 20100 9569 20102
rect 9593 20100 9649 20102
rect 9353 19066 9409 19068
rect 9433 19066 9489 19068
rect 9513 19066 9569 19068
rect 9593 19066 9649 19068
rect 9353 19014 9399 19066
rect 9399 19014 9409 19066
rect 9433 19014 9463 19066
rect 9463 19014 9475 19066
rect 9475 19014 9489 19066
rect 9513 19014 9527 19066
rect 9527 19014 9539 19066
rect 9539 19014 9569 19066
rect 9593 19014 9603 19066
rect 9603 19014 9649 19066
rect 9353 19012 9409 19014
rect 9433 19012 9489 19014
rect 9513 19012 9569 19014
rect 9593 19012 9649 19014
rect 9353 17978 9409 17980
rect 9433 17978 9489 17980
rect 9513 17978 9569 17980
rect 9593 17978 9649 17980
rect 9353 17926 9399 17978
rect 9399 17926 9409 17978
rect 9433 17926 9463 17978
rect 9463 17926 9475 17978
rect 9475 17926 9489 17978
rect 9513 17926 9527 17978
rect 9527 17926 9539 17978
rect 9539 17926 9569 17978
rect 9593 17926 9603 17978
rect 9603 17926 9649 17978
rect 9353 17924 9409 17926
rect 9433 17924 9489 17926
rect 9513 17924 9569 17926
rect 9593 17924 9649 17926
rect 9353 16890 9409 16892
rect 9433 16890 9489 16892
rect 9513 16890 9569 16892
rect 9593 16890 9649 16892
rect 9353 16838 9399 16890
rect 9399 16838 9409 16890
rect 9433 16838 9463 16890
rect 9463 16838 9475 16890
rect 9475 16838 9489 16890
rect 9513 16838 9527 16890
rect 9527 16838 9539 16890
rect 9539 16838 9569 16890
rect 9593 16838 9603 16890
rect 9603 16838 9649 16890
rect 9353 16836 9409 16838
rect 9433 16836 9489 16838
rect 9513 16836 9569 16838
rect 9593 16836 9649 16838
rect 6554 14170 6610 14172
rect 6634 14170 6690 14172
rect 6714 14170 6770 14172
rect 6794 14170 6850 14172
rect 6554 14118 6600 14170
rect 6600 14118 6610 14170
rect 6634 14118 6664 14170
rect 6664 14118 6676 14170
rect 6676 14118 6690 14170
rect 6714 14118 6728 14170
rect 6728 14118 6740 14170
rect 6740 14118 6770 14170
rect 6794 14118 6804 14170
rect 6804 14118 6850 14170
rect 6554 14116 6610 14118
rect 6634 14116 6690 14118
rect 6714 14116 6770 14118
rect 6794 14116 6850 14118
rect 6554 13082 6610 13084
rect 6634 13082 6690 13084
rect 6714 13082 6770 13084
rect 6794 13082 6850 13084
rect 6554 13030 6600 13082
rect 6600 13030 6610 13082
rect 6634 13030 6664 13082
rect 6664 13030 6676 13082
rect 6676 13030 6690 13082
rect 6714 13030 6728 13082
rect 6728 13030 6740 13082
rect 6740 13030 6770 13082
rect 6794 13030 6804 13082
rect 6804 13030 6850 13082
rect 6554 13028 6610 13030
rect 6634 13028 6690 13030
rect 6714 13028 6770 13030
rect 6794 13028 6850 13030
rect 6554 11994 6610 11996
rect 6634 11994 6690 11996
rect 6714 11994 6770 11996
rect 6794 11994 6850 11996
rect 6554 11942 6600 11994
rect 6600 11942 6610 11994
rect 6634 11942 6664 11994
rect 6664 11942 6676 11994
rect 6676 11942 6690 11994
rect 6714 11942 6728 11994
rect 6728 11942 6740 11994
rect 6740 11942 6770 11994
rect 6794 11942 6804 11994
rect 6804 11942 6850 11994
rect 6554 11940 6610 11942
rect 6634 11940 6690 11942
rect 6714 11940 6770 11942
rect 6794 11940 6850 11942
rect 3755 9274 3811 9276
rect 3835 9274 3891 9276
rect 3915 9274 3971 9276
rect 3995 9274 4051 9276
rect 3755 9222 3801 9274
rect 3801 9222 3811 9274
rect 3835 9222 3865 9274
rect 3865 9222 3877 9274
rect 3877 9222 3891 9274
rect 3915 9222 3929 9274
rect 3929 9222 3941 9274
rect 3941 9222 3971 9274
rect 3995 9222 4005 9274
rect 4005 9222 4051 9274
rect 3755 9220 3811 9222
rect 3835 9220 3891 9222
rect 3915 9220 3971 9222
rect 3995 9220 4051 9222
rect 6554 10906 6610 10908
rect 6634 10906 6690 10908
rect 6714 10906 6770 10908
rect 6794 10906 6850 10908
rect 6554 10854 6600 10906
rect 6600 10854 6610 10906
rect 6634 10854 6664 10906
rect 6664 10854 6676 10906
rect 6676 10854 6690 10906
rect 6714 10854 6728 10906
rect 6728 10854 6740 10906
rect 6740 10854 6770 10906
rect 6794 10854 6804 10906
rect 6804 10854 6850 10906
rect 6554 10852 6610 10854
rect 6634 10852 6690 10854
rect 6714 10852 6770 10854
rect 6794 10852 6850 10854
rect 6826 10532 6882 10568
rect 6826 10512 6828 10532
rect 6828 10512 6880 10532
rect 6880 10512 6882 10532
rect 9353 15802 9409 15804
rect 9433 15802 9489 15804
rect 9513 15802 9569 15804
rect 9593 15802 9649 15804
rect 9353 15750 9399 15802
rect 9399 15750 9409 15802
rect 9433 15750 9463 15802
rect 9463 15750 9475 15802
rect 9475 15750 9489 15802
rect 9513 15750 9527 15802
rect 9527 15750 9539 15802
rect 9539 15750 9569 15802
rect 9593 15750 9603 15802
rect 9603 15750 9649 15802
rect 9353 15748 9409 15750
rect 9433 15748 9489 15750
rect 9513 15748 9569 15750
rect 9593 15748 9649 15750
rect 9353 14714 9409 14716
rect 9433 14714 9489 14716
rect 9513 14714 9569 14716
rect 9593 14714 9649 14716
rect 9353 14662 9399 14714
rect 9399 14662 9409 14714
rect 9433 14662 9463 14714
rect 9463 14662 9475 14714
rect 9475 14662 9489 14714
rect 9513 14662 9527 14714
rect 9527 14662 9539 14714
rect 9539 14662 9569 14714
rect 9593 14662 9603 14714
rect 9603 14662 9649 14714
rect 9353 14660 9409 14662
rect 9433 14660 9489 14662
rect 9513 14660 9569 14662
rect 9593 14660 9649 14662
rect 9353 13626 9409 13628
rect 9433 13626 9489 13628
rect 9513 13626 9569 13628
rect 9593 13626 9649 13628
rect 9353 13574 9399 13626
rect 9399 13574 9409 13626
rect 9433 13574 9463 13626
rect 9463 13574 9475 13626
rect 9475 13574 9489 13626
rect 9513 13574 9527 13626
rect 9527 13574 9539 13626
rect 9539 13574 9569 13626
rect 9593 13574 9603 13626
rect 9603 13574 9649 13626
rect 9353 13572 9409 13574
rect 9433 13572 9489 13574
rect 9513 13572 9569 13574
rect 9593 13572 9649 13574
rect 9353 12538 9409 12540
rect 9433 12538 9489 12540
rect 9513 12538 9569 12540
rect 9593 12538 9649 12540
rect 9353 12486 9399 12538
rect 9399 12486 9409 12538
rect 9433 12486 9463 12538
rect 9463 12486 9475 12538
rect 9475 12486 9489 12538
rect 9513 12486 9527 12538
rect 9527 12486 9539 12538
rect 9539 12486 9569 12538
rect 9593 12486 9603 12538
rect 9603 12486 9649 12538
rect 9353 12484 9409 12486
rect 9433 12484 9489 12486
rect 9513 12484 9569 12486
rect 9593 12484 9649 12486
rect 9353 11450 9409 11452
rect 9433 11450 9489 11452
rect 9513 11450 9569 11452
rect 9593 11450 9649 11452
rect 9353 11398 9399 11450
rect 9399 11398 9409 11450
rect 9433 11398 9463 11450
rect 9463 11398 9475 11450
rect 9475 11398 9489 11450
rect 9513 11398 9527 11450
rect 9527 11398 9539 11450
rect 9539 11398 9569 11450
rect 9593 11398 9603 11450
rect 9603 11398 9649 11450
rect 9353 11396 9409 11398
rect 9433 11396 9489 11398
rect 9513 11396 9569 11398
rect 9593 11396 9649 11398
rect 6554 9818 6610 9820
rect 6634 9818 6690 9820
rect 6714 9818 6770 9820
rect 6794 9818 6850 9820
rect 6554 9766 6600 9818
rect 6600 9766 6610 9818
rect 6634 9766 6664 9818
rect 6664 9766 6676 9818
rect 6676 9766 6690 9818
rect 6714 9766 6728 9818
rect 6728 9766 6740 9818
rect 6740 9766 6770 9818
rect 6794 9766 6804 9818
rect 6804 9766 6850 9818
rect 6554 9764 6610 9766
rect 6634 9764 6690 9766
rect 6714 9764 6770 9766
rect 6794 9764 6850 9766
rect 3755 8186 3811 8188
rect 3835 8186 3891 8188
rect 3915 8186 3971 8188
rect 3995 8186 4051 8188
rect 3755 8134 3801 8186
rect 3801 8134 3811 8186
rect 3835 8134 3865 8186
rect 3865 8134 3877 8186
rect 3877 8134 3891 8186
rect 3915 8134 3929 8186
rect 3929 8134 3941 8186
rect 3941 8134 3971 8186
rect 3995 8134 4005 8186
rect 4005 8134 4051 8186
rect 3755 8132 3811 8134
rect 3835 8132 3891 8134
rect 3915 8132 3971 8134
rect 3995 8132 4051 8134
rect 3755 7098 3811 7100
rect 3835 7098 3891 7100
rect 3915 7098 3971 7100
rect 3995 7098 4051 7100
rect 3755 7046 3801 7098
rect 3801 7046 3811 7098
rect 3835 7046 3865 7098
rect 3865 7046 3877 7098
rect 3877 7046 3891 7098
rect 3915 7046 3929 7098
rect 3929 7046 3941 7098
rect 3941 7046 3971 7098
rect 3995 7046 4005 7098
rect 4005 7046 4051 7098
rect 3755 7044 3811 7046
rect 3835 7044 3891 7046
rect 3915 7044 3971 7046
rect 3995 7044 4051 7046
rect 3755 6010 3811 6012
rect 3835 6010 3891 6012
rect 3915 6010 3971 6012
rect 3995 6010 4051 6012
rect 3755 5958 3801 6010
rect 3801 5958 3811 6010
rect 3835 5958 3865 6010
rect 3865 5958 3877 6010
rect 3877 5958 3891 6010
rect 3915 5958 3929 6010
rect 3929 5958 3941 6010
rect 3941 5958 3971 6010
rect 3995 5958 4005 6010
rect 4005 5958 4051 6010
rect 3755 5956 3811 5958
rect 3835 5956 3891 5958
rect 3915 5956 3971 5958
rect 3995 5956 4051 5958
rect 8114 10512 8170 10568
rect 9353 10362 9409 10364
rect 9433 10362 9489 10364
rect 9513 10362 9569 10364
rect 9593 10362 9649 10364
rect 9353 10310 9399 10362
rect 9399 10310 9409 10362
rect 9433 10310 9463 10362
rect 9463 10310 9475 10362
rect 9475 10310 9489 10362
rect 9513 10310 9527 10362
rect 9527 10310 9539 10362
rect 9539 10310 9569 10362
rect 9593 10310 9603 10362
rect 9603 10310 9649 10362
rect 9353 10308 9409 10310
rect 9433 10308 9489 10310
rect 9513 10308 9569 10310
rect 9593 10308 9649 10310
rect 6554 8730 6610 8732
rect 6634 8730 6690 8732
rect 6714 8730 6770 8732
rect 6794 8730 6850 8732
rect 6554 8678 6600 8730
rect 6600 8678 6610 8730
rect 6634 8678 6664 8730
rect 6664 8678 6676 8730
rect 6676 8678 6690 8730
rect 6714 8678 6728 8730
rect 6728 8678 6740 8730
rect 6740 8678 6770 8730
rect 6794 8678 6804 8730
rect 6804 8678 6850 8730
rect 6554 8676 6610 8678
rect 6634 8676 6690 8678
rect 6714 8676 6770 8678
rect 6794 8676 6850 8678
rect 6554 7642 6610 7644
rect 6634 7642 6690 7644
rect 6714 7642 6770 7644
rect 6794 7642 6850 7644
rect 6554 7590 6600 7642
rect 6600 7590 6610 7642
rect 6634 7590 6664 7642
rect 6664 7590 6676 7642
rect 6676 7590 6690 7642
rect 6714 7590 6728 7642
rect 6728 7590 6740 7642
rect 6740 7590 6770 7642
rect 6794 7590 6804 7642
rect 6804 7590 6850 7642
rect 6554 7588 6610 7590
rect 6634 7588 6690 7590
rect 6714 7588 6770 7590
rect 6794 7588 6850 7590
rect 6554 6554 6610 6556
rect 6634 6554 6690 6556
rect 6714 6554 6770 6556
rect 6794 6554 6850 6556
rect 6554 6502 6600 6554
rect 6600 6502 6610 6554
rect 6634 6502 6664 6554
rect 6664 6502 6676 6554
rect 6676 6502 6690 6554
rect 6714 6502 6728 6554
rect 6728 6502 6740 6554
rect 6740 6502 6770 6554
rect 6794 6502 6804 6554
rect 6804 6502 6850 6554
rect 6554 6500 6610 6502
rect 6634 6500 6690 6502
rect 6714 6500 6770 6502
rect 6794 6500 6850 6502
rect 6554 5466 6610 5468
rect 6634 5466 6690 5468
rect 6714 5466 6770 5468
rect 6794 5466 6850 5468
rect 6554 5414 6600 5466
rect 6600 5414 6610 5466
rect 6634 5414 6664 5466
rect 6664 5414 6676 5466
rect 6676 5414 6690 5466
rect 6714 5414 6728 5466
rect 6728 5414 6740 5466
rect 6740 5414 6770 5466
rect 6794 5414 6804 5466
rect 6804 5414 6850 5466
rect 6554 5412 6610 5414
rect 6634 5412 6690 5414
rect 6714 5412 6770 5414
rect 6794 5412 6850 5414
rect 3755 4922 3811 4924
rect 3835 4922 3891 4924
rect 3915 4922 3971 4924
rect 3995 4922 4051 4924
rect 3755 4870 3801 4922
rect 3801 4870 3811 4922
rect 3835 4870 3865 4922
rect 3865 4870 3877 4922
rect 3877 4870 3891 4922
rect 3915 4870 3929 4922
rect 3929 4870 3941 4922
rect 3941 4870 3971 4922
rect 3995 4870 4005 4922
rect 4005 4870 4051 4922
rect 3755 4868 3811 4870
rect 3835 4868 3891 4870
rect 3915 4868 3971 4870
rect 3995 4868 4051 4870
rect 6554 4378 6610 4380
rect 6634 4378 6690 4380
rect 6714 4378 6770 4380
rect 6794 4378 6850 4380
rect 6554 4326 6600 4378
rect 6600 4326 6610 4378
rect 6634 4326 6664 4378
rect 6664 4326 6676 4378
rect 6676 4326 6690 4378
rect 6714 4326 6728 4378
rect 6728 4326 6740 4378
rect 6740 4326 6770 4378
rect 6794 4326 6804 4378
rect 6804 4326 6850 4378
rect 6554 4324 6610 4326
rect 6634 4324 6690 4326
rect 6714 4324 6770 4326
rect 6794 4324 6850 4326
rect 9353 9274 9409 9276
rect 9433 9274 9489 9276
rect 9513 9274 9569 9276
rect 9593 9274 9649 9276
rect 9353 9222 9399 9274
rect 9399 9222 9409 9274
rect 9433 9222 9463 9274
rect 9463 9222 9475 9274
rect 9475 9222 9489 9274
rect 9513 9222 9527 9274
rect 9527 9222 9539 9274
rect 9539 9222 9569 9274
rect 9593 9222 9603 9274
rect 9603 9222 9649 9274
rect 9353 9220 9409 9222
rect 9433 9220 9489 9222
rect 9513 9220 9569 9222
rect 9593 9220 9649 9222
rect 9353 8186 9409 8188
rect 9433 8186 9489 8188
rect 9513 8186 9569 8188
rect 9593 8186 9649 8188
rect 9353 8134 9399 8186
rect 9399 8134 9409 8186
rect 9433 8134 9463 8186
rect 9463 8134 9475 8186
rect 9475 8134 9489 8186
rect 9513 8134 9527 8186
rect 9527 8134 9539 8186
rect 9539 8134 9569 8186
rect 9593 8134 9603 8186
rect 9603 8134 9649 8186
rect 9353 8132 9409 8134
rect 9433 8132 9489 8134
rect 9513 8132 9569 8134
rect 9593 8132 9649 8134
rect 9353 7098 9409 7100
rect 9433 7098 9489 7100
rect 9513 7098 9569 7100
rect 9593 7098 9649 7100
rect 9353 7046 9399 7098
rect 9399 7046 9409 7098
rect 9433 7046 9463 7098
rect 9463 7046 9475 7098
rect 9475 7046 9489 7098
rect 9513 7046 9527 7098
rect 9527 7046 9539 7098
rect 9539 7046 9569 7098
rect 9593 7046 9603 7098
rect 9603 7046 9649 7098
rect 9353 7044 9409 7046
rect 9433 7044 9489 7046
rect 9513 7044 9569 7046
rect 9593 7044 9649 7046
rect 9353 6010 9409 6012
rect 9433 6010 9489 6012
rect 9513 6010 9569 6012
rect 9593 6010 9649 6012
rect 9353 5958 9399 6010
rect 9399 5958 9409 6010
rect 9433 5958 9463 6010
rect 9463 5958 9475 6010
rect 9475 5958 9489 6010
rect 9513 5958 9527 6010
rect 9527 5958 9539 6010
rect 9539 5958 9569 6010
rect 9593 5958 9603 6010
rect 9603 5958 9649 6010
rect 9353 5956 9409 5958
rect 9433 5956 9489 5958
rect 9513 5956 9569 5958
rect 9593 5956 9649 5958
rect 11426 21392 11482 21448
rect 11334 19372 11390 19408
rect 11334 19352 11336 19372
rect 11336 19352 11388 19372
rect 11388 19352 11390 19372
rect 11426 17720 11482 17776
rect 11334 17584 11390 17640
rect 11150 16496 11206 16552
rect 10690 16088 10746 16144
rect 12152 21786 12208 21788
rect 12232 21786 12288 21788
rect 12312 21786 12368 21788
rect 12392 21786 12448 21788
rect 12152 21734 12198 21786
rect 12198 21734 12208 21786
rect 12232 21734 12262 21786
rect 12262 21734 12274 21786
rect 12274 21734 12288 21786
rect 12312 21734 12326 21786
rect 12326 21734 12338 21786
rect 12338 21734 12368 21786
rect 12392 21734 12402 21786
rect 12402 21734 12448 21786
rect 12152 21732 12208 21734
rect 12232 21732 12288 21734
rect 12312 21732 12368 21734
rect 12392 21732 12448 21734
rect 12152 20698 12208 20700
rect 12232 20698 12288 20700
rect 12312 20698 12368 20700
rect 12392 20698 12448 20700
rect 12152 20646 12198 20698
rect 12198 20646 12208 20698
rect 12232 20646 12262 20698
rect 12262 20646 12274 20698
rect 12274 20646 12288 20698
rect 12312 20646 12326 20698
rect 12326 20646 12338 20698
rect 12338 20646 12368 20698
rect 12392 20646 12402 20698
rect 12402 20646 12448 20698
rect 12152 20644 12208 20646
rect 12232 20644 12288 20646
rect 12312 20644 12368 20646
rect 12392 20644 12448 20646
rect 11058 12708 11114 12744
rect 11058 12688 11060 12708
rect 11060 12688 11112 12708
rect 11112 12688 11114 12708
rect 11702 12280 11758 12336
rect 10782 7248 10838 7304
rect 10690 6840 10746 6896
rect 9353 4922 9409 4924
rect 9433 4922 9489 4924
rect 9513 4922 9569 4924
rect 9593 4922 9649 4924
rect 9353 4870 9399 4922
rect 9399 4870 9409 4922
rect 9433 4870 9463 4922
rect 9463 4870 9475 4922
rect 9475 4870 9489 4922
rect 9513 4870 9527 4922
rect 9527 4870 9539 4922
rect 9539 4870 9569 4922
rect 9593 4870 9603 4922
rect 9603 4870 9649 4922
rect 9353 4868 9409 4870
rect 9433 4868 9489 4870
rect 9513 4868 9569 4870
rect 9593 4868 9649 4870
rect 3755 3834 3811 3836
rect 3835 3834 3891 3836
rect 3915 3834 3971 3836
rect 3995 3834 4051 3836
rect 3755 3782 3801 3834
rect 3801 3782 3811 3834
rect 3835 3782 3865 3834
rect 3865 3782 3877 3834
rect 3877 3782 3891 3834
rect 3915 3782 3929 3834
rect 3929 3782 3941 3834
rect 3941 3782 3971 3834
rect 3995 3782 4005 3834
rect 4005 3782 4051 3834
rect 3755 3780 3811 3782
rect 3835 3780 3891 3782
rect 3915 3780 3971 3782
rect 3995 3780 4051 3782
rect 9353 3834 9409 3836
rect 9433 3834 9489 3836
rect 9513 3834 9569 3836
rect 9593 3834 9649 3836
rect 9353 3782 9399 3834
rect 9399 3782 9409 3834
rect 9433 3782 9463 3834
rect 9463 3782 9475 3834
rect 9475 3782 9489 3834
rect 9513 3782 9527 3834
rect 9527 3782 9539 3834
rect 9539 3782 9569 3834
rect 9593 3782 9603 3834
rect 9603 3782 9649 3834
rect 9353 3780 9409 3782
rect 9433 3780 9489 3782
rect 9513 3780 9569 3782
rect 9593 3780 9649 3782
rect 12152 19610 12208 19612
rect 12232 19610 12288 19612
rect 12312 19610 12368 19612
rect 12392 19610 12448 19612
rect 12152 19558 12198 19610
rect 12198 19558 12208 19610
rect 12232 19558 12262 19610
rect 12262 19558 12274 19610
rect 12274 19558 12288 19610
rect 12312 19558 12326 19610
rect 12326 19558 12338 19610
rect 12338 19558 12368 19610
rect 12392 19558 12402 19610
rect 12402 19558 12448 19610
rect 12152 19556 12208 19558
rect 12232 19556 12288 19558
rect 12312 19556 12368 19558
rect 12392 19556 12448 19558
rect 12152 18522 12208 18524
rect 12232 18522 12288 18524
rect 12312 18522 12368 18524
rect 12392 18522 12448 18524
rect 12152 18470 12198 18522
rect 12198 18470 12208 18522
rect 12232 18470 12262 18522
rect 12262 18470 12274 18522
rect 12274 18470 12288 18522
rect 12312 18470 12326 18522
rect 12326 18470 12338 18522
rect 12338 18470 12368 18522
rect 12392 18470 12402 18522
rect 12402 18470 12448 18522
rect 12152 18468 12208 18470
rect 12232 18468 12288 18470
rect 12312 18468 12368 18470
rect 12392 18468 12448 18470
rect 13174 22208 13230 22264
rect 12714 19896 12770 19952
rect 12898 19488 12954 19544
rect 13266 21800 13322 21856
rect 13266 21528 13322 21584
rect 13726 21020 13728 21040
rect 13728 21020 13780 21040
rect 13780 21020 13782 21040
rect 13726 20984 13782 21020
rect 13634 20576 13690 20632
rect 13266 19896 13322 19952
rect 13082 18400 13138 18456
rect 12990 18264 13046 18320
rect 13726 17720 13782 17776
rect 12152 17434 12208 17436
rect 12232 17434 12288 17436
rect 12312 17434 12368 17436
rect 12392 17434 12448 17436
rect 12152 17382 12198 17434
rect 12198 17382 12208 17434
rect 12232 17382 12262 17434
rect 12262 17382 12274 17434
rect 12274 17382 12288 17434
rect 12312 17382 12326 17434
rect 12326 17382 12338 17434
rect 12338 17382 12368 17434
rect 12392 17382 12402 17434
rect 12402 17382 12448 17434
rect 12152 17380 12208 17382
rect 12232 17380 12288 17382
rect 12312 17380 12368 17382
rect 12392 17380 12448 17382
rect 12152 16346 12208 16348
rect 12232 16346 12288 16348
rect 12312 16346 12368 16348
rect 12392 16346 12448 16348
rect 12152 16294 12198 16346
rect 12198 16294 12208 16346
rect 12232 16294 12262 16346
rect 12262 16294 12274 16346
rect 12274 16294 12288 16346
rect 12312 16294 12326 16346
rect 12326 16294 12338 16346
rect 12338 16294 12368 16346
rect 12392 16294 12402 16346
rect 12402 16294 12448 16346
rect 12152 16292 12208 16294
rect 12232 16292 12288 16294
rect 12312 16292 12368 16294
rect 12392 16292 12448 16294
rect 12254 15544 12310 15600
rect 12152 15258 12208 15260
rect 12232 15258 12288 15260
rect 12312 15258 12368 15260
rect 12392 15258 12448 15260
rect 12152 15206 12198 15258
rect 12198 15206 12208 15258
rect 12232 15206 12262 15258
rect 12262 15206 12274 15258
rect 12274 15206 12288 15258
rect 12312 15206 12326 15258
rect 12326 15206 12338 15258
rect 12338 15206 12368 15258
rect 12392 15206 12402 15258
rect 12402 15206 12448 15258
rect 12152 15204 12208 15206
rect 12232 15204 12288 15206
rect 12312 15204 12368 15206
rect 12392 15204 12448 15206
rect 12152 14170 12208 14172
rect 12232 14170 12288 14172
rect 12312 14170 12368 14172
rect 12392 14170 12448 14172
rect 12152 14118 12198 14170
rect 12198 14118 12208 14170
rect 12232 14118 12262 14170
rect 12262 14118 12274 14170
rect 12274 14118 12288 14170
rect 12312 14118 12326 14170
rect 12326 14118 12338 14170
rect 12338 14118 12368 14170
rect 12392 14118 12402 14170
rect 12402 14118 12448 14170
rect 12152 14116 12208 14118
rect 12232 14116 12288 14118
rect 12312 14116 12368 14118
rect 12392 14116 12448 14118
rect 12152 13082 12208 13084
rect 12232 13082 12288 13084
rect 12312 13082 12368 13084
rect 12392 13082 12448 13084
rect 12152 13030 12198 13082
rect 12198 13030 12208 13082
rect 12232 13030 12262 13082
rect 12262 13030 12274 13082
rect 12274 13030 12288 13082
rect 12312 13030 12326 13082
rect 12326 13030 12338 13082
rect 12338 13030 12368 13082
rect 12392 13030 12402 13082
rect 12402 13030 12448 13082
rect 12152 13028 12208 13030
rect 12232 13028 12288 13030
rect 12312 13028 12368 13030
rect 12392 13028 12448 13030
rect 12152 11994 12208 11996
rect 12232 11994 12288 11996
rect 12312 11994 12368 11996
rect 12392 11994 12448 11996
rect 12152 11942 12198 11994
rect 12198 11942 12208 11994
rect 12232 11942 12262 11994
rect 12262 11942 12274 11994
rect 12274 11942 12288 11994
rect 12312 11942 12326 11994
rect 12326 11942 12338 11994
rect 12338 11942 12368 11994
rect 12392 11942 12402 11994
rect 12402 11942 12448 11994
rect 12152 11940 12208 11942
rect 12232 11940 12288 11942
rect 12312 11940 12368 11942
rect 12392 11940 12448 11942
rect 12152 10906 12208 10908
rect 12232 10906 12288 10908
rect 12312 10906 12368 10908
rect 12392 10906 12448 10908
rect 12152 10854 12198 10906
rect 12198 10854 12208 10906
rect 12232 10854 12262 10906
rect 12262 10854 12274 10906
rect 12274 10854 12288 10906
rect 12312 10854 12326 10906
rect 12326 10854 12338 10906
rect 12338 10854 12368 10906
rect 12392 10854 12402 10906
rect 12402 10854 12448 10906
rect 12152 10852 12208 10854
rect 12232 10852 12288 10854
rect 12312 10852 12368 10854
rect 12392 10852 12448 10854
rect 12152 9818 12208 9820
rect 12232 9818 12288 9820
rect 12312 9818 12368 9820
rect 12392 9818 12448 9820
rect 12152 9766 12198 9818
rect 12198 9766 12208 9818
rect 12232 9766 12262 9818
rect 12262 9766 12274 9818
rect 12274 9766 12288 9818
rect 12312 9766 12326 9818
rect 12326 9766 12338 9818
rect 12338 9766 12368 9818
rect 12392 9766 12402 9818
rect 12402 9766 12448 9818
rect 12152 9764 12208 9766
rect 12232 9764 12288 9766
rect 12312 9764 12368 9766
rect 12392 9764 12448 9766
rect 12152 8730 12208 8732
rect 12232 8730 12288 8732
rect 12312 8730 12368 8732
rect 12392 8730 12448 8732
rect 12152 8678 12198 8730
rect 12198 8678 12208 8730
rect 12232 8678 12262 8730
rect 12262 8678 12274 8730
rect 12274 8678 12288 8730
rect 12312 8678 12326 8730
rect 12326 8678 12338 8730
rect 12338 8678 12368 8730
rect 12392 8678 12402 8730
rect 12402 8678 12448 8730
rect 12152 8676 12208 8678
rect 12232 8676 12288 8678
rect 12312 8676 12368 8678
rect 12392 8676 12448 8678
rect 12070 7792 12126 7848
rect 12152 7642 12208 7644
rect 12232 7642 12288 7644
rect 12312 7642 12368 7644
rect 12392 7642 12448 7644
rect 12152 7590 12198 7642
rect 12198 7590 12208 7642
rect 12232 7590 12262 7642
rect 12262 7590 12274 7642
rect 12274 7590 12288 7642
rect 12312 7590 12326 7642
rect 12326 7590 12338 7642
rect 12338 7590 12368 7642
rect 12392 7590 12402 7642
rect 12402 7590 12448 7642
rect 12152 7588 12208 7590
rect 12232 7588 12288 7590
rect 12312 7588 12368 7590
rect 12392 7588 12448 7590
rect 12152 6554 12208 6556
rect 12232 6554 12288 6556
rect 12312 6554 12368 6556
rect 12392 6554 12448 6556
rect 12152 6502 12198 6554
rect 12198 6502 12208 6554
rect 12232 6502 12262 6554
rect 12262 6502 12274 6554
rect 12274 6502 12288 6554
rect 12312 6502 12326 6554
rect 12326 6502 12338 6554
rect 12338 6502 12368 6554
rect 12392 6502 12402 6554
rect 12402 6502 12448 6554
rect 12152 6500 12208 6502
rect 12232 6500 12288 6502
rect 12312 6500 12368 6502
rect 12392 6500 12448 6502
rect 13266 14320 13322 14376
rect 14951 22330 15007 22332
rect 15031 22330 15087 22332
rect 15111 22330 15167 22332
rect 15191 22330 15247 22332
rect 14951 22278 14997 22330
rect 14997 22278 15007 22330
rect 15031 22278 15061 22330
rect 15061 22278 15073 22330
rect 15073 22278 15087 22330
rect 15111 22278 15125 22330
rect 15125 22278 15137 22330
rect 15137 22278 15167 22330
rect 15191 22278 15201 22330
rect 15201 22278 15247 22330
rect 14951 22276 15007 22278
rect 15031 22276 15087 22278
rect 15111 22276 15167 22278
rect 15191 22276 15247 22278
rect 14462 20712 14518 20768
rect 14554 19352 14610 19408
rect 14278 18400 14334 18456
rect 14278 18284 14334 18320
rect 14278 18264 14280 18284
rect 14280 18264 14332 18284
rect 14332 18264 14334 18284
rect 12806 6160 12862 6216
rect 13542 7384 13598 7440
rect 14462 18672 14518 18728
rect 15290 21800 15346 21856
rect 14951 21242 15007 21244
rect 15031 21242 15087 21244
rect 15111 21242 15167 21244
rect 15191 21242 15247 21244
rect 14951 21190 14997 21242
rect 14997 21190 15007 21242
rect 15031 21190 15061 21242
rect 15061 21190 15073 21242
rect 15073 21190 15087 21242
rect 15111 21190 15125 21242
rect 15125 21190 15137 21242
rect 15137 21190 15167 21242
rect 15191 21190 15201 21242
rect 15201 21190 15247 21242
rect 14951 21188 15007 21190
rect 15031 21188 15087 21190
rect 15111 21188 15167 21190
rect 15191 21188 15247 21190
rect 15382 20884 15384 20904
rect 15384 20884 15436 20904
rect 15436 20884 15438 20904
rect 15382 20848 15438 20884
rect 14951 20154 15007 20156
rect 15031 20154 15087 20156
rect 15111 20154 15167 20156
rect 15191 20154 15247 20156
rect 14951 20102 14997 20154
rect 14997 20102 15007 20154
rect 15031 20102 15061 20154
rect 15061 20102 15073 20154
rect 15073 20102 15087 20154
rect 15111 20102 15125 20154
rect 15125 20102 15137 20154
rect 15137 20102 15167 20154
rect 15191 20102 15201 20154
rect 15201 20102 15247 20154
rect 14951 20100 15007 20102
rect 15031 20100 15087 20102
rect 15111 20100 15167 20102
rect 15191 20100 15247 20102
rect 14951 19066 15007 19068
rect 15031 19066 15087 19068
rect 15111 19066 15167 19068
rect 15191 19066 15247 19068
rect 14951 19014 14997 19066
rect 14997 19014 15007 19066
rect 15031 19014 15061 19066
rect 15061 19014 15073 19066
rect 15073 19014 15087 19066
rect 15111 19014 15125 19066
rect 15125 19014 15137 19066
rect 15137 19014 15167 19066
rect 15191 19014 15201 19066
rect 15201 19014 15247 19066
rect 14951 19012 15007 19014
rect 15031 19012 15087 19014
rect 15111 19012 15167 19014
rect 15191 19012 15247 19014
rect 14922 18400 14978 18456
rect 15290 18264 15346 18320
rect 14951 17978 15007 17980
rect 15031 17978 15087 17980
rect 15111 17978 15167 17980
rect 15191 17978 15247 17980
rect 14951 17926 14997 17978
rect 14997 17926 15007 17978
rect 15031 17926 15061 17978
rect 15061 17926 15073 17978
rect 15073 17926 15087 17978
rect 15111 17926 15125 17978
rect 15125 17926 15137 17978
rect 15137 17926 15167 17978
rect 15191 17926 15201 17978
rect 15201 17926 15247 17978
rect 14951 17924 15007 17926
rect 15031 17924 15087 17926
rect 15111 17924 15167 17926
rect 15191 17924 15247 17926
rect 14462 17060 14518 17096
rect 14462 17040 14464 17060
rect 14464 17040 14516 17060
rect 14516 17040 14518 17060
rect 14951 16890 15007 16892
rect 15031 16890 15087 16892
rect 15111 16890 15167 16892
rect 15191 16890 15247 16892
rect 14951 16838 14997 16890
rect 14997 16838 15007 16890
rect 15031 16838 15061 16890
rect 15061 16838 15073 16890
rect 15073 16838 15087 16890
rect 15111 16838 15125 16890
rect 15125 16838 15137 16890
rect 15137 16838 15167 16890
rect 15191 16838 15201 16890
rect 15201 16838 15247 16890
rect 14951 16836 15007 16838
rect 15031 16836 15087 16838
rect 15111 16836 15167 16838
rect 15191 16836 15247 16838
rect 14951 15802 15007 15804
rect 15031 15802 15087 15804
rect 15111 15802 15167 15804
rect 15191 15802 15247 15804
rect 14951 15750 14997 15802
rect 14997 15750 15007 15802
rect 15031 15750 15061 15802
rect 15061 15750 15073 15802
rect 15073 15750 15087 15802
rect 15111 15750 15125 15802
rect 15125 15750 15137 15802
rect 15137 15750 15167 15802
rect 15191 15750 15201 15802
rect 15201 15750 15247 15802
rect 14951 15748 15007 15750
rect 15031 15748 15087 15750
rect 15111 15748 15167 15750
rect 15191 15748 15247 15750
rect 14951 14714 15007 14716
rect 15031 14714 15087 14716
rect 15111 14714 15167 14716
rect 15191 14714 15247 14716
rect 14951 14662 14997 14714
rect 14997 14662 15007 14714
rect 15031 14662 15061 14714
rect 15061 14662 15073 14714
rect 15073 14662 15087 14714
rect 15111 14662 15125 14714
rect 15125 14662 15137 14714
rect 15137 14662 15167 14714
rect 15191 14662 15201 14714
rect 15201 14662 15247 14714
rect 14951 14660 15007 14662
rect 15031 14660 15087 14662
rect 15111 14660 15167 14662
rect 15191 14660 15247 14662
rect 15014 14456 15070 14512
rect 15658 20032 15714 20088
rect 15934 21800 15990 21856
rect 15842 21664 15898 21720
rect 15934 21120 15990 21176
rect 16118 19488 16174 19544
rect 16302 21528 16358 21584
rect 16210 17176 16266 17232
rect 15198 13932 15254 13968
rect 15198 13912 15200 13932
rect 15200 13912 15252 13932
rect 15252 13912 15254 13932
rect 14951 13626 15007 13628
rect 15031 13626 15087 13628
rect 15111 13626 15167 13628
rect 15191 13626 15247 13628
rect 14951 13574 14997 13626
rect 14997 13574 15007 13626
rect 15031 13574 15061 13626
rect 15061 13574 15073 13626
rect 15073 13574 15087 13626
rect 15111 13574 15125 13626
rect 15125 13574 15137 13626
rect 15137 13574 15167 13626
rect 15191 13574 15201 13626
rect 15201 13574 15247 13626
rect 14951 13572 15007 13574
rect 15031 13572 15087 13574
rect 15111 13572 15167 13574
rect 15191 13572 15247 13574
rect 15106 13404 15108 13424
rect 15108 13404 15160 13424
rect 15160 13404 15162 13424
rect 15106 13368 15162 13404
rect 14646 13232 14702 13288
rect 14951 12538 15007 12540
rect 15031 12538 15087 12540
rect 15111 12538 15167 12540
rect 15191 12538 15247 12540
rect 14951 12486 14997 12538
rect 14997 12486 15007 12538
rect 15031 12486 15061 12538
rect 15061 12486 15073 12538
rect 15073 12486 15087 12538
rect 15111 12486 15125 12538
rect 15125 12486 15137 12538
rect 15137 12486 15167 12538
rect 15191 12486 15201 12538
rect 15201 12486 15247 12538
rect 14951 12484 15007 12486
rect 15031 12484 15087 12486
rect 15111 12484 15167 12486
rect 15191 12484 15247 12486
rect 14951 11450 15007 11452
rect 15031 11450 15087 11452
rect 15111 11450 15167 11452
rect 15191 11450 15247 11452
rect 14951 11398 14997 11450
rect 14997 11398 15007 11450
rect 15031 11398 15061 11450
rect 15061 11398 15073 11450
rect 15073 11398 15087 11450
rect 15111 11398 15125 11450
rect 15125 11398 15137 11450
rect 15137 11398 15167 11450
rect 15191 11398 15201 11450
rect 15201 11398 15247 11450
rect 14951 11396 15007 11398
rect 15031 11396 15087 11398
rect 15111 11396 15167 11398
rect 15191 11396 15247 11398
rect 14951 10362 15007 10364
rect 15031 10362 15087 10364
rect 15111 10362 15167 10364
rect 15191 10362 15247 10364
rect 14951 10310 14997 10362
rect 14997 10310 15007 10362
rect 15031 10310 15061 10362
rect 15061 10310 15073 10362
rect 15073 10310 15087 10362
rect 15111 10310 15125 10362
rect 15125 10310 15137 10362
rect 15137 10310 15167 10362
rect 15191 10310 15201 10362
rect 15201 10310 15247 10362
rect 14951 10308 15007 10310
rect 15031 10308 15087 10310
rect 15111 10308 15167 10310
rect 15191 10308 15247 10310
rect 14951 9274 15007 9276
rect 15031 9274 15087 9276
rect 15111 9274 15167 9276
rect 15191 9274 15247 9276
rect 14951 9222 14997 9274
rect 14997 9222 15007 9274
rect 15031 9222 15061 9274
rect 15061 9222 15073 9274
rect 15073 9222 15087 9274
rect 15111 9222 15125 9274
rect 15125 9222 15137 9274
rect 15137 9222 15167 9274
rect 15191 9222 15201 9274
rect 15201 9222 15247 9274
rect 14951 9220 15007 9222
rect 15031 9220 15087 9222
rect 15111 9220 15167 9222
rect 15191 9220 15247 9222
rect 14951 8186 15007 8188
rect 15031 8186 15087 8188
rect 15111 8186 15167 8188
rect 15191 8186 15247 8188
rect 14951 8134 14997 8186
rect 14997 8134 15007 8186
rect 15031 8134 15061 8186
rect 15061 8134 15073 8186
rect 15073 8134 15087 8186
rect 15111 8134 15125 8186
rect 15125 8134 15137 8186
rect 15137 8134 15167 8186
rect 15191 8134 15201 8186
rect 15201 8134 15247 8186
rect 14951 8132 15007 8134
rect 15031 8132 15087 8134
rect 15111 8132 15167 8134
rect 15191 8132 15247 8134
rect 11242 5752 11298 5808
rect 12152 5466 12208 5468
rect 12232 5466 12288 5468
rect 12312 5466 12368 5468
rect 12392 5466 12448 5468
rect 12152 5414 12198 5466
rect 12198 5414 12208 5466
rect 12232 5414 12262 5466
rect 12262 5414 12274 5466
rect 12274 5414 12288 5466
rect 12312 5414 12326 5466
rect 12326 5414 12338 5466
rect 12338 5414 12368 5466
rect 12392 5414 12402 5466
rect 12402 5414 12448 5466
rect 12152 5412 12208 5414
rect 12232 5412 12288 5414
rect 12312 5412 12368 5414
rect 12392 5412 12448 5414
rect 6554 3290 6610 3292
rect 6634 3290 6690 3292
rect 6714 3290 6770 3292
rect 6794 3290 6850 3292
rect 6554 3238 6600 3290
rect 6600 3238 6610 3290
rect 6634 3238 6664 3290
rect 6664 3238 6676 3290
rect 6676 3238 6690 3290
rect 6714 3238 6728 3290
rect 6728 3238 6740 3290
rect 6740 3238 6770 3290
rect 6794 3238 6804 3290
rect 6804 3238 6850 3290
rect 6554 3236 6610 3238
rect 6634 3236 6690 3238
rect 6714 3236 6770 3238
rect 6794 3236 6850 3238
rect 1398 3032 1454 3088
rect 12152 4378 12208 4380
rect 12232 4378 12288 4380
rect 12312 4378 12368 4380
rect 12392 4378 12448 4380
rect 12152 4326 12198 4378
rect 12198 4326 12208 4378
rect 12232 4326 12262 4378
rect 12262 4326 12274 4378
rect 12274 4326 12288 4378
rect 12312 4326 12326 4378
rect 12326 4326 12338 4378
rect 12338 4326 12368 4378
rect 12392 4326 12402 4378
rect 12402 4326 12448 4378
rect 12152 4324 12208 4326
rect 12232 4324 12288 4326
rect 12312 4324 12368 4326
rect 12392 4324 12448 4326
rect 12152 3290 12208 3292
rect 12232 3290 12288 3292
rect 12312 3290 12368 3292
rect 12392 3290 12448 3292
rect 12152 3238 12198 3290
rect 12198 3238 12208 3290
rect 12232 3238 12262 3290
rect 12262 3238 12274 3290
rect 12274 3238 12288 3290
rect 12312 3238 12326 3290
rect 12326 3238 12338 3290
rect 12338 3238 12368 3290
rect 12392 3238 12402 3290
rect 12402 3238 12448 3290
rect 12152 3236 12208 3238
rect 12232 3236 12288 3238
rect 12312 3236 12368 3238
rect 12392 3236 12448 3238
rect 14951 7098 15007 7100
rect 15031 7098 15087 7100
rect 15111 7098 15167 7100
rect 15191 7098 15247 7100
rect 14951 7046 14997 7098
rect 14997 7046 15007 7098
rect 15031 7046 15061 7098
rect 15061 7046 15073 7098
rect 15073 7046 15087 7098
rect 15111 7046 15125 7098
rect 15125 7046 15137 7098
rect 15137 7046 15167 7098
rect 15191 7046 15201 7098
rect 15201 7046 15247 7098
rect 14951 7044 15007 7046
rect 15031 7044 15087 7046
rect 15111 7044 15167 7046
rect 15191 7044 15247 7046
rect 15198 6724 15254 6760
rect 15198 6704 15200 6724
rect 15200 6704 15252 6724
rect 15252 6704 15254 6724
rect 14951 6010 15007 6012
rect 15031 6010 15087 6012
rect 15111 6010 15167 6012
rect 15191 6010 15247 6012
rect 14951 5958 14997 6010
rect 14997 5958 15007 6010
rect 15031 5958 15061 6010
rect 15061 5958 15073 6010
rect 15073 5958 15087 6010
rect 15111 5958 15125 6010
rect 15125 5958 15137 6010
rect 15137 5958 15167 6010
rect 15191 5958 15201 6010
rect 15201 5958 15247 6010
rect 14951 5956 15007 5958
rect 15031 5956 15087 5958
rect 15111 5956 15167 5958
rect 15191 5956 15247 5958
rect 16486 20168 16542 20224
rect 16670 20868 16726 20904
rect 16670 20848 16672 20868
rect 16672 20848 16724 20868
rect 16724 20848 16726 20868
rect 16486 19488 16542 19544
rect 16394 19372 16450 19408
rect 18234 22480 18290 22536
rect 17130 21528 17186 21584
rect 17038 20712 17094 20768
rect 16946 20440 17002 20496
rect 16394 19352 16396 19372
rect 16396 19352 16448 19372
rect 16448 19352 16450 19372
rect 16578 19352 16634 19408
rect 16578 19216 16634 19272
rect 16486 15972 16542 16008
rect 16486 15952 16488 15972
rect 16488 15952 16540 15972
rect 16540 15952 16542 15972
rect 16670 15408 16726 15464
rect 16578 15136 16634 15192
rect 16486 14220 16488 14240
rect 16488 14220 16540 14240
rect 16540 14220 16542 14240
rect 16486 14184 16542 14220
rect 15474 10648 15530 10704
rect 14951 4922 15007 4924
rect 15031 4922 15087 4924
rect 15111 4922 15167 4924
rect 15191 4922 15247 4924
rect 14951 4870 14997 4922
rect 14997 4870 15007 4922
rect 15031 4870 15061 4922
rect 15061 4870 15073 4922
rect 15073 4870 15087 4922
rect 15111 4870 15125 4922
rect 15125 4870 15137 4922
rect 15137 4870 15167 4922
rect 15191 4870 15201 4922
rect 15201 4870 15247 4922
rect 14951 4868 15007 4870
rect 15031 4868 15087 4870
rect 15111 4868 15167 4870
rect 15191 4868 15247 4870
rect 14951 3834 15007 3836
rect 15031 3834 15087 3836
rect 15111 3834 15167 3836
rect 15191 3834 15247 3836
rect 14951 3782 14997 3834
rect 14997 3782 15007 3834
rect 15031 3782 15061 3834
rect 15061 3782 15073 3834
rect 15073 3782 15087 3834
rect 15111 3782 15125 3834
rect 15125 3782 15137 3834
rect 15137 3782 15167 3834
rect 15191 3782 15201 3834
rect 15201 3782 15247 3834
rect 14951 3780 15007 3782
rect 15031 3780 15087 3782
rect 15111 3780 15167 3782
rect 15191 3780 15247 3782
rect 3755 2746 3811 2748
rect 3835 2746 3891 2748
rect 3915 2746 3971 2748
rect 3995 2746 4051 2748
rect 3755 2694 3801 2746
rect 3801 2694 3811 2746
rect 3835 2694 3865 2746
rect 3865 2694 3877 2746
rect 3877 2694 3891 2746
rect 3915 2694 3929 2746
rect 3929 2694 3941 2746
rect 3941 2694 3971 2746
rect 3995 2694 4005 2746
rect 4005 2694 4051 2746
rect 3755 2692 3811 2694
rect 3835 2692 3891 2694
rect 3915 2692 3971 2694
rect 3995 2692 4051 2694
rect 9353 2746 9409 2748
rect 9433 2746 9489 2748
rect 9513 2746 9569 2748
rect 9593 2746 9649 2748
rect 9353 2694 9399 2746
rect 9399 2694 9409 2746
rect 9433 2694 9463 2746
rect 9463 2694 9475 2746
rect 9475 2694 9489 2746
rect 9513 2694 9527 2746
rect 9527 2694 9539 2746
rect 9539 2694 9569 2746
rect 9593 2694 9603 2746
rect 9603 2694 9649 2746
rect 9353 2692 9409 2694
rect 9433 2692 9489 2694
rect 9513 2692 9569 2694
rect 9593 2692 9649 2694
rect 18234 21836 18236 21856
rect 18236 21836 18288 21856
rect 18288 21836 18290 21856
rect 18234 21800 18290 21836
rect 17750 21786 17806 21788
rect 17830 21786 17886 21788
rect 17910 21786 17966 21788
rect 17990 21786 18046 21788
rect 17750 21734 17796 21786
rect 17796 21734 17806 21786
rect 17830 21734 17860 21786
rect 17860 21734 17872 21786
rect 17872 21734 17886 21786
rect 17910 21734 17924 21786
rect 17924 21734 17936 21786
rect 17936 21734 17966 21786
rect 17990 21734 18000 21786
rect 18000 21734 18046 21786
rect 17750 21732 17806 21734
rect 17830 21732 17886 21734
rect 17910 21732 17966 21734
rect 17990 21732 18046 21734
rect 18142 21664 18198 21720
rect 17750 20698 17806 20700
rect 17830 20698 17886 20700
rect 17910 20698 17966 20700
rect 17990 20698 18046 20700
rect 17750 20646 17796 20698
rect 17796 20646 17806 20698
rect 17830 20646 17860 20698
rect 17860 20646 17872 20698
rect 17872 20646 17886 20698
rect 17910 20646 17924 20698
rect 17924 20646 17936 20698
rect 17936 20646 17966 20698
rect 17990 20646 18000 20698
rect 18000 20646 18046 20698
rect 17750 20644 17806 20646
rect 17830 20644 17886 20646
rect 17910 20644 17966 20646
rect 17990 20644 18046 20646
rect 17682 20440 17738 20496
rect 17866 20476 17868 20496
rect 17868 20476 17920 20496
rect 17920 20476 17922 20496
rect 17866 20440 17922 20476
rect 17958 20168 18014 20224
rect 17222 19352 17278 19408
rect 16946 18128 17002 18184
rect 17958 19780 18014 19816
rect 17958 19760 17960 19780
rect 17960 19760 18012 19780
rect 18012 19760 18014 19780
rect 17750 19610 17806 19612
rect 17830 19610 17886 19612
rect 17910 19610 17966 19612
rect 17990 19610 18046 19612
rect 17750 19558 17796 19610
rect 17796 19558 17806 19610
rect 17830 19558 17860 19610
rect 17860 19558 17872 19610
rect 17872 19558 17886 19610
rect 17910 19558 17924 19610
rect 17924 19558 17936 19610
rect 17936 19558 17966 19610
rect 17990 19558 18000 19610
rect 18000 19558 18046 19610
rect 17750 19556 17806 19558
rect 17830 19556 17886 19558
rect 17910 19556 17966 19558
rect 17990 19556 18046 19558
rect 18418 20848 18474 20904
rect 18326 20576 18382 20632
rect 18326 20304 18382 20360
rect 18326 19508 18382 19544
rect 18326 19488 18328 19508
rect 18328 19488 18380 19508
rect 18380 19488 18382 19508
rect 17406 17484 17408 17504
rect 17408 17484 17460 17504
rect 17460 17484 17462 17504
rect 17406 17448 17462 17484
rect 17750 18522 17806 18524
rect 17830 18522 17886 18524
rect 17910 18522 17966 18524
rect 17990 18522 18046 18524
rect 17750 18470 17796 18522
rect 17796 18470 17806 18522
rect 17830 18470 17860 18522
rect 17860 18470 17872 18522
rect 17872 18470 17886 18522
rect 17910 18470 17924 18522
rect 17924 18470 17936 18522
rect 17936 18470 17966 18522
rect 17990 18470 18000 18522
rect 18000 18470 18046 18522
rect 17750 18468 17806 18470
rect 17830 18468 17886 18470
rect 17910 18468 17966 18470
rect 17990 18468 18046 18470
rect 17750 17434 17806 17436
rect 17830 17434 17886 17436
rect 17910 17434 17966 17436
rect 17990 17434 18046 17436
rect 17750 17382 17796 17434
rect 17796 17382 17806 17434
rect 17830 17382 17860 17434
rect 17860 17382 17872 17434
rect 17872 17382 17886 17434
rect 17910 17382 17924 17434
rect 17924 17382 17936 17434
rect 17936 17382 17966 17434
rect 17990 17382 18000 17434
rect 18000 17382 18046 17434
rect 17750 17380 17806 17382
rect 17830 17380 17886 17382
rect 17910 17380 17966 17382
rect 17990 17380 18046 17382
rect 17750 16346 17806 16348
rect 17830 16346 17886 16348
rect 17910 16346 17966 16348
rect 17990 16346 18046 16348
rect 17750 16294 17796 16346
rect 17796 16294 17806 16346
rect 17830 16294 17860 16346
rect 17860 16294 17872 16346
rect 17872 16294 17886 16346
rect 17910 16294 17924 16346
rect 17924 16294 17936 16346
rect 17936 16294 17966 16346
rect 17990 16294 18000 16346
rect 18000 16294 18046 16346
rect 17750 16292 17806 16294
rect 17830 16292 17886 16294
rect 17910 16292 17966 16294
rect 17990 16292 18046 16294
rect 18878 20168 18934 20224
rect 20549 22330 20605 22332
rect 20629 22330 20685 22332
rect 20709 22330 20765 22332
rect 20789 22330 20845 22332
rect 20549 22278 20595 22330
rect 20595 22278 20605 22330
rect 20629 22278 20659 22330
rect 20659 22278 20671 22330
rect 20671 22278 20685 22330
rect 20709 22278 20723 22330
rect 20723 22278 20735 22330
rect 20735 22278 20765 22330
rect 20789 22278 20799 22330
rect 20799 22278 20845 22330
rect 20549 22276 20605 22278
rect 20629 22276 20685 22278
rect 20709 22276 20765 22278
rect 20789 22276 20845 22278
rect 20810 22108 20812 22128
rect 20812 22108 20864 22128
rect 20864 22108 20866 22128
rect 19246 21664 19302 21720
rect 19430 21528 19486 21584
rect 19246 21256 19302 21312
rect 19062 20576 19118 20632
rect 19246 20848 19302 20904
rect 19246 19760 19302 19816
rect 19614 20576 19670 20632
rect 19430 19624 19486 19680
rect 19430 19488 19486 19544
rect 18786 17584 18842 17640
rect 17222 15544 17278 15600
rect 17590 15544 17646 15600
rect 17750 15258 17806 15260
rect 17830 15258 17886 15260
rect 17910 15258 17966 15260
rect 17990 15258 18046 15260
rect 17750 15206 17796 15258
rect 17796 15206 17806 15258
rect 17830 15206 17860 15258
rect 17860 15206 17872 15258
rect 17872 15206 17886 15258
rect 17910 15206 17924 15258
rect 17924 15206 17936 15258
rect 17936 15206 17966 15258
rect 17990 15206 18000 15258
rect 18000 15206 18046 15258
rect 17750 15204 17806 15206
rect 17830 15204 17886 15206
rect 17910 15204 17966 15206
rect 17990 15204 18046 15206
rect 17750 14170 17806 14172
rect 17830 14170 17886 14172
rect 17910 14170 17966 14172
rect 17990 14170 18046 14172
rect 17750 14118 17796 14170
rect 17796 14118 17806 14170
rect 17830 14118 17860 14170
rect 17860 14118 17872 14170
rect 17872 14118 17886 14170
rect 17910 14118 17924 14170
rect 17924 14118 17936 14170
rect 17936 14118 17966 14170
rect 17990 14118 18000 14170
rect 18000 14118 18046 14170
rect 17750 14116 17806 14118
rect 17830 14116 17886 14118
rect 17910 14116 17966 14118
rect 17990 14116 18046 14118
rect 19338 16632 19394 16688
rect 19706 18536 19762 18592
rect 18694 16224 18750 16280
rect 18786 15136 18842 15192
rect 19338 15000 19394 15056
rect 20074 21528 20130 21584
rect 20074 21120 20130 21176
rect 20810 22072 20866 22108
rect 20549 21242 20605 21244
rect 20629 21242 20685 21244
rect 20709 21242 20765 21244
rect 20789 21242 20845 21244
rect 20549 21190 20595 21242
rect 20595 21190 20605 21242
rect 20629 21190 20659 21242
rect 20659 21190 20671 21242
rect 20671 21190 20685 21242
rect 20709 21190 20723 21242
rect 20723 21190 20735 21242
rect 20735 21190 20765 21242
rect 20789 21190 20799 21242
rect 20799 21190 20845 21242
rect 20549 21188 20605 21190
rect 20629 21188 20685 21190
rect 20709 21188 20765 21190
rect 20789 21188 20845 21190
rect 21086 20984 21142 21040
rect 20549 20154 20605 20156
rect 20629 20154 20685 20156
rect 20709 20154 20765 20156
rect 20789 20154 20845 20156
rect 20549 20102 20595 20154
rect 20595 20102 20605 20154
rect 20629 20102 20659 20154
rect 20659 20102 20671 20154
rect 20671 20102 20685 20154
rect 20709 20102 20723 20154
rect 20723 20102 20735 20154
rect 20735 20102 20765 20154
rect 20789 20102 20799 20154
rect 20799 20102 20845 20154
rect 20549 20100 20605 20102
rect 20629 20100 20685 20102
rect 20709 20100 20765 20102
rect 20789 20100 20845 20102
rect 20718 19796 20720 19816
rect 20720 19796 20772 19816
rect 20772 19796 20774 19816
rect 20718 19760 20774 19796
rect 21086 19624 21142 19680
rect 20994 19488 21050 19544
rect 20549 19066 20605 19068
rect 20629 19066 20685 19068
rect 20709 19066 20765 19068
rect 20789 19066 20845 19068
rect 20549 19014 20595 19066
rect 20595 19014 20605 19066
rect 20629 19014 20659 19066
rect 20659 19014 20671 19066
rect 20671 19014 20685 19066
rect 20709 19014 20723 19066
rect 20723 19014 20735 19066
rect 20735 19014 20765 19066
rect 20789 19014 20799 19066
rect 20799 19014 20845 19066
rect 20549 19012 20605 19014
rect 20629 19012 20685 19014
rect 20709 19012 20765 19014
rect 20789 19012 20845 19014
rect 20810 18128 20866 18184
rect 19706 15544 19762 15600
rect 17750 13082 17806 13084
rect 17830 13082 17886 13084
rect 17910 13082 17966 13084
rect 17990 13082 18046 13084
rect 17750 13030 17796 13082
rect 17796 13030 17806 13082
rect 17830 13030 17860 13082
rect 17860 13030 17872 13082
rect 17872 13030 17886 13082
rect 17910 13030 17924 13082
rect 17924 13030 17936 13082
rect 17936 13030 17966 13082
rect 17990 13030 18000 13082
rect 18000 13030 18046 13082
rect 17750 13028 17806 13030
rect 17830 13028 17886 13030
rect 17910 13028 17966 13030
rect 17990 13028 18046 13030
rect 18326 12980 18382 13016
rect 18326 12960 18328 12980
rect 18328 12960 18380 12980
rect 18380 12960 18382 12980
rect 17958 12144 18014 12200
rect 17750 11994 17806 11996
rect 17830 11994 17886 11996
rect 17910 11994 17966 11996
rect 17990 11994 18046 11996
rect 17750 11942 17796 11994
rect 17796 11942 17806 11994
rect 17830 11942 17860 11994
rect 17860 11942 17872 11994
rect 17872 11942 17886 11994
rect 17910 11942 17924 11994
rect 17924 11942 17936 11994
rect 17936 11942 17966 11994
rect 17990 11942 18000 11994
rect 18000 11942 18046 11994
rect 17750 11940 17806 11942
rect 17830 11940 17886 11942
rect 17910 11940 17966 11942
rect 17990 11940 18046 11942
rect 18326 11756 18382 11792
rect 18326 11736 18328 11756
rect 18328 11736 18380 11756
rect 18380 11736 18382 11756
rect 18142 11192 18198 11248
rect 18050 11056 18106 11112
rect 16946 9968 17002 10024
rect 17130 8880 17186 8936
rect 15934 8356 15990 8392
rect 15934 8336 15936 8356
rect 15936 8336 15988 8356
rect 15988 8336 15990 8356
rect 15842 6296 15898 6352
rect 16026 6296 16082 6352
rect 16302 5752 16358 5808
rect 16670 4020 16672 4040
rect 16672 4020 16724 4040
rect 16724 4020 16726 4040
rect 16670 3984 16726 4020
rect 17314 8336 17370 8392
rect 17750 10906 17806 10908
rect 17830 10906 17886 10908
rect 17910 10906 17966 10908
rect 17990 10906 18046 10908
rect 17750 10854 17796 10906
rect 17796 10854 17806 10906
rect 17830 10854 17860 10906
rect 17860 10854 17872 10906
rect 17872 10854 17886 10906
rect 17910 10854 17924 10906
rect 17924 10854 17936 10906
rect 17936 10854 17966 10906
rect 17990 10854 18000 10906
rect 18000 10854 18046 10906
rect 17750 10852 17806 10854
rect 17830 10852 17886 10854
rect 17910 10852 17966 10854
rect 17990 10852 18046 10854
rect 17750 9818 17806 9820
rect 17830 9818 17886 9820
rect 17910 9818 17966 9820
rect 17990 9818 18046 9820
rect 17750 9766 17796 9818
rect 17796 9766 17806 9818
rect 17830 9766 17860 9818
rect 17860 9766 17872 9818
rect 17872 9766 17886 9818
rect 17910 9766 17924 9818
rect 17924 9766 17936 9818
rect 17936 9766 17966 9818
rect 17990 9766 18000 9818
rect 18000 9766 18046 9818
rect 17750 9764 17806 9766
rect 17830 9764 17886 9766
rect 17910 9764 17966 9766
rect 17990 9764 18046 9766
rect 18326 9696 18382 9752
rect 17774 9580 17830 9616
rect 17774 9560 17776 9580
rect 17776 9560 17828 9580
rect 17828 9560 17830 9580
rect 17590 9424 17646 9480
rect 17750 8730 17806 8732
rect 17830 8730 17886 8732
rect 17910 8730 17966 8732
rect 17990 8730 18046 8732
rect 17750 8678 17796 8730
rect 17796 8678 17806 8730
rect 17830 8678 17860 8730
rect 17860 8678 17872 8730
rect 17872 8678 17886 8730
rect 17910 8678 17924 8730
rect 17924 8678 17936 8730
rect 17936 8678 17966 8730
rect 17990 8678 18000 8730
rect 18000 8678 18046 8730
rect 17750 8676 17806 8678
rect 17830 8676 17886 8678
rect 17910 8676 17966 8678
rect 17990 8676 18046 8678
rect 17750 7642 17806 7644
rect 17830 7642 17886 7644
rect 17910 7642 17966 7644
rect 17990 7642 18046 7644
rect 17750 7590 17796 7642
rect 17796 7590 17806 7642
rect 17830 7590 17860 7642
rect 17860 7590 17872 7642
rect 17872 7590 17886 7642
rect 17910 7590 17924 7642
rect 17924 7590 17936 7642
rect 17936 7590 17966 7642
rect 17990 7590 18000 7642
rect 18000 7590 18046 7642
rect 17750 7588 17806 7590
rect 17830 7588 17886 7590
rect 17910 7588 17966 7590
rect 17990 7588 18046 7590
rect 18326 7928 18382 7984
rect 18142 7268 18198 7304
rect 18142 7248 18144 7268
rect 18144 7248 18196 7268
rect 18196 7248 18198 7268
rect 18142 6568 18198 6624
rect 17750 6554 17806 6556
rect 17830 6554 17886 6556
rect 17910 6554 17966 6556
rect 17990 6554 18046 6556
rect 17750 6502 17796 6554
rect 17796 6502 17806 6554
rect 17830 6502 17860 6554
rect 17860 6502 17872 6554
rect 17872 6502 17886 6554
rect 17910 6502 17924 6554
rect 17924 6502 17936 6554
rect 17936 6502 17966 6554
rect 17990 6502 18000 6554
rect 18000 6502 18046 6554
rect 17750 6500 17806 6502
rect 17830 6500 17886 6502
rect 17910 6500 17966 6502
rect 17990 6500 18046 6502
rect 17750 5466 17806 5468
rect 17830 5466 17886 5468
rect 17910 5466 17966 5468
rect 17990 5466 18046 5468
rect 17750 5414 17796 5466
rect 17796 5414 17806 5466
rect 17830 5414 17860 5466
rect 17860 5414 17872 5466
rect 17872 5414 17886 5466
rect 17910 5414 17924 5466
rect 17924 5414 17936 5466
rect 17936 5414 17966 5466
rect 17990 5414 18000 5466
rect 18000 5414 18046 5466
rect 17750 5412 17806 5414
rect 17830 5412 17886 5414
rect 17910 5412 17966 5414
rect 17990 5412 18046 5414
rect 17750 4378 17806 4380
rect 17830 4378 17886 4380
rect 17910 4378 17966 4380
rect 17990 4378 18046 4380
rect 17750 4326 17796 4378
rect 17796 4326 17806 4378
rect 17830 4326 17860 4378
rect 17860 4326 17872 4378
rect 17872 4326 17886 4378
rect 17910 4326 17924 4378
rect 17924 4326 17936 4378
rect 17936 4326 17966 4378
rect 17990 4326 18000 4378
rect 18000 4326 18046 4378
rect 17750 4324 17806 4326
rect 17830 4324 17886 4326
rect 17910 4324 17966 4326
rect 17990 4324 18046 4326
rect 19338 13368 19394 13424
rect 19430 13096 19486 13152
rect 19062 12824 19118 12880
rect 19062 12688 19118 12744
rect 19338 12280 19394 12336
rect 19338 11228 19340 11248
rect 19340 11228 19392 11248
rect 19392 11228 19394 11248
rect 18510 7520 18566 7576
rect 19338 11192 19394 11228
rect 19338 10784 19394 10840
rect 19246 10104 19302 10160
rect 19798 14864 19854 14920
rect 19706 13912 19762 13968
rect 19798 11872 19854 11928
rect 19338 9832 19394 9888
rect 19706 9696 19762 9752
rect 19338 9016 19394 9072
rect 19154 8744 19210 8800
rect 19338 8472 19394 8528
rect 19062 7112 19118 7168
rect 19154 6976 19210 7032
rect 19522 8628 19578 8664
rect 19522 8608 19524 8628
rect 19524 8608 19576 8628
rect 19576 8608 19578 8628
rect 19338 7112 19394 7168
rect 18970 6060 18972 6080
rect 18972 6060 19024 6080
rect 19024 6060 19026 6080
rect 18970 6024 19026 6060
rect 19062 5888 19118 5944
rect 19430 6432 19486 6488
rect 19338 5344 19394 5400
rect 19246 4120 19302 4176
rect 18510 3340 18512 3360
rect 18512 3340 18564 3360
rect 18564 3340 18566 3360
rect 18510 3304 18566 3340
rect 17750 3290 17806 3292
rect 17830 3290 17886 3292
rect 17910 3290 17966 3292
rect 17990 3290 18046 3292
rect 17750 3238 17796 3290
rect 17796 3238 17806 3290
rect 17830 3238 17860 3290
rect 17860 3238 17872 3290
rect 17872 3238 17886 3290
rect 17910 3238 17924 3290
rect 17924 3238 17936 3290
rect 17936 3238 17966 3290
rect 17990 3238 18000 3290
rect 18000 3238 18046 3290
rect 17750 3236 17806 3238
rect 17830 3236 17886 3238
rect 17910 3236 17966 3238
rect 17990 3236 18046 3238
rect 14951 2746 15007 2748
rect 15031 2746 15087 2748
rect 15111 2746 15167 2748
rect 15191 2746 15247 2748
rect 14951 2694 14997 2746
rect 14997 2694 15007 2746
rect 15031 2694 15061 2746
rect 15061 2694 15073 2746
rect 15073 2694 15087 2746
rect 15111 2694 15125 2746
rect 15125 2694 15137 2746
rect 15137 2694 15167 2746
rect 15191 2694 15201 2746
rect 15201 2694 15247 2746
rect 14951 2692 15007 2694
rect 15031 2692 15087 2694
rect 15111 2692 15167 2694
rect 15191 2692 15247 2694
rect 20549 17978 20605 17980
rect 20629 17978 20685 17980
rect 20709 17978 20765 17980
rect 20789 17978 20845 17980
rect 20549 17926 20595 17978
rect 20595 17926 20605 17978
rect 20629 17926 20659 17978
rect 20659 17926 20671 17978
rect 20671 17926 20685 17978
rect 20709 17926 20723 17978
rect 20723 17926 20735 17978
rect 20735 17926 20765 17978
rect 20789 17926 20799 17978
rect 20799 17926 20845 17978
rect 20549 17924 20605 17926
rect 20629 17924 20685 17926
rect 20709 17924 20765 17926
rect 20789 17924 20845 17926
rect 20549 16890 20605 16892
rect 20629 16890 20685 16892
rect 20709 16890 20765 16892
rect 20789 16890 20845 16892
rect 20549 16838 20595 16890
rect 20595 16838 20605 16890
rect 20629 16838 20659 16890
rect 20659 16838 20671 16890
rect 20671 16838 20685 16890
rect 20709 16838 20723 16890
rect 20723 16838 20735 16890
rect 20735 16838 20765 16890
rect 20789 16838 20799 16890
rect 20799 16838 20845 16890
rect 20549 16836 20605 16838
rect 20629 16836 20685 16838
rect 20709 16836 20765 16838
rect 20789 16836 20845 16838
rect 21086 16496 21142 16552
rect 20626 16360 20682 16416
rect 21362 21392 21418 21448
rect 21362 20460 21418 20496
rect 21362 20440 21364 20460
rect 21364 20440 21416 20460
rect 21416 20440 21418 20460
rect 21546 20596 21602 20632
rect 21546 20576 21548 20596
rect 21548 20576 21600 20596
rect 21600 20576 21602 20596
rect 21270 19372 21326 19408
rect 21270 19352 21272 19372
rect 21272 19352 21324 19372
rect 21324 19352 21326 19372
rect 22374 22072 22430 22128
rect 21822 21972 21824 21992
rect 21824 21972 21876 21992
rect 21876 21972 21878 21992
rect 21822 21936 21878 21972
rect 22098 20848 22154 20904
rect 22558 21800 22614 21856
rect 22466 21548 22522 21584
rect 22466 21528 22468 21548
rect 22468 21528 22520 21548
rect 22520 21528 22522 21548
rect 22650 21528 22706 21584
rect 21178 16224 21234 16280
rect 21362 16224 21418 16280
rect 21086 16088 21142 16144
rect 21270 16108 21326 16144
rect 21270 16088 21272 16108
rect 21272 16088 21324 16108
rect 21324 16088 21326 16108
rect 20549 15802 20605 15804
rect 20629 15802 20685 15804
rect 20709 15802 20765 15804
rect 20789 15802 20845 15804
rect 20549 15750 20595 15802
rect 20595 15750 20605 15802
rect 20629 15750 20659 15802
rect 20659 15750 20671 15802
rect 20671 15750 20685 15802
rect 20709 15750 20723 15802
rect 20723 15750 20735 15802
rect 20735 15750 20765 15802
rect 20789 15750 20799 15802
rect 20799 15750 20845 15802
rect 20549 15748 20605 15750
rect 20629 15748 20685 15750
rect 20709 15748 20765 15750
rect 20789 15748 20845 15750
rect 20549 14714 20605 14716
rect 20629 14714 20685 14716
rect 20709 14714 20765 14716
rect 20789 14714 20845 14716
rect 20549 14662 20595 14714
rect 20595 14662 20605 14714
rect 20629 14662 20659 14714
rect 20659 14662 20671 14714
rect 20671 14662 20685 14714
rect 20709 14662 20723 14714
rect 20723 14662 20735 14714
rect 20735 14662 20765 14714
rect 20789 14662 20799 14714
rect 20799 14662 20845 14714
rect 20549 14660 20605 14662
rect 20629 14660 20685 14662
rect 20709 14660 20765 14662
rect 20789 14660 20845 14662
rect 20258 14456 20314 14512
rect 21822 17720 21878 17776
rect 21546 16496 21602 16552
rect 21822 17448 21878 17504
rect 23018 20984 23074 21040
rect 23018 20440 23074 20496
rect 22282 18672 22338 18728
rect 22374 18264 22430 18320
rect 22190 17584 22246 17640
rect 22374 16396 22376 16416
rect 22376 16396 22428 16416
rect 22428 16396 22430 16416
rect 22374 16360 22430 16396
rect 22374 16224 22430 16280
rect 22834 19896 22890 19952
rect 22742 17584 22798 17640
rect 22650 17176 22706 17232
rect 22742 17040 22798 17096
rect 21546 15136 21602 15192
rect 21730 15020 21786 15056
rect 21730 15000 21732 15020
rect 21732 15000 21784 15020
rect 21784 15000 21786 15020
rect 20549 13626 20605 13628
rect 20629 13626 20685 13628
rect 20709 13626 20765 13628
rect 20789 13626 20845 13628
rect 20549 13574 20595 13626
rect 20595 13574 20605 13626
rect 20629 13574 20659 13626
rect 20659 13574 20671 13626
rect 20671 13574 20685 13626
rect 20709 13574 20723 13626
rect 20723 13574 20735 13626
rect 20735 13574 20765 13626
rect 20789 13574 20799 13626
rect 20799 13574 20845 13626
rect 20549 13572 20605 13574
rect 20629 13572 20685 13574
rect 20709 13572 20765 13574
rect 20789 13572 20845 13574
rect 21362 14320 21418 14376
rect 21086 13252 21142 13288
rect 21086 13232 21088 13252
rect 21088 13232 21140 13252
rect 21140 13232 21142 13252
rect 21086 12960 21142 13016
rect 19982 11600 20038 11656
rect 20549 12538 20605 12540
rect 20629 12538 20685 12540
rect 20709 12538 20765 12540
rect 20789 12538 20845 12540
rect 20549 12486 20595 12538
rect 20595 12486 20605 12538
rect 20629 12486 20659 12538
rect 20659 12486 20671 12538
rect 20671 12486 20685 12538
rect 20709 12486 20723 12538
rect 20723 12486 20735 12538
rect 20735 12486 20765 12538
rect 20789 12486 20799 12538
rect 20799 12486 20845 12538
rect 20549 12484 20605 12486
rect 20629 12484 20685 12486
rect 20709 12484 20765 12486
rect 20789 12484 20845 12486
rect 20994 12008 21050 12064
rect 21178 12824 21234 12880
rect 20549 11450 20605 11452
rect 20629 11450 20685 11452
rect 20709 11450 20765 11452
rect 20789 11450 20845 11452
rect 20549 11398 20595 11450
rect 20595 11398 20605 11450
rect 20629 11398 20659 11450
rect 20659 11398 20671 11450
rect 20671 11398 20685 11450
rect 20709 11398 20723 11450
rect 20723 11398 20735 11450
rect 20735 11398 20765 11450
rect 20789 11398 20799 11450
rect 20799 11398 20845 11450
rect 20549 11396 20605 11398
rect 20629 11396 20685 11398
rect 20709 11396 20765 11398
rect 20789 11396 20845 11398
rect 20902 11056 20958 11112
rect 20549 10362 20605 10364
rect 20629 10362 20685 10364
rect 20709 10362 20765 10364
rect 20789 10362 20845 10364
rect 20549 10310 20595 10362
rect 20595 10310 20605 10362
rect 20629 10310 20659 10362
rect 20659 10310 20671 10362
rect 20671 10310 20685 10362
rect 20709 10310 20723 10362
rect 20723 10310 20735 10362
rect 20735 10310 20765 10362
rect 20789 10310 20799 10362
rect 20799 10310 20845 10362
rect 20549 10308 20605 10310
rect 20629 10308 20685 10310
rect 20709 10308 20765 10310
rect 20789 10308 20845 10310
rect 20718 10140 20720 10160
rect 20720 10140 20772 10160
rect 20772 10140 20774 10160
rect 20718 10104 20774 10140
rect 19890 7656 19946 7712
rect 19706 7384 19762 7440
rect 19614 7112 19670 7168
rect 19706 5616 19762 5672
rect 19522 3576 19578 3632
rect 19522 2916 19578 2952
rect 19522 2896 19524 2916
rect 19524 2896 19576 2916
rect 19576 2896 19578 2916
rect 20166 8472 20222 8528
rect 20074 7792 20130 7848
rect 19982 6160 20038 6216
rect 20549 9274 20605 9276
rect 20629 9274 20685 9276
rect 20709 9274 20765 9276
rect 20789 9274 20845 9276
rect 20549 9222 20595 9274
rect 20595 9222 20605 9274
rect 20629 9222 20659 9274
rect 20659 9222 20671 9274
rect 20671 9222 20685 9274
rect 20709 9222 20723 9274
rect 20723 9222 20735 9274
rect 20735 9222 20765 9274
rect 20789 9222 20799 9274
rect 20799 9222 20845 9274
rect 20549 9220 20605 9222
rect 20629 9220 20685 9222
rect 20709 9220 20765 9222
rect 20789 9220 20845 9222
rect 20258 6296 20314 6352
rect 20074 5516 20076 5536
rect 20076 5516 20128 5536
rect 20128 5516 20130 5536
rect 20074 5480 20130 5516
rect 20074 5208 20130 5264
rect 20258 4548 20314 4584
rect 20258 4528 20260 4548
rect 20260 4528 20312 4548
rect 20312 4528 20314 4548
rect 20534 8472 20590 8528
rect 20549 8186 20605 8188
rect 20629 8186 20685 8188
rect 20709 8186 20765 8188
rect 20789 8186 20845 8188
rect 20549 8134 20595 8186
rect 20595 8134 20605 8186
rect 20629 8134 20659 8186
rect 20659 8134 20671 8186
rect 20671 8134 20685 8186
rect 20709 8134 20723 8186
rect 20723 8134 20735 8186
rect 20735 8134 20765 8186
rect 20789 8134 20799 8186
rect 20799 8134 20845 8186
rect 20549 8132 20605 8134
rect 20629 8132 20685 8134
rect 20709 8132 20765 8134
rect 20789 8132 20845 8134
rect 20442 7656 20498 7712
rect 20810 7656 20866 7712
rect 20549 7098 20605 7100
rect 20629 7098 20685 7100
rect 20709 7098 20765 7100
rect 20789 7098 20845 7100
rect 20549 7046 20595 7098
rect 20595 7046 20605 7098
rect 20629 7046 20659 7098
rect 20659 7046 20671 7098
rect 20671 7046 20685 7098
rect 20709 7046 20723 7098
rect 20723 7046 20735 7098
rect 20735 7046 20765 7098
rect 20789 7046 20799 7098
rect 20799 7046 20845 7098
rect 20549 7044 20605 7046
rect 20629 7044 20685 7046
rect 20709 7044 20765 7046
rect 20789 7044 20845 7046
rect 20994 9560 21050 9616
rect 20994 9288 21050 9344
rect 21270 12688 21326 12744
rect 21730 13912 21786 13968
rect 21638 11600 21694 11656
rect 21914 10104 21970 10160
rect 21270 9560 21326 9616
rect 22098 10684 22100 10704
rect 22100 10684 22152 10704
rect 22152 10684 22154 10704
rect 22098 10648 22154 10684
rect 21822 8900 21878 8936
rect 21822 8880 21824 8900
rect 21824 8880 21876 8900
rect 21876 8880 21878 8900
rect 20442 6432 20498 6488
rect 20626 6432 20682 6488
rect 20902 6740 20904 6760
rect 20904 6740 20956 6760
rect 20956 6740 20958 6760
rect 20902 6704 20958 6740
rect 20902 6568 20958 6624
rect 20549 6010 20605 6012
rect 20629 6010 20685 6012
rect 20709 6010 20765 6012
rect 20789 6010 20845 6012
rect 20549 5958 20595 6010
rect 20595 5958 20605 6010
rect 20629 5958 20659 6010
rect 20659 5958 20671 6010
rect 20671 5958 20685 6010
rect 20709 5958 20723 6010
rect 20723 5958 20735 6010
rect 20735 5958 20765 6010
rect 20789 5958 20799 6010
rect 20799 5958 20845 6010
rect 20549 5956 20605 5958
rect 20629 5956 20685 5958
rect 20709 5956 20765 5958
rect 20789 5956 20845 5958
rect 20534 5344 20590 5400
rect 20549 4922 20605 4924
rect 20629 4922 20685 4924
rect 20709 4922 20765 4924
rect 20789 4922 20845 4924
rect 20549 4870 20595 4922
rect 20595 4870 20605 4922
rect 20629 4870 20659 4922
rect 20659 4870 20671 4922
rect 20671 4870 20685 4922
rect 20709 4870 20723 4922
rect 20723 4870 20735 4922
rect 20735 4870 20765 4922
rect 20789 4870 20799 4922
rect 20799 4870 20845 4922
rect 20549 4868 20605 4870
rect 20629 4868 20685 4870
rect 20709 4868 20765 4870
rect 20789 4868 20845 4870
rect 20810 4664 20866 4720
rect 20549 3834 20605 3836
rect 20629 3834 20685 3836
rect 20709 3834 20765 3836
rect 20789 3834 20845 3836
rect 20549 3782 20595 3834
rect 20595 3782 20605 3834
rect 20629 3782 20659 3834
rect 20659 3782 20671 3834
rect 20671 3782 20685 3834
rect 20709 3782 20723 3834
rect 20723 3782 20735 3834
rect 20735 3782 20765 3834
rect 20789 3782 20799 3834
rect 20799 3782 20845 3834
rect 20549 3780 20605 3782
rect 20629 3780 20685 3782
rect 20709 3780 20765 3782
rect 20789 3780 20845 3782
rect 21178 5344 21234 5400
rect 21178 5072 21234 5128
rect 20549 2746 20605 2748
rect 20629 2746 20685 2748
rect 20709 2746 20765 2748
rect 20789 2746 20845 2748
rect 20549 2694 20595 2746
rect 20595 2694 20605 2746
rect 20629 2694 20659 2746
rect 20659 2694 20671 2746
rect 20671 2694 20685 2746
rect 20709 2694 20723 2746
rect 20723 2694 20735 2746
rect 20735 2694 20765 2746
rect 20789 2694 20799 2746
rect 20799 2694 20845 2746
rect 20549 2692 20605 2694
rect 20629 2692 20685 2694
rect 20709 2692 20765 2694
rect 20789 2692 20845 2694
rect 21454 7384 21510 7440
rect 21822 7928 21878 7984
rect 22006 7928 22062 7984
rect 21454 7148 21456 7168
rect 21456 7148 21508 7168
rect 21508 7148 21510 7168
rect 21454 7112 21510 7148
rect 21546 6296 21602 6352
rect 22098 7792 22154 7848
rect 21822 6568 21878 6624
rect 21730 5752 21786 5808
rect 21270 3984 21326 4040
rect 21546 3576 21602 3632
rect 21914 5888 21970 5944
rect 21730 2896 21786 2952
rect 22282 6976 22338 7032
rect 22190 6568 22246 6624
rect 22282 6332 22284 6352
rect 22284 6332 22336 6352
rect 22336 6332 22338 6352
rect 22282 6296 22338 6332
rect 22190 6160 22246 6216
rect 22098 6024 22154 6080
rect 23110 19896 23166 19952
rect 23110 19252 23112 19272
rect 23112 19252 23164 19272
rect 23164 19252 23166 19272
rect 23110 19216 23166 19252
rect 23018 18808 23074 18864
rect 23294 19352 23350 19408
rect 23202 18536 23258 18592
rect 23110 18264 23166 18320
rect 23110 17176 23166 17232
rect 22926 15000 22982 15056
rect 23202 14456 23258 14512
rect 22650 12144 22706 12200
rect 22742 12044 22744 12064
rect 22744 12044 22796 12064
rect 22796 12044 22798 12064
rect 22742 12008 22798 12044
rect 22834 11872 22890 11928
rect 22834 9968 22890 10024
rect 22742 9560 22798 9616
rect 22558 9424 22614 9480
rect 22834 7520 22890 7576
rect 23662 15952 23718 16008
rect 23570 15408 23626 15464
rect 22742 7248 22798 7304
rect 22650 6840 22706 6896
rect 22466 6296 22522 6352
rect 22374 6024 22430 6080
rect 22558 5616 22614 5672
rect 22466 5480 22522 5536
rect 22650 5364 22706 5400
rect 22650 5344 22652 5364
rect 22652 5344 22704 5364
rect 22704 5344 22706 5364
rect 22650 5208 22706 5264
rect 22558 4120 22614 4176
rect 23110 8492 23166 8528
rect 23110 8472 23112 8492
rect 23112 8472 23164 8492
rect 23164 8472 23166 8492
rect 22834 5752 22890 5808
rect 23110 6840 23166 6896
rect 23018 6296 23074 6352
rect 23294 8608 23350 8664
rect 23202 5752 23258 5808
rect 22466 3304 22522 3360
rect 22742 3712 22798 3768
rect 23110 5480 23166 5536
rect 22926 5208 22982 5264
rect 23018 4664 23074 4720
rect 23110 4120 23166 4176
rect 23662 8336 23718 8392
rect 23018 3032 23074 3088
rect 22650 2488 22706 2544
rect 6554 2202 6610 2204
rect 6634 2202 6690 2204
rect 6714 2202 6770 2204
rect 6794 2202 6850 2204
rect 6554 2150 6600 2202
rect 6600 2150 6610 2202
rect 6634 2150 6664 2202
rect 6664 2150 6676 2202
rect 6676 2150 6690 2202
rect 6714 2150 6728 2202
rect 6728 2150 6740 2202
rect 6740 2150 6770 2202
rect 6794 2150 6804 2202
rect 6804 2150 6850 2202
rect 6554 2148 6610 2150
rect 6634 2148 6690 2150
rect 6714 2148 6770 2150
rect 6794 2148 6850 2150
rect 12152 2202 12208 2204
rect 12232 2202 12288 2204
rect 12312 2202 12368 2204
rect 12392 2202 12448 2204
rect 12152 2150 12198 2202
rect 12198 2150 12208 2202
rect 12232 2150 12262 2202
rect 12262 2150 12274 2202
rect 12274 2150 12288 2202
rect 12312 2150 12326 2202
rect 12326 2150 12338 2202
rect 12338 2150 12368 2202
rect 12392 2150 12402 2202
rect 12402 2150 12448 2202
rect 12152 2148 12208 2150
rect 12232 2148 12288 2150
rect 12312 2148 12368 2150
rect 12392 2148 12448 2150
rect 17750 2202 17806 2204
rect 17830 2202 17886 2204
rect 17910 2202 17966 2204
rect 17990 2202 18046 2204
rect 17750 2150 17796 2202
rect 17796 2150 17806 2202
rect 17830 2150 17860 2202
rect 17860 2150 17872 2202
rect 17872 2150 17886 2202
rect 17910 2150 17924 2202
rect 17924 2150 17936 2202
rect 17936 2150 17966 2202
rect 17990 2150 18000 2202
rect 18000 2150 18046 2202
rect 17750 2148 17806 2150
rect 17830 2148 17886 2150
rect 17910 2148 17966 2150
rect 17990 2148 18046 2150
<< metal3 >>
rect 3325 22538 3391 22541
rect 18229 22538 18295 22541
rect 3325 22536 18295 22538
rect 3325 22480 3330 22536
rect 3386 22480 18234 22536
rect 18290 22480 18295 22536
rect 3325 22478 18295 22480
rect 3325 22475 3391 22478
rect 18229 22475 18295 22478
rect 5349 22402 5415 22405
rect 8753 22402 8819 22405
rect 5349 22400 8819 22402
rect 5349 22344 5354 22400
rect 5410 22344 8758 22400
rect 8814 22344 8819 22400
rect 5349 22342 8819 22344
rect 5349 22339 5415 22342
rect 8753 22339 8819 22342
rect 3745 22336 4061 22337
rect 3745 22272 3751 22336
rect 3815 22272 3831 22336
rect 3895 22272 3911 22336
rect 3975 22272 3991 22336
rect 4055 22272 4061 22336
rect 3745 22271 4061 22272
rect 9343 22336 9659 22337
rect 9343 22272 9349 22336
rect 9413 22272 9429 22336
rect 9493 22272 9509 22336
rect 9573 22272 9589 22336
rect 9653 22272 9659 22336
rect 9343 22271 9659 22272
rect 14941 22336 15257 22337
rect 14941 22272 14947 22336
rect 15011 22272 15027 22336
rect 15091 22272 15107 22336
rect 15171 22272 15187 22336
rect 15251 22272 15257 22336
rect 14941 22271 15257 22272
rect 20539 22336 20855 22337
rect 20539 22272 20545 22336
rect 20609 22272 20625 22336
rect 20689 22272 20705 22336
rect 20769 22272 20785 22336
rect 20849 22272 20855 22336
rect 20539 22271 20855 22272
rect 4429 22266 4495 22269
rect 7189 22266 7255 22269
rect 4429 22264 7255 22266
rect 4429 22208 4434 22264
rect 4490 22208 7194 22264
rect 7250 22208 7255 22264
rect 4429 22206 7255 22208
rect 4429 22203 4495 22206
rect 7189 22203 7255 22206
rect 10225 22266 10291 22269
rect 13169 22266 13235 22269
rect 10225 22264 13235 22266
rect 10225 22208 10230 22264
rect 10286 22208 13174 22264
rect 13230 22208 13235 22264
rect 10225 22206 13235 22208
rect 10225 22203 10291 22206
rect 13169 22203 13235 22206
rect 2957 22130 3023 22133
rect 3785 22130 3851 22133
rect 20805 22130 20871 22133
rect 2957 22128 20871 22130
rect 2957 22072 2962 22128
rect 3018 22072 3790 22128
rect 3846 22072 20810 22128
rect 20866 22072 20871 22128
rect 2957 22070 20871 22072
rect 2957 22067 3023 22070
rect 3785 22067 3851 22070
rect 20805 22067 20871 22070
rect 22369 22130 22435 22133
rect 23800 22130 24600 22160
rect 22369 22128 24600 22130
rect 22369 22072 22374 22128
rect 22430 22072 24600 22128
rect 22369 22070 24600 22072
rect 22369 22067 22435 22070
rect 23800 22040 24600 22070
rect 3601 21994 3667 21997
rect 3601 21992 5458 21994
rect 3601 21936 3606 21992
rect 3662 21936 5458 21992
rect 3601 21934 5458 21936
rect 3601 21931 3667 21934
rect 2773 21858 2839 21861
rect 4521 21858 4587 21861
rect 2773 21856 4587 21858
rect 2773 21800 2778 21856
rect 2834 21800 4526 21856
rect 4582 21800 4587 21856
rect 2773 21798 4587 21800
rect 5398 21858 5458 21934
rect 5574 21932 5580 21996
rect 5644 21994 5650 21996
rect 6545 21994 6611 21997
rect 5644 21992 6611 21994
rect 5644 21936 6550 21992
rect 6606 21936 6611 21992
rect 5644 21934 6611 21936
rect 5644 21932 5650 21934
rect 6545 21931 6611 21934
rect 6729 21994 6795 21997
rect 9857 21994 9923 21997
rect 6729 21992 9923 21994
rect 6729 21936 6734 21992
rect 6790 21936 9862 21992
rect 9918 21936 9923 21992
rect 6729 21934 9923 21936
rect 6729 21931 6795 21934
rect 9857 21931 9923 21934
rect 10041 21994 10107 21997
rect 21817 21994 21883 21997
rect 10041 21992 21883 21994
rect 10041 21936 10046 21992
rect 10102 21936 21822 21992
rect 21878 21936 21883 21992
rect 10041 21934 21883 21936
rect 10041 21931 10107 21934
rect 21817 21931 21883 21934
rect 6177 21858 6243 21861
rect 5398 21856 6243 21858
rect 5398 21800 6182 21856
rect 6238 21800 6243 21856
rect 5398 21798 6243 21800
rect 2773 21795 2839 21798
rect 4521 21795 4587 21798
rect 6177 21795 6243 21798
rect 7005 21858 7071 21861
rect 8569 21858 8635 21861
rect 7005 21856 8635 21858
rect 7005 21800 7010 21856
rect 7066 21800 8574 21856
rect 8630 21800 8635 21856
rect 7005 21798 8635 21800
rect 7005 21795 7071 21798
rect 8569 21795 8635 21798
rect 8753 21858 8819 21861
rect 9397 21858 9463 21861
rect 13261 21860 13327 21861
rect 13261 21858 13308 21860
rect 8753 21856 9463 21858
rect 8753 21800 8758 21856
rect 8814 21800 9402 21856
rect 9458 21800 9463 21856
rect 8753 21798 9463 21800
rect 13216 21856 13308 21858
rect 13216 21800 13266 21856
rect 13216 21798 13308 21800
rect 8753 21795 8819 21798
rect 9397 21795 9463 21798
rect 13261 21796 13308 21798
rect 13372 21796 13378 21860
rect 15285 21858 15351 21861
rect 15929 21858 15995 21861
rect 18229 21860 18295 21861
rect 18229 21858 18276 21860
rect 15285 21856 15995 21858
rect 15285 21800 15290 21856
rect 15346 21800 15934 21856
rect 15990 21800 15995 21856
rect 15285 21798 15995 21800
rect 18184 21856 18276 21858
rect 18340 21858 18346 21860
rect 22553 21858 22619 21861
rect 18340 21856 22619 21858
rect 18184 21800 18234 21856
rect 18340 21800 22558 21856
rect 22614 21800 22619 21856
rect 18184 21798 18276 21800
rect 13261 21795 13327 21796
rect 15285 21795 15351 21798
rect 15929 21795 15995 21798
rect 18229 21796 18276 21798
rect 18340 21798 22619 21800
rect 18340 21796 18346 21798
rect 18229 21795 18295 21796
rect 22553 21795 22619 21798
rect 6544 21792 6860 21793
rect 6544 21728 6550 21792
rect 6614 21728 6630 21792
rect 6694 21728 6710 21792
rect 6774 21728 6790 21792
rect 6854 21728 6860 21792
rect 6544 21727 6860 21728
rect 12142 21792 12458 21793
rect 12142 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12458 21792
rect 12142 21727 12458 21728
rect 17740 21792 18056 21793
rect 17740 21728 17746 21792
rect 17810 21728 17826 21792
rect 17890 21728 17906 21792
rect 17970 21728 17986 21792
rect 18050 21728 18056 21792
rect 17740 21727 18056 21728
rect 2313 21722 2379 21725
rect 3049 21722 3115 21725
rect 6361 21722 6427 21725
rect 2313 21720 2790 21722
rect 2313 21664 2318 21720
rect 2374 21664 2790 21720
rect 2313 21662 2790 21664
rect 2313 21659 2379 21662
rect 2730 21586 2790 21662
rect 3049 21720 6427 21722
rect 3049 21664 3054 21720
rect 3110 21664 6366 21720
rect 6422 21664 6427 21720
rect 3049 21662 6427 21664
rect 3049 21659 3115 21662
rect 6361 21659 6427 21662
rect 7097 21722 7163 21725
rect 15326 21722 15332 21724
rect 7097 21720 12082 21722
rect 7097 21664 7102 21720
rect 7158 21664 12082 21720
rect 7097 21662 12082 21664
rect 7097 21659 7163 21662
rect 10041 21586 10107 21589
rect 2730 21584 10107 21586
rect 2730 21528 10046 21584
rect 10102 21528 10107 21584
rect 2730 21526 10107 21528
rect 12022 21586 12082 21662
rect 13126 21662 15332 21722
rect 13126 21586 13186 21662
rect 15326 21660 15332 21662
rect 15396 21722 15402 21724
rect 15837 21722 15903 21725
rect 15396 21720 15903 21722
rect 15396 21664 15842 21720
rect 15898 21664 15903 21720
rect 15396 21662 15903 21664
rect 15396 21660 15402 21662
rect 15837 21659 15903 21662
rect 18137 21722 18203 21725
rect 19241 21722 19307 21725
rect 18137 21720 19307 21722
rect 18137 21664 18142 21720
rect 18198 21664 19246 21720
rect 19302 21664 19307 21720
rect 18137 21662 19307 21664
rect 18137 21659 18203 21662
rect 19241 21659 19307 21662
rect 12022 21526 13186 21586
rect 13261 21586 13327 21589
rect 16297 21586 16363 21589
rect 13261 21584 16363 21586
rect 13261 21528 13266 21584
rect 13322 21528 16302 21584
rect 16358 21528 16363 21584
rect 13261 21526 16363 21528
rect 10041 21523 10107 21526
rect 13261 21523 13327 21526
rect 16297 21523 16363 21526
rect 17125 21586 17191 21589
rect 19425 21586 19491 21589
rect 17125 21584 19491 21586
rect 17125 21528 17130 21584
rect 17186 21528 19430 21584
rect 19486 21528 19491 21584
rect 17125 21526 19491 21528
rect 17125 21523 17191 21526
rect 19425 21523 19491 21526
rect 20069 21586 20135 21589
rect 22461 21586 22527 21589
rect 20069 21584 22527 21586
rect 20069 21528 20074 21584
rect 20130 21528 22466 21584
rect 22522 21528 22527 21584
rect 20069 21526 22527 21528
rect 20069 21523 20135 21526
rect 22461 21523 22527 21526
rect 22645 21586 22711 21589
rect 23800 21586 24600 21616
rect 22645 21584 24600 21586
rect 22645 21528 22650 21584
rect 22706 21528 24600 21584
rect 22645 21526 24600 21528
rect 22645 21523 22711 21526
rect 23800 21496 24600 21526
rect 0 21360 800 21480
rect 3417 21450 3483 21453
rect 9121 21450 9187 21453
rect 11421 21450 11487 21453
rect 21357 21450 21423 21453
rect 3417 21448 11487 21450
rect 3417 21392 3422 21448
rect 3478 21392 9126 21448
rect 9182 21392 11426 21448
rect 11482 21392 11487 21448
rect 3417 21390 11487 21392
rect 3417 21387 3483 21390
rect 9121 21387 9187 21390
rect 11421 21387 11487 21390
rect 12390 21448 21423 21450
rect 12390 21392 21362 21448
rect 21418 21392 21423 21448
rect 12390 21390 21423 21392
rect 4521 21314 4587 21317
rect 7097 21314 7163 21317
rect 4521 21312 7163 21314
rect 4521 21256 4526 21312
rect 4582 21256 7102 21312
rect 7158 21256 7163 21312
rect 4521 21254 7163 21256
rect 4521 21251 4587 21254
rect 7097 21251 7163 21254
rect 9765 21314 9831 21317
rect 12390 21314 12450 21390
rect 21357 21387 21423 21390
rect 19241 21314 19307 21317
rect 9765 21312 12450 21314
rect 9765 21256 9770 21312
rect 9826 21256 12450 21312
rect 9765 21254 12450 21256
rect 15334 21312 19307 21314
rect 15334 21256 19246 21312
rect 19302 21256 19307 21312
rect 15334 21254 19307 21256
rect 9765 21251 9831 21254
rect 3745 21248 4061 21249
rect 3745 21184 3751 21248
rect 3815 21184 3831 21248
rect 3895 21184 3911 21248
rect 3975 21184 3991 21248
rect 4055 21184 4061 21248
rect 3745 21183 4061 21184
rect 9343 21248 9659 21249
rect 9343 21184 9349 21248
rect 9413 21184 9429 21248
rect 9493 21184 9509 21248
rect 9573 21184 9589 21248
rect 9653 21184 9659 21248
rect 9343 21183 9659 21184
rect 14941 21248 15257 21249
rect 14941 21184 14947 21248
rect 15011 21184 15027 21248
rect 15091 21184 15107 21248
rect 15171 21184 15187 21248
rect 15251 21184 15257 21248
rect 14941 21183 15257 21184
rect 6085 21178 6151 21181
rect 8753 21178 8819 21181
rect 9121 21178 9187 21181
rect 6085 21176 9187 21178
rect 6085 21120 6090 21176
rect 6146 21120 8758 21176
rect 8814 21120 9126 21176
rect 9182 21120 9187 21176
rect 6085 21118 9187 21120
rect 6085 21115 6151 21118
rect 8753 21115 8819 21118
rect 9121 21115 9187 21118
rect 3417 21042 3483 21045
rect 12566 21042 12572 21044
rect 3417 21040 12572 21042
rect 3417 20984 3422 21040
rect 3478 20984 12572 21040
rect 3417 20982 12572 20984
rect 3417 20979 3483 20982
rect 12566 20980 12572 20982
rect 12636 21042 12642 21044
rect 13721 21042 13787 21045
rect 15334 21042 15394 21254
rect 19241 21251 19307 21254
rect 20539 21248 20855 21249
rect 20539 21184 20545 21248
rect 20609 21184 20625 21248
rect 20689 21184 20705 21248
rect 20769 21184 20785 21248
rect 20849 21184 20855 21248
rect 20539 21183 20855 21184
rect 15929 21178 15995 21181
rect 20069 21178 20135 21181
rect 15929 21176 20135 21178
rect 15929 21120 15934 21176
rect 15990 21120 20074 21176
rect 20130 21120 20135 21176
rect 15929 21118 20135 21120
rect 15929 21115 15995 21118
rect 20069 21115 20135 21118
rect 21081 21042 21147 21045
rect 12636 21040 15394 21042
rect 12636 20984 13726 21040
rect 13782 20984 15394 21040
rect 12636 20982 15394 20984
rect 16070 21040 21147 21042
rect 16070 20984 21086 21040
rect 21142 20984 21147 21040
rect 16070 20982 21147 20984
rect 12636 20980 12642 20982
rect 13721 20979 13787 20982
rect 2037 20906 2103 20909
rect 2681 20906 2747 20909
rect 4245 20906 4311 20909
rect 4838 20906 4844 20908
rect 2037 20904 2790 20906
rect 2037 20848 2042 20904
rect 2098 20848 2686 20904
rect 2742 20848 2790 20904
rect 2037 20846 2790 20848
rect 2037 20843 2103 20846
rect 2681 20843 2790 20846
rect 4245 20904 4844 20906
rect 4245 20848 4250 20904
rect 4306 20848 4844 20904
rect 4245 20846 4844 20848
rect 4245 20843 4311 20846
rect 4838 20844 4844 20846
rect 4908 20844 4914 20908
rect 6310 20844 6316 20908
rect 6380 20906 6386 20908
rect 6637 20906 6703 20909
rect 6380 20904 6703 20906
rect 6380 20848 6642 20904
rect 6698 20848 6703 20904
rect 6380 20846 6703 20848
rect 6380 20844 6386 20846
rect 6637 20843 6703 20846
rect 6821 20906 6887 20909
rect 10133 20906 10199 20909
rect 6821 20904 10199 20906
rect 6821 20848 6826 20904
rect 6882 20848 10138 20904
rect 10194 20848 10199 20904
rect 6821 20846 10199 20848
rect 6821 20843 6887 20846
rect 10133 20843 10199 20846
rect 15377 20906 15443 20909
rect 16070 20906 16130 20982
rect 21081 20979 21147 20982
rect 23013 21042 23079 21045
rect 23800 21042 24600 21072
rect 23013 21040 24600 21042
rect 23013 20984 23018 21040
rect 23074 20984 24600 21040
rect 23013 20982 24600 20984
rect 23013 20979 23079 20982
rect 23800 20952 24600 20982
rect 15377 20904 16130 20906
rect 15377 20848 15382 20904
rect 15438 20848 16130 20904
rect 15377 20846 16130 20848
rect 16665 20906 16731 20909
rect 18413 20906 18479 20909
rect 16665 20904 18479 20906
rect 16665 20848 16670 20904
rect 16726 20848 18418 20904
rect 18474 20848 18479 20904
rect 16665 20846 18479 20848
rect 15377 20843 15443 20846
rect 16665 20843 16731 20846
rect 18413 20843 18479 20846
rect 19241 20906 19307 20909
rect 22093 20906 22159 20909
rect 19241 20904 22159 20906
rect 19241 20848 19246 20904
rect 19302 20848 22098 20904
rect 22154 20848 22159 20904
rect 19241 20846 22159 20848
rect 19241 20843 19307 20846
rect 22093 20843 22159 20846
rect 2730 20770 2790 20843
rect 6085 20770 6151 20773
rect 14457 20770 14523 20773
rect 17033 20770 17099 20773
rect 2730 20768 6151 20770
rect 2730 20712 6090 20768
rect 6146 20712 6151 20768
rect 2730 20710 6151 20712
rect 6085 20707 6151 20710
rect 12758 20768 14523 20770
rect 12758 20712 14462 20768
rect 14518 20712 14523 20768
rect 12758 20710 14523 20712
rect 6544 20704 6860 20705
rect 6544 20640 6550 20704
rect 6614 20640 6630 20704
rect 6694 20640 6710 20704
rect 6774 20640 6790 20704
rect 6854 20640 6860 20704
rect 6544 20639 6860 20640
rect 12142 20704 12458 20705
rect 12142 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12458 20704
rect 12142 20639 12458 20640
rect 3141 20634 3207 20637
rect 4797 20634 4863 20637
rect 3141 20632 4863 20634
rect 3141 20576 3146 20632
rect 3202 20576 4802 20632
rect 4858 20576 4863 20632
rect 3141 20574 4863 20576
rect 3141 20571 3207 20574
rect 4797 20571 4863 20574
rect 4981 20634 5047 20637
rect 6269 20634 6335 20637
rect 4981 20632 6335 20634
rect 4981 20576 4986 20632
rect 5042 20576 6274 20632
rect 6330 20576 6335 20632
rect 4981 20574 6335 20576
rect 4981 20571 5047 20574
rect 6269 20571 6335 20574
rect 3233 20498 3299 20501
rect 12758 20498 12818 20710
rect 14457 20707 14523 20710
rect 15150 20768 17099 20770
rect 15150 20712 17038 20768
rect 17094 20712 17099 20768
rect 15150 20710 17099 20712
rect 13629 20634 13695 20637
rect 15150 20634 15210 20710
rect 17033 20707 17099 20710
rect 17740 20704 18056 20705
rect 17740 20640 17746 20704
rect 17810 20640 17826 20704
rect 17890 20640 17906 20704
rect 17970 20640 17986 20704
rect 18050 20640 18056 20704
rect 17740 20639 18056 20640
rect 13629 20632 15210 20634
rect 13629 20576 13634 20632
rect 13690 20576 15210 20632
rect 13629 20574 15210 20576
rect 18321 20634 18387 20637
rect 19057 20634 19123 20637
rect 18321 20632 19123 20634
rect 18321 20576 18326 20632
rect 18382 20576 19062 20632
rect 19118 20576 19123 20632
rect 18321 20574 19123 20576
rect 13629 20571 13695 20574
rect 18321 20571 18387 20574
rect 19057 20571 19123 20574
rect 19609 20634 19675 20637
rect 21541 20634 21607 20637
rect 19609 20632 21607 20634
rect 19609 20576 19614 20632
rect 19670 20576 21546 20632
rect 21602 20576 21607 20632
rect 19609 20574 21607 20576
rect 19609 20571 19675 20574
rect 21541 20571 21607 20574
rect 16941 20500 17007 20501
rect 16941 20498 16988 20500
rect 3233 20496 12818 20498
rect 3233 20440 3238 20496
rect 3294 20440 12818 20496
rect 3233 20438 12818 20440
rect 16860 20496 16988 20498
rect 17052 20498 17058 20500
rect 17677 20498 17743 20501
rect 17052 20496 17743 20498
rect 16860 20440 16946 20496
rect 17052 20440 17682 20496
rect 17738 20440 17743 20496
rect 16860 20438 16988 20440
rect 3233 20435 3299 20438
rect 16941 20436 16988 20438
rect 17052 20438 17743 20440
rect 17052 20436 17058 20438
rect 16941 20435 17007 20436
rect 17677 20435 17743 20438
rect 17861 20498 17927 20501
rect 21357 20498 21423 20501
rect 17861 20496 21423 20498
rect 17861 20440 17866 20496
rect 17922 20440 21362 20496
rect 21418 20440 21423 20496
rect 17861 20438 21423 20440
rect 17861 20435 17927 20438
rect 21357 20435 21423 20438
rect 23013 20498 23079 20501
rect 23800 20498 24600 20528
rect 23013 20496 24600 20498
rect 23013 20440 23018 20496
rect 23074 20440 24600 20496
rect 23013 20438 24600 20440
rect 23013 20435 23079 20438
rect 23800 20408 24600 20438
rect 7281 20362 7347 20365
rect 18321 20362 18387 20365
rect 7281 20360 18387 20362
rect 7281 20304 7286 20360
rect 7342 20304 18326 20360
rect 18382 20304 18387 20360
rect 7281 20302 18387 20304
rect 7281 20299 7347 20302
rect 18321 20299 18387 20302
rect 16481 20226 16547 20229
rect 17953 20226 18019 20229
rect 18873 20226 18939 20229
rect 16481 20224 18939 20226
rect 16481 20168 16486 20224
rect 16542 20168 17958 20224
rect 18014 20168 18878 20224
rect 18934 20168 18939 20224
rect 16481 20166 18939 20168
rect 16481 20163 16547 20166
rect 17953 20163 18019 20166
rect 18873 20163 18939 20166
rect 3745 20160 4061 20161
rect 3745 20096 3751 20160
rect 3815 20096 3831 20160
rect 3895 20096 3911 20160
rect 3975 20096 3991 20160
rect 4055 20096 4061 20160
rect 3745 20095 4061 20096
rect 9343 20160 9659 20161
rect 9343 20096 9349 20160
rect 9413 20096 9429 20160
rect 9493 20096 9509 20160
rect 9573 20096 9589 20160
rect 9653 20096 9659 20160
rect 9343 20095 9659 20096
rect 14941 20160 15257 20161
rect 14941 20096 14947 20160
rect 15011 20096 15027 20160
rect 15091 20096 15107 20160
rect 15171 20096 15187 20160
rect 15251 20096 15257 20160
rect 14941 20095 15257 20096
rect 20539 20160 20855 20161
rect 20539 20096 20545 20160
rect 20609 20096 20625 20160
rect 20689 20096 20705 20160
rect 20769 20096 20785 20160
rect 20849 20096 20855 20160
rect 20539 20095 20855 20096
rect 15653 20090 15719 20093
rect 16430 20090 16436 20092
rect 15653 20088 16436 20090
rect 15653 20032 15658 20088
rect 15714 20032 16436 20088
rect 15653 20030 16436 20032
rect 15653 20027 15719 20030
rect 16430 20028 16436 20030
rect 16500 20028 16506 20092
rect 5717 19954 5783 19957
rect 12709 19954 12775 19957
rect 5717 19952 12775 19954
rect 5717 19896 5722 19952
rect 5778 19896 12714 19952
rect 12770 19896 12775 19952
rect 5717 19894 12775 19896
rect 5717 19891 5783 19894
rect 12709 19891 12775 19894
rect 13261 19954 13327 19957
rect 22829 19954 22895 19957
rect 13261 19952 22895 19954
rect 13261 19896 13266 19952
rect 13322 19896 22834 19952
rect 22890 19896 22895 19952
rect 13261 19894 22895 19896
rect 13261 19891 13327 19894
rect 22829 19891 22895 19894
rect 23105 19954 23171 19957
rect 23800 19954 24600 19984
rect 23105 19952 24600 19954
rect 23105 19896 23110 19952
rect 23166 19896 24600 19952
rect 23105 19894 24600 19896
rect 23105 19891 23171 19894
rect 23800 19864 24600 19894
rect 17953 19818 18019 19821
rect 19241 19818 19307 19821
rect 20713 19818 20779 19821
rect 17953 19816 20779 19818
rect 17953 19760 17958 19816
rect 18014 19760 19246 19816
rect 19302 19760 20718 19816
rect 20774 19760 20779 19816
rect 17953 19758 20779 19760
rect 17953 19755 18019 19758
rect 19241 19755 19307 19758
rect 20713 19755 20779 19758
rect 19425 19682 19491 19685
rect 21081 19682 21147 19685
rect 19425 19680 21147 19682
rect 19425 19624 19430 19680
rect 19486 19624 21086 19680
rect 21142 19624 21147 19680
rect 19425 19622 21147 19624
rect 19425 19619 19491 19622
rect 21081 19619 21147 19622
rect 6544 19616 6860 19617
rect 6544 19552 6550 19616
rect 6614 19552 6630 19616
rect 6694 19552 6710 19616
rect 6774 19552 6790 19616
rect 6854 19552 6860 19616
rect 6544 19551 6860 19552
rect 12142 19616 12458 19617
rect 12142 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12458 19616
rect 12142 19551 12458 19552
rect 17740 19616 18056 19617
rect 17740 19552 17746 19616
rect 17810 19552 17826 19616
rect 17890 19552 17906 19616
rect 17970 19552 17986 19616
rect 18050 19552 18056 19616
rect 17740 19551 18056 19552
rect 12893 19546 12959 19549
rect 16113 19546 16179 19549
rect 16481 19548 16547 19549
rect 12528 19544 16179 19546
rect 12528 19488 12898 19544
rect 12954 19488 16118 19544
rect 16174 19488 16179 19544
rect 12528 19486 16179 19488
rect 11329 19410 11395 19413
rect 12528 19410 12588 19486
rect 12893 19483 12959 19486
rect 16113 19483 16179 19486
rect 16430 19484 16436 19548
rect 16500 19546 16547 19548
rect 18321 19546 18387 19549
rect 18454 19546 18460 19548
rect 16500 19544 16592 19546
rect 16542 19488 16592 19544
rect 16500 19486 16592 19488
rect 18321 19544 18460 19546
rect 18321 19488 18326 19544
rect 18382 19488 18460 19544
rect 18321 19486 18460 19488
rect 16500 19484 16547 19486
rect 16481 19483 16547 19484
rect 18321 19483 18387 19486
rect 18454 19484 18460 19486
rect 18524 19484 18530 19548
rect 19425 19546 19491 19549
rect 20989 19546 21055 19549
rect 19425 19544 21055 19546
rect 19425 19488 19430 19544
rect 19486 19488 20994 19544
rect 21050 19488 21055 19544
rect 19425 19486 21055 19488
rect 19425 19483 19491 19486
rect 20989 19483 21055 19486
rect 11329 19408 12588 19410
rect 11329 19352 11334 19408
rect 11390 19352 12588 19408
rect 11329 19350 12588 19352
rect 14549 19410 14615 19413
rect 16389 19410 16455 19413
rect 16573 19412 16639 19413
rect 14549 19408 16498 19410
rect 14549 19352 14554 19408
rect 14610 19352 16394 19408
rect 16450 19352 16498 19408
rect 14549 19350 16498 19352
rect 11329 19347 11395 19350
rect 14549 19347 14615 19350
rect 16389 19347 16498 19350
rect 16573 19408 16620 19412
rect 16684 19410 16690 19412
rect 16573 19352 16578 19408
rect 16573 19348 16620 19352
rect 16684 19350 16730 19410
rect 16684 19348 16690 19350
rect 16982 19348 16988 19412
rect 17052 19348 17058 19412
rect 17217 19410 17283 19413
rect 21265 19410 21331 19413
rect 17217 19408 21331 19410
rect 17217 19352 17222 19408
rect 17278 19352 21270 19408
rect 21326 19352 21331 19408
rect 17217 19350 21331 19352
rect 16573 19347 16639 19348
rect 16438 19138 16498 19347
rect 16573 19274 16639 19277
rect 16990 19274 17050 19348
rect 17217 19347 17283 19350
rect 21265 19347 21331 19350
rect 23289 19410 23355 19413
rect 23800 19410 24600 19440
rect 23289 19408 24600 19410
rect 23289 19352 23294 19408
rect 23350 19352 24600 19408
rect 23289 19350 24600 19352
rect 23289 19347 23355 19350
rect 23800 19320 24600 19350
rect 23105 19274 23171 19277
rect 16573 19272 17050 19274
rect 16573 19216 16578 19272
rect 16634 19216 17050 19272
rect 16573 19214 17050 19216
rect 17542 19272 23171 19274
rect 17542 19216 23110 19272
rect 23166 19216 23171 19272
rect 17542 19214 23171 19216
rect 16573 19211 16639 19214
rect 17542 19138 17602 19214
rect 23105 19211 23171 19214
rect 16438 19078 17602 19138
rect 3745 19072 4061 19073
rect 3745 19008 3751 19072
rect 3815 19008 3831 19072
rect 3895 19008 3911 19072
rect 3975 19008 3991 19072
rect 4055 19008 4061 19072
rect 3745 19007 4061 19008
rect 9343 19072 9659 19073
rect 9343 19008 9349 19072
rect 9413 19008 9429 19072
rect 9493 19008 9509 19072
rect 9573 19008 9589 19072
rect 9653 19008 9659 19072
rect 9343 19007 9659 19008
rect 14941 19072 15257 19073
rect 14941 19008 14947 19072
rect 15011 19008 15027 19072
rect 15091 19008 15107 19072
rect 15171 19008 15187 19072
rect 15251 19008 15257 19072
rect 14941 19007 15257 19008
rect 20539 19072 20855 19073
rect 20539 19008 20545 19072
rect 20609 19008 20625 19072
rect 20689 19008 20705 19072
rect 20769 19008 20785 19072
rect 20849 19008 20855 19072
rect 20539 19007 20855 19008
rect 5441 18866 5507 18869
rect 5625 18866 5691 18869
rect 5441 18864 5691 18866
rect 5441 18808 5446 18864
rect 5502 18808 5630 18864
rect 5686 18808 5691 18864
rect 5441 18806 5691 18808
rect 5441 18803 5507 18806
rect 5625 18803 5691 18806
rect 13302 18804 13308 18868
rect 13372 18866 13378 18868
rect 19926 18866 19932 18868
rect 13372 18806 19932 18866
rect 13372 18804 13378 18806
rect 19926 18804 19932 18806
rect 19996 18804 20002 18868
rect 23013 18866 23079 18869
rect 23800 18866 24600 18896
rect 23013 18864 24600 18866
rect 23013 18808 23018 18864
rect 23074 18808 24600 18864
rect 23013 18806 24600 18808
rect 23013 18803 23079 18806
rect 23800 18776 24600 18806
rect 3509 18730 3575 18733
rect 6085 18730 6151 18733
rect 3509 18728 6151 18730
rect 3509 18672 3514 18728
rect 3570 18672 6090 18728
rect 6146 18672 6151 18728
rect 3509 18670 6151 18672
rect 3509 18667 3575 18670
rect 6085 18667 6151 18670
rect 14457 18730 14523 18733
rect 22277 18730 22343 18733
rect 14457 18728 22343 18730
rect 14457 18672 14462 18728
rect 14518 18672 22282 18728
rect 22338 18672 22343 18728
rect 14457 18670 22343 18672
rect 14457 18667 14523 18670
rect 22277 18667 22343 18670
rect 3877 18594 3943 18597
rect 5165 18594 5231 18597
rect 3877 18592 5231 18594
rect 3877 18536 3882 18592
rect 3938 18536 5170 18592
rect 5226 18536 5231 18592
rect 3877 18534 5231 18536
rect 3877 18531 3943 18534
rect 5165 18531 5231 18534
rect 19701 18594 19767 18597
rect 23197 18594 23263 18597
rect 19701 18592 23263 18594
rect 19701 18536 19706 18592
rect 19762 18536 23202 18592
rect 23258 18536 23263 18592
rect 19701 18534 23263 18536
rect 19701 18531 19767 18534
rect 23197 18531 23263 18534
rect 6544 18528 6860 18529
rect 6544 18464 6550 18528
rect 6614 18464 6630 18528
rect 6694 18464 6710 18528
rect 6774 18464 6790 18528
rect 6854 18464 6860 18528
rect 6544 18463 6860 18464
rect 12142 18528 12458 18529
rect 12142 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12458 18528
rect 12142 18463 12458 18464
rect 17740 18528 18056 18529
rect 17740 18464 17746 18528
rect 17810 18464 17826 18528
rect 17890 18464 17906 18528
rect 17970 18464 17986 18528
rect 18050 18464 18056 18528
rect 17740 18463 18056 18464
rect 3417 18458 3483 18461
rect 5257 18458 5323 18461
rect 3417 18456 5323 18458
rect 3417 18400 3422 18456
rect 3478 18400 5262 18456
rect 5318 18400 5323 18456
rect 3417 18398 5323 18400
rect 3417 18395 3483 18398
rect 5257 18395 5323 18398
rect 13077 18458 13143 18461
rect 14273 18458 14339 18461
rect 14917 18458 14983 18461
rect 13077 18456 14983 18458
rect 13077 18400 13082 18456
rect 13138 18400 14278 18456
rect 14334 18400 14922 18456
rect 14978 18400 14983 18456
rect 13077 18398 14983 18400
rect 13077 18395 13143 18398
rect 14273 18395 14339 18398
rect 14917 18395 14983 18398
rect 2773 18322 2839 18325
rect 7189 18322 7255 18325
rect 2773 18320 7255 18322
rect 2773 18264 2778 18320
rect 2834 18264 7194 18320
rect 7250 18264 7255 18320
rect 2773 18262 7255 18264
rect 2773 18259 2839 18262
rect 7189 18259 7255 18262
rect 12985 18322 13051 18325
rect 14273 18322 14339 18325
rect 12985 18320 14339 18322
rect 12985 18264 12990 18320
rect 13046 18264 14278 18320
rect 14334 18264 14339 18320
rect 12985 18262 14339 18264
rect 12985 18259 13051 18262
rect 14273 18259 14339 18262
rect 15285 18322 15351 18325
rect 22369 18322 22435 18325
rect 15285 18320 22435 18322
rect 15285 18264 15290 18320
rect 15346 18264 22374 18320
rect 22430 18264 22435 18320
rect 15285 18262 22435 18264
rect 15285 18259 15351 18262
rect 22369 18259 22435 18262
rect 23105 18322 23171 18325
rect 23800 18322 24600 18352
rect 23105 18320 24600 18322
rect 23105 18264 23110 18320
rect 23166 18264 24600 18320
rect 23105 18262 24600 18264
rect 23105 18259 23171 18262
rect 23800 18232 24600 18262
rect 4981 18186 5047 18189
rect 8661 18186 8727 18189
rect 4981 18184 8727 18186
rect 4981 18128 4986 18184
rect 5042 18128 8666 18184
rect 8722 18128 8727 18184
rect 4981 18126 8727 18128
rect 4981 18123 5047 18126
rect 8661 18123 8727 18126
rect 16941 18186 17007 18189
rect 20805 18186 20871 18189
rect 16941 18184 20871 18186
rect 16941 18128 16946 18184
rect 17002 18128 20810 18184
rect 20866 18128 20871 18184
rect 16941 18126 20871 18128
rect 16941 18123 17007 18126
rect 20805 18123 20871 18126
rect 4153 18050 4219 18053
rect 5165 18050 5231 18053
rect 6453 18050 6519 18053
rect 4153 18048 6519 18050
rect 4153 17992 4158 18048
rect 4214 17992 5170 18048
rect 5226 17992 6458 18048
rect 6514 17992 6519 18048
rect 4153 17990 6519 17992
rect 4153 17987 4219 17990
rect 5165 17987 5231 17990
rect 6453 17987 6519 17990
rect 3745 17984 4061 17985
rect 3745 17920 3751 17984
rect 3815 17920 3831 17984
rect 3895 17920 3911 17984
rect 3975 17920 3991 17984
rect 4055 17920 4061 17984
rect 3745 17919 4061 17920
rect 9343 17984 9659 17985
rect 9343 17920 9349 17984
rect 9413 17920 9429 17984
rect 9493 17920 9509 17984
rect 9573 17920 9589 17984
rect 9653 17920 9659 17984
rect 9343 17919 9659 17920
rect 14941 17984 15257 17985
rect 14941 17920 14947 17984
rect 15011 17920 15027 17984
rect 15091 17920 15107 17984
rect 15171 17920 15187 17984
rect 15251 17920 15257 17984
rect 14941 17919 15257 17920
rect 20539 17984 20855 17985
rect 20539 17920 20545 17984
rect 20609 17920 20625 17984
rect 20689 17920 20705 17984
rect 20769 17920 20785 17984
rect 20849 17920 20855 17984
rect 20539 17919 20855 17920
rect 6913 17778 6979 17781
rect 11421 17778 11487 17781
rect 6913 17776 11487 17778
rect 6913 17720 6918 17776
rect 6974 17720 11426 17776
rect 11482 17720 11487 17776
rect 6913 17718 11487 17720
rect 6913 17715 6979 17718
rect 11421 17715 11487 17718
rect 13721 17778 13787 17781
rect 21817 17778 21883 17781
rect 23800 17778 24600 17808
rect 13721 17776 21883 17778
rect 13721 17720 13726 17776
rect 13782 17720 21822 17776
rect 21878 17720 21883 17776
rect 13721 17718 21883 17720
rect 13721 17715 13787 17718
rect 21817 17715 21883 17718
rect 22050 17718 24600 17778
rect 4061 17642 4127 17645
rect 7465 17642 7531 17645
rect 4061 17640 7531 17642
rect 4061 17584 4066 17640
rect 4122 17584 7470 17640
rect 7526 17584 7531 17640
rect 4061 17582 7531 17584
rect 4061 17579 4127 17582
rect 7465 17579 7531 17582
rect 11329 17642 11395 17645
rect 15326 17642 15332 17644
rect 11329 17640 15332 17642
rect 11329 17584 11334 17640
rect 11390 17584 15332 17640
rect 11329 17582 15332 17584
rect 11329 17579 11395 17582
rect 15326 17580 15332 17582
rect 15396 17580 15402 17644
rect 18781 17642 18847 17645
rect 17588 17640 18847 17642
rect 17588 17584 18786 17640
rect 18842 17584 18847 17640
rect 17588 17582 18847 17584
rect 17401 17506 17467 17509
rect 17588 17506 17648 17582
rect 18781 17579 18847 17582
rect 17401 17504 17648 17506
rect 17401 17448 17406 17504
rect 17462 17448 17648 17504
rect 17401 17446 17648 17448
rect 21817 17506 21883 17509
rect 22050 17506 22110 17718
rect 23800 17688 24600 17718
rect 22185 17642 22251 17645
rect 22737 17642 22803 17645
rect 22185 17640 22803 17642
rect 22185 17584 22190 17640
rect 22246 17584 22742 17640
rect 22798 17584 22803 17640
rect 22185 17582 22803 17584
rect 22185 17579 22251 17582
rect 22737 17579 22803 17582
rect 21817 17504 22110 17506
rect 21817 17448 21822 17504
rect 21878 17448 22110 17504
rect 21817 17446 22110 17448
rect 17401 17443 17467 17446
rect 21817 17443 21883 17446
rect 6544 17440 6860 17441
rect 6544 17376 6550 17440
rect 6614 17376 6630 17440
rect 6694 17376 6710 17440
rect 6774 17376 6790 17440
rect 6854 17376 6860 17440
rect 6544 17375 6860 17376
rect 12142 17440 12458 17441
rect 12142 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12458 17440
rect 12142 17375 12458 17376
rect 17740 17440 18056 17441
rect 17740 17376 17746 17440
rect 17810 17376 17826 17440
rect 17890 17376 17906 17440
rect 17970 17376 17986 17440
rect 18050 17376 18056 17440
rect 17740 17375 18056 17376
rect 16205 17234 16271 17237
rect 22645 17234 22711 17237
rect 16205 17232 22711 17234
rect 16205 17176 16210 17232
rect 16266 17176 22650 17232
rect 22706 17176 22711 17232
rect 16205 17174 22711 17176
rect 16205 17171 16271 17174
rect 22645 17171 22711 17174
rect 23105 17234 23171 17237
rect 23800 17234 24600 17264
rect 23105 17232 24600 17234
rect 23105 17176 23110 17232
rect 23166 17176 24600 17232
rect 23105 17174 24600 17176
rect 23105 17171 23171 17174
rect 23800 17144 24600 17174
rect 14457 17098 14523 17101
rect 22737 17098 22803 17101
rect 14457 17096 22803 17098
rect 14457 17040 14462 17096
rect 14518 17040 22742 17096
rect 22798 17040 22803 17096
rect 14457 17038 22803 17040
rect 14457 17035 14523 17038
rect 22737 17035 22803 17038
rect 3745 16896 4061 16897
rect 3745 16832 3751 16896
rect 3815 16832 3831 16896
rect 3895 16832 3911 16896
rect 3975 16832 3991 16896
rect 4055 16832 4061 16896
rect 3745 16831 4061 16832
rect 9343 16896 9659 16897
rect 9343 16832 9349 16896
rect 9413 16832 9429 16896
rect 9493 16832 9509 16896
rect 9573 16832 9589 16896
rect 9653 16832 9659 16896
rect 9343 16831 9659 16832
rect 14941 16896 15257 16897
rect 14941 16832 14947 16896
rect 15011 16832 15027 16896
rect 15091 16832 15107 16896
rect 15171 16832 15187 16896
rect 15251 16832 15257 16896
rect 14941 16831 15257 16832
rect 20539 16896 20855 16897
rect 20539 16832 20545 16896
rect 20609 16832 20625 16896
rect 20689 16832 20705 16896
rect 20769 16832 20785 16896
rect 20849 16832 20855 16896
rect 20539 16831 20855 16832
rect 19333 16690 19399 16693
rect 23800 16690 24600 16720
rect 19333 16688 24600 16690
rect 19333 16632 19338 16688
rect 19394 16632 24600 16688
rect 19333 16630 24600 16632
rect 19333 16627 19399 16630
rect 23800 16600 24600 16630
rect 11145 16554 11211 16557
rect 12566 16554 12572 16556
rect 11145 16552 12572 16554
rect 11145 16496 11150 16552
rect 11206 16496 12572 16552
rect 11145 16494 12572 16496
rect 11145 16491 11211 16494
rect 12566 16492 12572 16494
rect 12636 16492 12642 16556
rect 21081 16554 21147 16557
rect 21541 16554 21607 16557
rect 21081 16552 21607 16554
rect 21081 16496 21086 16552
rect 21142 16496 21546 16552
rect 21602 16496 21607 16552
rect 21081 16494 21607 16496
rect 21081 16491 21147 16494
rect 21541 16491 21607 16494
rect 20621 16418 20687 16421
rect 22369 16418 22435 16421
rect 20621 16416 22435 16418
rect 20621 16360 20626 16416
rect 20682 16360 22374 16416
rect 22430 16360 22435 16416
rect 20621 16358 22435 16360
rect 20621 16355 20687 16358
rect 22369 16355 22435 16358
rect 6544 16352 6860 16353
rect 6544 16288 6550 16352
rect 6614 16288 6630 16352
rect 6694 16288 6710 16352
rect 6774 16288 6790 16352
rect 6854 16288 6860 16352
rect 6544 16287 6860 16288
rect 12142 16352 12458 16353
rect 12142 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12458 16352
rect 12142 16287 12458 16288
rect 17740 16352 18056 16353
rect 17740 16288 17746 16352
rect 17810 16288 17826 16352
rect 17890 16288 17906 16352
rect 17970 16288 17986 16352
rect 18050 16288 18056 16352
rect 17740 16287 18056 16288
rect 18689 16282 18755 16285
rect 21173 16282 21239 16285
rect 18689 16280 21239 16282
rect 18689 16224 18694 16280
rect 18750 16224 21178 16280
rect 21234 16224 21239 16280
rect 18689 16222 21239 16224
rect 18689 16219 18755 16222
rect 21173 16219 21239 16222
rect 21357 16282 21423 16285
rect 22369 16282 22435 16285
rect 21357 16280 22435 16282
rect 21357 16224 21362 16280
rect 21418 16224 22374 16280
rect 22430 16224 22435 16280
rect 21357 16222 22435 16224
rect 21357 16219 21423 16222
rect 22369 16219 22435 16222
rect 10685 16146 10751 16149
rect 21081 16146 21147 16149
rect 10685 16144 21147 16146
rect 10685 16088 10690 16144
rect 10746 16088 21086 16144
rect 21142 16088 21147 16144
rect 10685 16086 21147 16088
rect 10685 16083 10751 16086
rect 21081 16083 21147 16086
rect 21265 16146 21331 16149
rect 23800 16146 24600 16176
rect 21265 16144 24600 16146
rect 21265 16088 21270 16144
rect 21326 16088 24600 16144
rect 21265 16086 24600 16088
rect 21265 16083 21331 16086
rect 23800 16056 24600 16086
rect 16481 16010 16547 16013
rect 23657 16010 23723 16013
rect 16481 16008 23723 16010
rect 16481 15952 16486 16008
rect 16542 15952 23662 16008
rect 23718 15952 23723 16008
rect 16481 15950 23723 15952
rect 16481 15947 16547 15950
rect 23657 15947 23723 15950
rect 3745 15808 4061 15809
rect 3745 15744 3751 15808
rect 3815 15744 3831 15808
rect 3895 15744 3911 15808
rect 3975 15744 3991 15808
rect 4055 15744 4061 15808
rect 3745 15743 4061 15744
rect 9343 15808 9659 15809
rect 9343 15744 9349 15808
rect 9413 15744 9429 15808
rect 9493 15744 9509 15808
rect 9573 15744 9589 15808
rect 9653 15744 9659 15808
rect 9343 15743 9659 15744
rect 14941 15808 15257 15809
rect 14941 15744 14947 15808
rect 15011 15744 15027 15808
rect 15091 15744 15107 15808
rect 15171 15744 15187 15808
rect 15251 15744 15257 15808
rect 14941 15743 15257 15744
rect 20539 15808 20855 15809
rect 20539 15744 20545 15808
rect 20609 15744 20625 15808
rect 20689 15744 20705 15808
rect 20769 15744 20785 15808
rect 20849 15744 20855 15808
rect 20539 15743 20855 15744
rect 12249 15602 12315 15605
rect 17217 15602 17283 15605
rect 12249 15600 17283 15602
rect 12249 15544 12254 15600
rect 12310 15544 17222 15600
rect 17278 15544 17283 15600
rect 12249 15542 17283 15544
rect 12249 15539 12315 15542
rect 17217 15539 17283 15542
rect 17585 15602 17651 15605
rect 19701 15602 19767 15605
rect 23800 15602 24600 15632
rect 17585 15600 24600 15602
rect 17585 15544 17590 15600
rect 17646 15544 19706 15600
rect 19762 15544 24600 15600
rect 17585 15542 24600 15544
rect 17585 15539 17651 15542
rect 19701 15539 19767 15542
rect 23800 15512 24600 15542
rect 16665 15466 16731 15469
rect 23565 15466 23631 15469
rect 16665 15464 23631 15466
rect 16665 15408 16670 15464
rect 16726 15408 23570 15464
rect 23626 15408 23631 15464
rect 16665 15406 23631 15408
rect 16665 15403 16731 15406
rect 23565 15403 23631 15406
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 4245 15332 4311 15333
rect 4245 15328 4292 15332
rect 4356 15330 4362 15332
rect 4245 15272 4250 15328
rect 4245 15268 4292 15272
rect 4356 15270 4402 15330
rect 4356 15268 4362 15270
rect 4245 15267 4311 15268
rect 6544 15264 6860 15265
rect 6544 15200 6550 15264
rect 6614 15200 6630 15264
rect 6694 15200 6710 15264
rect 6774 15200 6790 15264
rect 6854 15200 6860 15264
rect 6544 15199 6860 15200
rect 12142 15264 12458 15265
rect 12142 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12458 15264
rect 12142 15199 12458 15200
rect 17740 15264 18056 15265
rect 17740 15200 17746 15264
rect 17810 15200 17826 15264
rect 17890 15200 17906 15264
rect 17970 15200 17986 15264
rect 18050 15200 18056 15264
rect 17740 15199 18056 15200
rect 16573 15196 16639 15197
rect 16573 15194 16620 15196
rect 16528 15192 16620 15194
rect 16528 15136 16578 15192
rect 16528 15134 16620 15136
rect 16573 15132 16620 15134
rect 16684 15132 16690 15196
rect 18781 15194 18847 15197
rect 21541 15194 21607 15197
rect 18781 15192 21607 15194
rect 18781 15136 18786 15192
rect 18842 15136 21546 15192
rect 21602 15136 21607 15192
rect 18781 15134 21607 15136
rect 16573 15131 16639 15132
rect 18781 15131 18847 15134
rect 21541 15131 21607 15134
rect 4889 15060 4955 15061
rect 4838 14996 4844 15060
rect 4908 15058 4955 15060
rect 19333 15058 19399 15061
rect 21725 15058 21791 15061
rect 4908 15056 5000 15058
rect 4950 15000 5000 15056
rect 4908 14998 5000 15000
rect 19333 15056 21791 15058
rect 19333 15000 19338 15056
rect 19394 15000 21730 15056
rect 21786 15000 21791 15056
rect 19333 14998 21791 15000
rect 4908 14996 4955 14998
rect 4889 14995 4955 14996
rect 19333 14995 19399 14998
rect 21725 14995 21791 14998
rect 22921 15058 22987 15061
rect 23800 15058 24600 15088
rect 22921 15056 24600 15058
rect 22921 15000 22926 15056
rect 22982 15000 24600 15056
rect 22921 14998 24600 15000
rect 22921 14995 22987 14998
rect 23800 14968 24600 14998
rect 19793 14922 19859 14925
rect 19793 14920 22110 14922
rect 19793 14864 19798 14920
rect 19854 14864 22110 14920
rect 19793 14862 22110 14864
rect 19793 14859 19859 14862
rect 3745 14720 4061 14721
rect 3745 14656 3751 14720
rect 3815 14656 3831 14720
rect 3895 14656 3911 14720
rect 3975 14656 3991 14720
rect 4055 14656 4061 14720
rect 3745 14655 4061 14656
rect 9343 14720 9659 14721
rect 9343 14656 9349 14720
rect 9413 14656 9429 14720
rect 9493 14656 9509 14720
rect 9573 14656 9589 14720
rect 9653 14656 9659 14720
rect 9343 14655 9659 14656
rect 14941 14720 15257 14721
rect 14941 14656 14947 14720
rect 15011 14656 15027 14720
rect 15091 14656 15107 14720
rect 15171 14656 15187 14720
rect 15251 14656 15257 14720
rect 14941 14655 15257 14656
rect 20539 14720 20855 14721
rect 20539 14656 20545 14720
rect 20609 14656 20625 14720
rect 20689 14656 20705 14720
rect 20769 14656 20785 14720
rect 20849 14656 20855 14720
rect 20539 14655 20855 14656
rect 15009 14514 15075 14517
rect 20253 14514 20319 14517
rect 15009 14512 20319 14514
rect 15009 14456 15014 14512
rect 15070 14456 20258 14512
rect 20314 14456 20319 14512
rect 15009 14454 20319 14456
rect 22050 14514 22110 14862
rect 23197 14514 23263 14517
rect 23800 14514 24600 14544
rect 22050 14512 24600 14514
rect 22050 14456 23202 14512
rect 23258 14456 24600 14512
rect 22050 14454 24600 14456
rect 15009 14451 15075 14454
rect 20253 14451 20319 14454
rect 23197 14451 23263 14454
rect 23800 14424 24600 14454
rect 13261 14378 13327 14381
rect 21357 14378 21423 14381
rect 13261 14376 21423 14378
rect 13261 14320 13266 14376
rect 13322 14320 21362 14376
rect 21418 14320 21423 14376
rect 13261 14318 21423 14320
rect 13261 14315 13327 14318
rect 21357 14315 21423 14318
rect 16481 14242 16547 14245
rect 17166 14242 17172 14244
rect 16481 14240 17172 14242
rect 16481 14184 16486 14240
rect 16542 14184 17172 14240
rect 16481 14182 17172 14184
rect 16481 14179 16547 14182
rect 17166 14180 17172 14182
rect 17236 14180 17242 14244
rect 6544 14176 6860 14177
rect 6544 14112 6550 14176
rect 6614 14112 6630 14176
rect 6694 14112 6710 14176
rect 6774 14112 6790 14176
rect 6854 14112 6860 14176
rect 6544 14111 6860 14112
rect 12142 14176 12458 14177
rect 12142 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12458 14176
rect 12142 14111 12458 14112
rect 17740 14176 18056 14177
rect 17740 14112 17746 14176
rect 17810 14112 17826 14176
rect 17890 14112 17906 14176
rect 17970 14112 17986 14176
rect 18050 14112 18056 14176
rect 17740 14111 18056 14112
rect 15193 13970 15259 13973
rect 19701 13970 19767 13973
rect 15193 13968 19767 13970
rect 15193 13912 15198 13968
rect 15254 13912 19706 13968
rect 19762 13912 19767 13968
rect 15193 13910 19767 13912
rect 15193 13907 15259 13910
rect 19701 13907 19767 13910
rect 21725 13970 21791 13973
rect 23800 13970 24600 14000
rect 21725 13968 24600 13970
rect 21725 13912 21730 13968
rect 21786 13912 24600 13968
rect 21725 13910 24600 13912
rect 21725 13907 21791 13910
rect 23800 13880 24600 13910
rect 3745 13632 4061 13633
rect 3745 13568 3751 13632
rect 3815 13568 3831 13632
rect 3895 13568 3911 13632
rect 3975 13568 3991 13632
rect 4055 13568 4061 13632
rect 3745 13567 4061 13568
rect 9343 13632 9659 13633
rect 9343 13568 9349 13632
rect 9413 13568 9429 13632
rect 9493 13568 9509 13632
rect 9573 13568 9589 13632
rect 9653 13568 9659 13632
rect 9343 13567 9659 13568
rect 14941 13632 15257 13633
rect 14941 13568 14947 13632
rect 15011 13568 15027 13632
rect 15091 13568 15107 13632
rect 15171 13568 15187 13632
rect 15251 13568 15257 13632
rect 14941 13567 15257 13568
rect 20539 13632 20855 13633
rect 20539 13568 20545 13632
rect 20609 13568 20625 13632
rect 20689 13568 20705 13632
rect 20769 13568 20785 13632
rect 20849 13568 20855 13632
rect 20539 13567 20855 13568
rect 5349 13426 5415 13429
rect 5574 13426 5580 13428
rect 5349 13424 5580 13426
rect 5349 13368 5354 13424
rect 5410 13368 5580 13424
rect 5349 13366 5580 13368
rect 5349 13363 5415 13366
rect 5574 13364 5580 13366
rect 5644 13364 5650 13428
rect 15101 13426 15167 13429
rect 18270 13426 18276 13428
rect 15101 13424 18276 13426
rect 15101 13368 15106 13424
rect 15162 13368 18276 13424
rect 15101 13366 18276 13368
rect 15101 13363 15167 13366
rect 18270 13364 18276 13366
rect 18340 13364 18346 13428
rect 19333 13426 19399 13429
rect 23800 13426 24600 13456
rect 19333 13424 24600 13426
rect 19333 13368 19338 13424
rect 19394 13368 24600 13424
rect 19333 13366 24600 13368
rect 19333 13363 19399 13366
rect 23800 13336 24600 13366
rect 14641 13290 14707 13293
rect 21081 13290 21147 13293
rect 14641 13288 21147 13290
rect 14641 13232 14646 13288
rect 14702 13232 21086 13288
rect 21142 13232 21147 13288
rect 14641 13230 21147 13232
rect 14641 13227 14707 13230
rect 21081 13227 21147 13230
rect 19425 13154 19491 13157
rect 19425 13152 22110 13154
rect 19425 13096 19430 13152
rect 19486 13096 22110 13152
rect 19425 13094 22110 13096
rect 19425 13091 19491 13094
rect 6544 13088 6860 13089
rect 6544 13024 6550 13088
rect 6614 13024 6630 13088
rect 6694 13024 6710 13088
rect 6774 13024 6790 13088
rect 6854 13024 6860 13088
rect 6544 13023 6860 13024
rect 12142 13088 12458 13089
rect 12142 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12458 13088
rect 12142 13023 12458 13024
rect 17740 13088 18056 13089
rect 17740 13024 17746 13088
rect 17810 13024 17826 13088
rect 17890 13024 17906 13088
rect 17970 13024 17986 13088
rect 18050 13024 18056 13088
rect 17740 13023 18056 13024
rect 18321 13018 18387 13021
rect 21081 13018 21147 13021
rect 18321 13016 21147 13018
rect 18321 12960 18326 13016
rect 18382 12960 21086 13016
rect 21142 12960 21147 13016
rect 18321 12958 21147 12960
rect 18321 12955 18387 12958
rect 21081 12955 21147 12958
rect 4153 12882 4219 12885
rect 4286 12882 4292 12884
rect 4153 12880 4292 12882
rect 4153 12824 4158 12880
rect 4214 12824 4292 12880
rect 4153 12822 4292 12824
rect 4153 12819 4219 12822
rect 4286 12820 4292 12822
rect 4356 12820 4362 12884
rect 19057 12882 19123 12885
rect 21173 12882 21239 12885
rect 19057 12880 21239 12882
rect 19057 12824 19062 12880
rect 19118 12824 21178 12880
rect 21234 12824 21239 12880
rect 19057 12822 21239 12824
rect 22050 12882 22110 13094
rect 23800 12882 24600 12912
rect 22050 12822 24600 12882
rect 19057 12819 19123 12822
rect 21173 12819 21239 12822
rect 23800 12792 24600 12822
rect 11053 12746 11119 12749
rect 18822 12746 18828 12748
rect 11053 12744 18828 12746
rect 11053 12688 11058 12744
rect 11114 12688 18828 12744
rect 11053 12686 18828 12688
rect 11053 12683 11119 12686
rect 18822 12684 18828 12686
rect 18892 12684 18898 12748
rect 19057 12746 19123 12749
rect 21265 12746 21331 12749
rect 19057 12744 21331 12746
rect 19057 12688 19062 12744
rect 19118 12688 21270 12744
rect 21326 12688 21331 12744
rect 19057 12686 21331 12688
rect 19057 12683 19123 12686
rect 21265 12683 21331 12686
rect 3745 12544 4061 12545
rect 3745 12480 3751 12544
rect 3815 12480 3831 12544
rect 3895 12480 3911 12544
rect 3975 12480 3991 12544
rect 4055 12480 4061 12544
rect 3745 12479 4061 12480
rect 9343 12544 9659 12545
rect 9343 12480 9349 12544
rect 9413 12480 9429 12544
rect 9493 12480 9509 12544
rect 9573 12480 9589 12544
rect 9653 12480 9659 12544
rect 9343 12479 9659 12480
rect 14941 12544 15257 12545
rect 14941 12480 14947 12544
rect 15011 12480 15027 12544
rect 15091 12480 15107 12544
rect 15171 12480 15187 12544
rect 15251 12480 15257 12544
rect 14941 12479 15257 12480
rect 20539 12544 20855 12545
rect 20539 12480 20545 12544
rect 20609 12480 20625 12544
rect 20689 12480 20705 12544
rect 20769 12480 20785 12544
rect 20849 12480 20855 12544
rect 20539 12479 20855 12480
rect 11697 12338 11763 12341
rect 18454 12338 18460 12340
rect 11697 12336 18460 12338
rect 11697 12280 11702 12336
rect 11758 12280 18460 12336
rect 11697 12278 18460 12280
rect 11697 12275 11763 12278
rect 18454 12276 18460 12278
rect 18524 12276 18530 12340
rect 19333 12338 19399 12341
rect 23800 12338 24600 12368
rect 19333 12336 24600 12338
rect 19333 12280 19338 12336
rect 19394 12280 24600 12336
rect 19333 12278 24600 12280
rect 19333 12275 19399 12278
rect 23800 12248 24600 12278
rect 17953 12202 18019 12205
rect 22645 12202 22711 12205
rect 17953 12200 22711 12202
rect 17953 12144 17958 12200
rect 18014 12144 22650 12200
rect 22706 12144 22711 12200
rect 17953 12142 22711 12144
rect 17953 12139 18019 12142
rect 22645 12139 22711 12142
rect 20989 12066 21055 12069
rect 22737 12066 22803 12069
rect 20989 12064 22803 12066
rect 20989 12008 20994 12064
rect 21050 12008 22742 12064
rect 22798 12008 22803 12064
rect 20989 12006 22803 12008
rect 20989 12003 21055 12006
rect 22737 12003 22803 12006
rect 6544 12000 6860 12001
rect 6544 11936 6550 12000
rect 6614 11936 6630 12000
rect 6694 11936 6710 12000
rect 6774 11936 6790 12000
rect 6854 11936 6860 12000
rect 6544 11935 6860 11936
rect 12142 12000 12458 12001
rect 12142 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12458 12000
rect 12142 11935 12458 11936
rect 17740 12000 18056 12001
rect 17740 11936 17746 12000
rect 17810 11936 17826 12000
rect 17890 11936 17906 12000
rect 17970 11936 17986 12000
rect 18050 11936 18056 12000
rect 17740 11935 18056 11936
rect 19793 11930 19859 11933
rect 22829 11930 22895 11933
rect 19793 11928 22895 11930
rect 19793 11872 19798 11928
rect 19854 11872 22834 11928
rect 22890 11872 22895 11928
rect 19793 11870 22895 11872
rect 19793 11867 19859 11870
rect 22829 11867 22895 11870
rect 3877 11794 3943 11797
rect 6310 11794 6316 11796
rect 3877 11792 6316 11794
rect 3877 11736 3882 11792
rect 3938 11736 6316 11792
rect 3877 11734 6316 11736
rect 3877 11731 3943 11734
rect 6310 11732 6316 11734
rect 6380 11732 6386 11796
rect 18321 11794 18387 11797
rect 23800 11794 24600 11824
rect 18321 11792 24600 11794
rect 18321 11736 18326 11792
rect 18382 11736 24600 11792
rect 18321 11734 24600 11736
rect 18321 11731 18387 11734
rect 23800 11704 24600 11734
rect 19977 11658 20043 11661
rect 21633 11658 21699 11661
rect 19977 11656 21699 11658
rect 19977 11600 19982 11656
rect 20038 11600 21638 11656
rect 21694 11600 21699 11656
rect 19977 11598 21699 11600
rect 19977 11595 20043 11598
rect 21633 11595 21699 11598
rect 3745 11456 4061 11457
rect 3745 11392 3751 11456
rect 3815 11392 3831 11456
rect 3895 11392 3911 11456
rect 3975 11392 3991 11456
rect 4055 11392 4061 11456
rect 3745 11391 4061 11392
rect 9343 11456 9659 11457
rect 9343 11392 9349 11456
rect 9413 11392 9429 11456
rect 9493 11392 9509 11456
rect 9573 11392 9589 11456
rect 9653 11392 9659 11456
rect 9343 11391 9659 11392
rect 14941 11456 15257 11457
rect 14941 11392 14947 11456
rect 15011 11392 15027 11456
rect 15091 11392 15107 11456
rect 15171 11392 15187 11456
rect 15251 11392 15257 11456
rect 14941 11391 15257 11392
rect 20539 11456 20855 11457
rect 20539 11392 20545 11456
rect 20609 11392 20625 11456
rect 20689 11392 20705 11456
rect 20769 11392 20785 11456
rect 20849 11392 20855 11456
rect 20539 11391 20855 11392
rect 18137 11250 18203 11253
rect 19190 11250 19196 11252
rect 18137 11248 19196 11250
rect 18137 11192 18142 11248
rect 18198 11192 19196 11248
rect 18137 11190 19196 11192
rect 18137 11187 18203 11190
rect 19190 11188 19196 11190
rect 19260 11188 19266 11252
rect 19333 11250 19399 11253
rect 23800 11250 24600 11280
rect 19333 11248 24600 11250
rect 19333 11192 19338 11248
rect 19394 11192 24600 11248
rect 19333 11190 24600 11192
rect 19333 11187 19399 11190
rect 23800 11160 24600 11190
rect 18045 11114 18111 11117
rect 20897 11114 20963 11117
rect 18045 11112 20963 11114
rect 18045 11056 18050 11112
rect 18106 11056 20902 11112
rect 20958 11056 20963 11112
rect 18045 11054 20963 11056
rect 18045 11051 18111 11054
rect 20897 11051 20963 11054
rect 6544 10912 6860 10913
rect 6544 10848 6550 10912
rect 6614 10848 6630 10912
rect 6694 10848 6710 10912
rect 6774 10848 6790 10912
rect 6854 10848 6860 10912
rect 6544 10847 6860 10848
rect 12142 10912 12458 10913
rect 12142 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12458 10912
rect 12142 10847 12458 10848
rect 17740 10912 18056 10913
rect 17740 10848 17746 10912
rect 17810 10848 17826 10912
rect 17890 10848 17906 10912
rect 17970 10848 17986 10912
rect 18050 10848 18056 10912
rect 17740 10847 18056 10848
rect 19333 10842 19399 10845
rect 19333 10840 23122 10842
rect 19333 10784 19338 10840
rect 19394 10784 23122 10840
rect 19333 10782 23122 10784
rect 19333 10779 19399 10782
rect 15469 10706 15535 10709
rect 22093 10706 22159 10709
rect 15469 10704 22159 10706
rect 15469 10648 15474 10704
rect 15530 10648 22098 10704
rect 22154 10648 22159 10704
rect 15469 10646 22159 10648
rect 23062 10706 23122 10782
rect 23800 10706 24600 10736
rect 23062 10646 24600 10706
rect 15469 10643 15535 10646
rect 22093 10643 22159 10646
rect 23800 10616 24600 10646
rect 6821 10570 6887 10573
rect 8109 10570 8175 10573
rect 6821 10568 8175 10570
rect 6821 10512 6826 10568
rect 6882 10512 8114 10568
rect 8170 10512 8175 10568
rect 6821 10510 8175 10512
rect 6821 10507 6887 10510
rect 8109 10507 8175 10510
rect 3745 10368 4061 10369
rect 3745 10304 3751 10368
rect 3815 10304 3831 10368
rect 3895 10304 3911 10368
rect 3975 10304 3991 10368
rect 4055 10304 4061 10368
rect 3745 10303 4061 10304
rect 9343 10368 9659 10369
rect 9343 10304 9349 10368
rect 9413 10304 9429 10368
rect 9493 10304 9509 10368
rect 9573 10304 9589 10368
rect 9653 10304 9659 10368
rect 9343 10303 9659 10304
rect 14941 10368 15257 10369
rect 14941 10304 14947 10368
rect 15011 10304 15027 10368
rect 15091 10304 15107 10368
rect 15171 10304 15187 10368
rect 15251 10304 15257 10368
rect 14941 10303 15257 10304
rect 20539 10368 20855 10369
rect 20539 10304 20545 10368
rect 20609 10304 20625 10368
rect 20689 10304 20705 10368
rect 20769 10304 20785 10368
rect 20849 10304 20855 10368
rect 20539 10303 20855 10304
rect 19241 10162 19307 10165
rect 20713 10162 20779 10165
rect 21909 10162 21975 10165
rect 23800 10162 24600 10192
rect 19241 10160 21975 10162
rect 19241 10104 19246 10160
rect 19302 10104 20718 10160
rect 20774 10104 21914 10160
rect 21970 10104 21975 10160
rect 19241 10102 21975 10104
rect 19241 10099 19307 10102
rect 20713 10099 20779 10102
rect 21909 10099 21975 10102
rect 23062 10102 24600 10162
rect 16941 10026 17007 10029
rect 22829 10026 22895 10029
rect 16941 10024 22895 10026
rect 16941 9968 16946 10024
rect 17002 9968 22834 10024
rect 22890 9968 22895 10024
rect 16941 9966 22895 9968
rect 16941 9963 17007 9966
rect 22829 9963 22895 9966
rect 19333 9890 19399 9893
rect 23062 9890 23122 10102
rect 23800 10072 24600 10102
rect 19333 9888 23122 9890
rect 19333 9832 19338 9888
rect 19394 9832 23122 9888
rect 19333 9830 23122 9832
rect 19333 9827 19399 9830
rect 6544 9824 6860 9825
rect 6544 9760 6550 9824
rect 6614 9760 6630 9824
rect 6694 9760 6710 9824
rect 6774 9760 6790 9824
rect 6854 9760 6860 9824
rect 6544 9759 6860 9760
rect 12142 9824 12458 9825
rect 12142 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12458 9824
rect 12142 9759 12458 9760
rect 17740 9824 18056 9825
rect 17740 9760 17746 9824
rect 17810 9760 17826 9824
rect 17890 9760 17906 9824
rect 17970 9760 17986 9824
rect 18050 9760 18056 9824
rect 17740 9759 18056 9760
rect 18321 9754 18387 9757
rect 19701 9754 19767 9757
rect 18321 9752 19767 9754
rect 18321 9696 18326 9752
rect 18382 9696 19706 9752
rect 19762 9696 19767 9752
rect 18321 9694 19767 9696
rect 18321 9691 18387 9694
rect 19701 9691 19767 9694
rect 17769 9618 17835 9621
rect 20989 9618 21055 9621
rect 17769 9616 21055 9618
rect 17769 9560 17774 9616
rect 17830 9560 20994 9616
rect 21050 9560 21055 9616
rect 17769 9558 21055 9560
rect 17769 9555 17835 9558
rect 20989 9555 21055 9558
rect 21265 9618 21331 9621
rect 22737 9618 22803 9621
rect 23800 9618 24600 9648
rect 21265 9616 22803 9618
rect 21265 9560 21270 9616
rect 21326 9560 22742 9616
rect 22798 9560 22803 9616
rect 21265 9558 22803 9560
rect 21265 9555 21331 9558
rect 22737 9555 22803 9558
rect 23062 9558 24600 9618
rect 17585 9482 17651 9485
rect 22553 9482 22619 9485
rect 17585 9480 22619 9482
rect 17585 9424 17590 9480
rect 17646 9424 22558 9480
rect 22614 9424 22619 9480
rect 17585 9422 22619 9424
rect 17585 9419 17651 9422
rect 22553 9419 22619 9422
rect 20989 9346 21055 9349
rect 23062 9346 23122 9558
rect 23800 9528 24600 9558
rect 20989 9344 23122 9346
rect 20989 9288 20994 9344
rect 21050 9288 23122 9344
rect 20989 9286 23122 9288
rect 20989 9283 21055 9286
rect 3745 9280 4061 9281
rect 0 9210 800 9240
rect 3745 9216 3751 9280
rect 3815 9216 3831 9280
rect 3895 9216 3911 9280
rect 3975 9216 3991 9280
rect 4055 9216 4061 9280
rect 3745 9215 4061 9216
rect 9343 9280 9659 9281
rect 9343 9216 9349 9280
rect 9413 9216 9429 9280
rect 9493 9216 9509 9280
rect 9573 9216 9589 9280
rect 9653 9216 9659 9280
rect 9343 9215 9659 9216
rect 14941 9280 15257 9281
rect 14941 9216 14947 9280
rect 15011 9216 15027 9280
rect 15091 9216 15107 9280
rect 15171 9216 15187 9280
rect 15251 9216 15257 9280
rect 14941 9215 15257 9216
rect 20539 9280 20855 9281
rect 20539 9216 20545 9280
rect 20609 9216 20625 9280
rect 20689 9216 20705 9280
rect 20769 9216 20785 9280
rect 20849 9216 20855 9280
rect 20539 9215 20855 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 19333 9074 19399 9077
rect 23800 9074 24600 9104
rect 19333 9072 24600 9074
rect 19333 9016 19338 9072
rect 19394 9016 24600 9072
rect 19333 9014 24600 9016
rect 19333 9011 19399 9014
rect 23800 8984 24600 9014
rect 17125 8938 17191 8941
rect 21817 8938 21883 8941
rect 17125 8936 21883 8938
rect 17125 8880 17130 8936
rect 17186 8880 21822 8936
rect 21878 8880 21883 8936
rect 17125 8878 21883 8880
rect 17125 8875 17191 8878
rect 21817 8875 21883 8878
rect 19006 8740 19012 8804
rect 19076 8802 19082 8804
rect 19149 8802 19215 8805
rect 19076 8800 19215 8802
rect 19076 8744 19154 8800
rect 19210 8744 19215 8800
rect 19076 8742 19215 8744
rect 19076 8740 19082 8742
rect 19149 8739 19215 8742
rect 6544 8736 6860 8737
rect 6544 8672 6550 8736
rect 6614 8672 6630 8736
rect 6694 8672 6710 8736
rect 6774 8672 6790 8736
rect 6854 8672 6860 8736
rect 6544 8671 6860 8672
rect 12142 8736 12458 8737
rect 12142 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12458 8736
rect 12142 8671 12458 8672
rect 17740 8736 18056 8737
rect 17740 8672 17746 8736
rect 17810 8672 17826 8736
rect 17890 8672 17906 8736
rect 17970 8672 17986 8736
rect 18050 8672 18056 8736
rect 17740 8671 18056 8672
rect 19517 8666 19583 8669
rect 23289 8666 23355 8669
rect 19517 8664 23355 8666
rect 19517 8608 19522 8664
rect 19578 8608 23294 8664
rect 23350 8608 23355 8664
rect 19517 8606 23355 8608
rect 19517 8603 19583 8606
rect 23289 8603 23355 8606
rect 19333 8530 19399 8533
rect 16622 8528 19399 8530
rect 16622 8472 19338 8528
rect 19394 8472 19399 8528
rect 16622 8470 19399 8472
rect 15929 8394 15995 8397
rect 16622 8396 16682 8470
rect 19333 8467 19399 8470
rect 20161 8530 20227 8533
rect 20529 8530 20595 8533
rect 20161 8528 20595 8530
rect 20161 8472 20166 8528
rect 20222 8472 20534 8528
rect 20590 8472 20595 8528
rect 20161 8470 20595 8472
rect 20161 8467 20227 8470
rect 20529 8467 20595 8470
rect 23105 8530 23171 8533
rect 23800 8530 24600 8560
rect 23105 8528 24600 8530
rect 23105 8472 23110 8528
rect 23166 8472 24600 8528
rect 23105 8470 24600 8472
rect 23105 8467 23171 8470
rect 23800 8440 24600 8470
rect 16614 8394 16620 8396
rect 15929 8392 16620 8394
rect 15929 8336 15934 8392
rect 15990 8336 16620 8392
rect 15929 8334 16620 8336
rect 15929 8331 15995 8334
rect 16614 8332 16620 8334
rect 16684 8332 16690 8396
rect 17309 8394 17375 8397
rect 23657 8394 23723 8397
rect 17309 8392 23723 8394
rect 17309 8336 17314 8392
rect 17370 8336 23662 8392
rect 23718 8336 23723 8392
rect 17309 8334 23723 8336
rect 17309 8331 17375 8334
rect 23657 8331 23723 8334
rect 3745 8192 4061 8193
rect 3745 8128 3751 8192
rect 3815 8128 3831 8192
rect 3895 8128 3911 8192
rect 3975 8128 3991 8192
rect 4055 8128 4061 8192
rect 3745 8127 4061 8128
rect 9343 8192 9659 8193
rect 9343 8128 9349 8192
rect 9413 8128 9429 8192
rect 9493 8128 9509 8192
rect 9573 8128 9589 8192
rect 9653 8128 9659 8192
rect 9343 8127 9659 8128
rect 14941 8192 15257 8193
rect 14941 8128 14947 8192
rect 15011 8128 15027 8192
rect 15091 8128 15107 8192
rect 15171 8128 15187 8192
rect 15251 8128 15257 8192
rect 14941 8127 15257 8128
rect 20539 8192 20855 8193
rect 20539 8128 20545 8192
rect 20609 8128 20625 8192
rect 20689 8128 20705 8192
rect 20769 8128 20785 8192
rect 20849 8128 20855 8192
rect 20539 8127 20855 8128
rect 18321 7986 18387 7989
rect 21817 7986 21883 7989
rect 18321 7984 21883 7986
rect 18321 7928 18326 7984
rect 18382 7928 21822 7984
rect 21878 7928 21883 7984
rect 18321 7926 21883 7928
rect 18321 7923 18387 7926
rect 21817 7923 21883 7926
rect 22001 7986 22067 7989
rect 23800 7986 24600 8016
rect 22001 7984 24600 7986
rect 22001 7928 22006 7984
rect 22062 7928 24600 7984
rect 22001 7926 24600 7928
rect 22001 7923 22067 7926
rect 23800 7896 24600 7926
rect 12065 7850 12131 7853
rect 20069 7850 20135 7853
rect 12065 7848 20135 7850
rect 12065 7792 12070 7848
rect 12126 7792 20074 7848
rect 20130 7792 20135 7848
rect 12065 7790 20135 7792
rect 12065 7787 12131 7790
rect 20069 7787 20135 7790
rect 20294 7788 20300 7852
rect 20364 7850 20370 7852
rect 22093 7850 22159 7853
rect 20364 7848 22159 7850
rect 20364 7792 22098 7848
rect 22154 7792 22159 7848
rect 20364 7790 22159 7792
rect 20364 7788 20370 7790
rect 22093 7787 22159 7790
rect 19885 7714 19951 7717
rect 20437 7714 20503 7717
rect 19885 7712 20503 7714
rect 19885 7656 19890 7712
rect 19946 7656 20442 7712
rect 20498 7656 20503 7712
rect 19885 7654 20503 7656
rect 19885 7651 19951 7654
rect 20437 7651 20503 7654
rect 20805 7714 20871 7717
rect 21030 7714 21036 7716
rect 20805 7712 21036 7714
rect 20805 7656 20810 7712
rect 20866 7656 21036 7712
rect 20805 7654 21036 7656
rect 20805 7651 20871 7654
rect 21030 7652 21036 7654
rect 21100 7652 21106 7716
rect 6544 7648 6860 7649
rect 6544 7584 6550 7648
rect 6614 7584 6630 7648
rect 6694 7584 6710 7648
rect 6774 7584 6790 7648
rect 6854 7584 6860 7648
rect 6544 7583 6860 7584
rect 12142 7648 12458 7649
rect 12142 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12458 7648
rect 12142 7583 12458 7584
rect 17740 7648 18056 7649
rect 17740 7584 17746 7648
rect 17810 7584 17826 7648
rect 17890 7584 17906 7648
rect 17970 7584 17986 7648
rect 18050 7584 18056 7648
rect 17740 7583 18056 7584
rect 18505 7578 18571 7581
rect 22829 7578 22895 7581
rect 18505 7576 22895 7578
rect 18505 7520 18510 7576
rect 18566 7520 22834 7576
rect 22890 7520 22895 7576
rect 18505 7518 22895 7520
rect 18505 7515 18571 7518
rect 22829 7515 22895 7518
rect 13537 7442 13603 7445
rect 19701 7442 19767 7445
rect 13537 7440 19767 7442
rect 13537 7384 13542 7440
rect 13598 7384 19706 7440
rect 19762 7384 19767 7440
rect 13537 7382 19767 7384
rect 13537 7379 13603 7382
rect 19701 7379 19767 7382
rect 21449 7442 21515 7445
rect 23800 7442 24600 7472
rect 21449 7440 24600 7442
rect 21449 7384 21454 7440
rect 21510 7384 24600 7440
rect 21449 7382 24600 7384
rect 21449 7379 21515 7382
rect 23800 7352 24600 7382
rect 10777 7306 10843 7309
rect 18137 7306 18203 7309
rect 22737 7306 22803 7309
rect 10777 7304 15394 7306
rect 10777 7248 10782 7304
rect 10838 7248 15394 7304
rect 10777 7246 15394 7248
rect 10777 7243 10843 7246
rect 15334 7170 15394 7246
rect 18137 7304 22803 7306
rect 18137 7248 18142 7304
rect 18198 7248 22742 7304
rect 22798 7248 22803 7304
rect 18137 7246 22803 7248
rect 18137 7243 18203 7246
rect 22737 7243 22803 7246
rect 19057 7170 19123 7173
rect 15334 7168 19123 7170
rect 15334 7112 19062 7168
rect 19118 7112 19123 7168
rect 15334 7110 19123 7112
rect 19057 7107 19123 7110
rect 19333 7170 19399 7173
rect 19609 7170 19675 7173
rect 21449 7172 21515 7173
rect 19333 7168 19675 7170
rect 19333 7112 19338 7168
rect 19394 7112 19614 7168
rect 19670 7112 19675 7168
rect 19333 7110 19675 7112
rect 19333 7107 19399 7110
rect 19609 7107 19675 7110
rect 21398 7108 21404 7172
rect 21468 7170 21515 7172
rect 21468 7168 21560 7170
rect 21510 7112 21560 7168
rect 21468 7110 21560 7112
rect 21468 7108 21515 7110
rect 21449 7107 21515 7108
rect 3745 7104 4061 7105
rect 3745 7040 3751 7104
rect 3815 7040 3831 7104
rect 3895 7040 3911 7104
rect 3975 7040 3991 7104
rect 4055 7040 4061 7104
rect 3745 7039 4061 7040
rect 9343 7104 9659 7105
rect 9343 7040 9349 7104
rect 9413 7040 9429 7104
rect 9493 7040 9509 7104
rect 9573 7040 9589 7104
rect 9653 7040 9659 7104
rect 9343 7039 9659 7040
rect 14941 7104 15257 7105
rect 14941 7040 14947 7104
rect 15011 7040 15027 7104
rect 15091 7040 15107 7104
rect 15171 7040 15187 7104
rect 15251 7040 15257 7104
rect 14941 7039 15257 7040
rect 20539 7104 20855 7105
rect 20539 7040 20545 7104
rect 20609 7040 20625 7104
rect 20689 7040 20705 7104
rect 20769 7040 20785 7104
rect 20849 7040 20855 7104
rect 20539 7039 20855 7040
rect 18638 6972 18644 7036
rect 18708 7034 18714 7036
rect 19149 7034 19215 7037
rect 18708 7032 19215 7034
rect 18708 6976 19154 7032
rect 19210 6976 19215 7032
rect 18708 6974 19215 6976
rect 18708 6972 18714 6974
rect 19149 6971 19215 6974
rect 22134 6972 22140 7036
rect 22204 7034 22210 7036
rect 22277 7034 22343 7037
rect 22204 7032 22343 7034
rect 22204 6976 22282 7032
rect 22338 6976 22343 7032
rect 22204 6974 22343 6976
rect 22204 6972 22210 6974
rect 22277 6971 22343 6974
rect 10685 6898 10751 6901
rect 22645 6898 22711 6901
rect 10685 6896 22711 6898
rect 10685 6840 10690 6896
rect 10746 6840 22650 6896
rect 22706 6840 22711 6896
rect 10685 6838 22711 6840
rect 10685 6835 10751 6838
rect 22645 6835 22711 6838
rect 23105 6898 23171 6901
rect 23800 6898 24600 6928
rect 23105 6896 24600 6898
rect 23105 6840 23110 6896
rect 23166 6840 24600 6896
rect 23105 6838 24600 6840
rect 23105 6835 23171 6838
rect 23800 6808 24600 6838
rect 15193 6762 15259 6765
rect 20897 6762 20963 6765
rect 15193 6760 20963 6762
rect 15193 6704 15198 6760
rect 15254 6704 20902 6760
rect 20958 6704 20963 6760
rect 15193 6702 20963 6704
rect 15193 6699 15259 6702
rect 20897 6699 20963 6702
rect 18137 6626 18203 6629
rect 20897 6626 20963 6629
rect 21817 6626 21883 6629
rect 18137 6624 21883 6626
rect 18137 6568 18142 6624
rect 18198 6568 20902 6624
rect 20958 6568 21822 6624
rect 21878 6568 21883 6624
rect 18137 6566 21883 6568
rect 18137 6563 18203 6566
rect 20897 6563 20963 6566
rect 21817 6563 21883 6566
rect 22185 6624 22251 6629
rect 22185 6568 22190 6624
rect 22246 6568 22251 6624
rect 22185 6563 22251 6568
rect 6544 6560 6860 6561
rect 6544 6496 6550 6560
rect 6614 6496 6630 6560
rect 6694 6496 6710 6560
rect 6774 6496 6790 6560
rect 6854 6496 6860 6560
rect 6544 6495 6860 6496
rect 12142 6560 12458 6561
rect 12142 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12458 6560
rect 12142 6495 12458 6496
rect 17740 6560 18056 6561
rect 17740 6496 17746 6560
rect 17810 6496 17826 6560
rect 17890 6496 17906 6560
rect 17970 6496 17986 6560
rect 18050 6496 18056 6560
rect 17740 6495 18056 6496
rect 19425 6490 19491 6493
rect 20294 6490 20300 6492
rect 19425 6488 20300 6490
rect 19425 6432 19430 6488
rect 19486 6432 20300 6488
rect 19425 6430 20300 6432
rect 19425 6427 19491 6430
rect 20294 6428 20300 6430
rect 20364 6490 20370 6492
rect 20437 6490 20503 6493
rect 20364 6488 20503 6490
rect 20364 6432 20442 6488
rect 20498 6432 20503 6488
rect 20364 6430 20503 6432
rect 20364 6428 20370 6430
rect 20437 6427 20503 6430
rect 20621 6490 20687 6493
rect 22188 6490 22248 6563
rect 20621 6488 22248 6490
rect 20621 6432 20626 6488
rect 20682 6432 22248 6488
rect 20621 6430 22248 6432
rect 20621 6427 20687 6430
rect 15837 6354 15903 6357
rect 16021 6354 16087 6357
rect 20253 6354 20319 6357
rect 15837 6352 20319 6354
rect 15837 6296 15842 6352
rect 15898 6296 16026 6352
rect 16082 6296 20258 6352
rect 20314 6296 20319 6352
rect 15837 6294 20319 6296
rect 15837 6291 15903 6294
rect 16021 6291 16087 6294
rect 20253 6291 20319 6294
rect 21398 6292 21404 6356
rect 21468 6354 21474 6356
rect 21541 6354 21607 6357
rect 21468 6352 21607 6354
rect 21468 6296 21546 6352
rect 21602 6296 21607 6352
rect 21468 6294 21607 6296
rect 21468 6292 21474 6294
rect 21541 6291 21607 6294
rect 22277 6354 22343 6357
rect 22461 6354 22527 6357
rect 22277 6352 22527 6354
rect 22277 6296 22282 6352
rect 22338 6296 22466 6352
rect 22522 6296 22527 6352
rect 22277 6294 22527 6296
rect 22277 6291 22343 6294
rect 22461 6291 22527 6294
rect 23013 6354 23079 6357
rect 23800 6354 24600 6384
rect 23013 6352 24600 6354
rect 23013 6296 23018 6352
rect 23074 6296 24600 6352
rect 23013 6294 24600 6296
rect 23013 6291 23079 6294
rect 23800 6264 24600 6294
rect 12801 6218 12867 6221
rect 19977 6218 20043 6221
rect 22185 6218 22251 6221
rect 12801 6216 18890 6218
rect 12801 6160 12806 6216
rect 12862 6160 18890 6216
rect 12801 6158 18890 6160
rect 12801 6155 12867 6158
rect 18830 6082 18890 6158
rect 19977 6216 22251 6218
rect 19977 6160 19982 6216
rect 20038 6160 22190 6216
rect 22246 6160 22251 6216
rect 19977 6158 22251 6160
rect 19977 6155 20043 6158
rect 22185 6155 22251 6158
rect 18965 6082 19031 6085
rect 18830 6080 19031 6082
rect 18830 6024 18970 6080
rect 19026 6024 19031 6080
rect 18830 6022 19031 6024
rect 18965 6019 19031 6022
rect 22093 6082 22159 6085
rect 22369 6082 22435 6085
rect 22093 6080 22435 6082
rect 22093 6024 22098 6080
rect 22154 6024 22374 6080
rect 22430 6024 22435 6080
rect 22093 6022 22435 6024
rect 22093 6019 22159 6022
rect 22369 6019 22435 6022
rect 3745 6016 4061 6017
rect 3745 5952 3751 6016
rect 3815 5952 3831 6016
rect 3895 5952 3911 6016
rect 3975 5952 3991 6016
rect 4055 5952 4061 6016
rect 3745 5951 4061 5952
rect 9343 6016 9659 6017
rect 9343 5952 9349 6016
rect 9413 5952 9429 6016
rect 9493 5952 9509 6016
rect 9573 5952 9589 6016
rect 9653 5952 9659 6016
rect 9343 5951 9659 5952
rect 14941 6016 15257 6017
rect 14941 5952 14947 6016
rect 15011 5952 15027 6016
rect 15091 5952 15107 6016
rect 15171 5952 15187 6016
rect 15251 5952 15257 6016
rect 14941 5951 15257 5952
rect 20539 6016 20855 6017
rect 20539 5952 20545 6016
rect 20609 5952 20625 6016
rect 20689 5952 20705 6016
rect 20769 5952 20785 6016
rect 20849 5952 20855 6016
rect 20539 5951 20855 5952
rect 18638 5884 18644 5948
rect 18708 5946 18714 5948
rect 19057 5946 19123 5949
rect 18708 5944 19123 5946
rect 18708 5888 19062 5944
rect 19118 5888 19123 5944
rect 18708 5886 19123 5888
rect 18708 5884 18714 5886
rect 19057 5883 19123 5886
rect 21909 5946 21975 5949
rect 22134 5946 22140 5948
rect 21909 5944 22140 5946
rect 21909 5888 21914 5944
rect 21970 5888 22140 5944
rect 21909 5886 22140 5888
rect 21909 5883 21975 5886
rect 22134 5884 22140 5886
rect 22204 5884 22210 5948
rect 11237 5810 11303 5813
rect 16297 5810 16363 5813
rect 11237 5808 16363 5810
rect 11237 5752 11242 5808
rect 11298 5752 16302 5808
rect 16358 5752 16363 5808
rect 11237 5750 16363 5752
rect 11237 5747 11303 5750
rect 16297 5747 16363 5750
rect 21725 5810 21791 5813
rect 22829 5810 22895 5813
rect 21725 5808 22895 5810
rect 21725 5752 21730 5808
rect 21786 5752 22834 5808
rect 22890 5752 22895 5808
rect 21725 5750 22895 5752
rect 21725 5747 21791 5750
rect 22829 5747 22895 5750
rect 23197 5810 23263 5813
rect 23800 5810 24600 5840
rect 23197 5808 24600 5810
rect 23197 5752 23202 5808
rect 23258 5752 24600 5808
rect 23197 5750 24600 5752
rect 23197 5747 23263 5750
rect 23800 5720 24600 5750
rect 19701 5674 19767 5677
rect 22553 5674 22619 5677
rect 19701 5672 22619 5674
rect 19701 5616 19706 5672
rect 19762 5616 22558 5672
rect 22614 5616 22619 5672
rect 19701 5614 22619 5616
rect 19701 5611 19767 5614
rect 22553 5611 22619 5614
rect 20069 5538 20135 5541
rect 22461 5538 22527 5541
rect 23105 5538 23171 5541
rect 20069 5536 23171 5538
rect 20069 5480 20074 5536
rect 20130 5480 22466 5536
rect 22522 5480 23110 5536
rect 23166 5480 23171 5536
rect 20069 5478 23171 5480
rect 20069 5475 20135 5478
rect 22461 5475 22527 5478
rect 23105 5475 23171 5478
rect 6544 5472 6860 5473
rect 6544 5408 6550 5472
rect 6614 5408 6630 5472
rect 6694 5408 6710 5472
rect 6774 5408 6790 5472
rect 6854 5408 6860 5472
rect 6544 5407 6860 5408
rect 12142 5472 12458 5473
rect 12142 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12458 5472
rect 12142 5407 12458 5408
rect 17740 5472 18056 5473
rect 17740 5408 17746 5472
rect 17810 5408 17826 5472
rect 17890 5408 17906 5472
rect 17970 5408 17986 5472
rect 18050 5408 18056 5472
rect 17740 5407 18056 5408
rect 19333 5402 19399 5405
rect 20529 5402 20595 5405
rect 19333 5400 20595 5402
rect 19333 5344 19338 5400
rect 19394 5344 20534 5400
rect 20590 5344 20595 5400
rect 19333 5342 20595 5344
rect 19333 5339 19399 5342
rect 20529 5339 20595 5342
rect 21173 5402 21239 5405
rect 22645 5402 22711 5405
rect 21173 5400 22711 5402
rect 21173 5344 21178 5400
rect 21234 5344 22650 5400
rect 22706 5344 22711 5400
rect 21173 5342 22711 5344
rect 21173 5339 21239 5342
rect 22645 5339 22711 5342
rect 20069 5266 20135 5269
rect 22645 5266 22711 5269
rect 20069 5264 22711 5266
rect 20069 5208 20074 5264
rect 20130 5208 22650 5264
rect 22706 5208 22711 5264
rect 20069 5206 22711 5208
rect 20069 5203 20135 5206
rect 22645 5203 22711 5206
rect 22921 5266 22987 5269
rect 23800 5266 24600 5296
rect 22921 5264 24600 5266
rect 22921 5208 22926 5264
rect 22982 5208 24600 5264
rect 22921 5206 24600 5208
rect 22921 5203 22987 5206
rect 23800 5176 24600 5206
rect 18822 5068 18828 5132
rect 18892 5130 18898 5132
rect 21173 5130 21239 5133
rect 18892 5128 21239 5130
rect 18892 5072 21178 5128
rect 21234 5072 21239 5128
rect 18892 5070 21239 5072
rect 18892 5068 18898 5070
rect 21173 5067 21239 5070
rect 3745 4928 4061 4929
rect 3745 4864 3751 4928
rect 3815 4864 3831 4928
rect 3895 4864 3911 4928
rect 3975 4864 3991 4928
rect 4055 4864 4061 4928
rect 3745 4863 4061 4864
rect 9343 4928 9659 4929
rect 9343 4864 9349 4928
rect 9413 4864 9429 4928
rect 9493 4864 9509 4928
rect 9573 4864 9589 4928
rect 9653 4864 9659 4928
rect 9343 4863 9659 4864
rect 14941 4928 15257 4929
rect 14941 4864 14947 4928
rect 15011 4864 15027 4928
rect 15091 4864 15107 4928
rect 15171 4864 15187 4928
rect 15251 4864 15257 4928
rect 14941 4863 15257 4864
rect 20539 4928 20855 4929
rect 20539 4864 20545 4928
rect 20609 4864 20625 4928
rect 20689 4864 20705 4928
rect 20769 4864 20785 4928
rect 20849 4864 20855 4928
rect 20539 4863 20855 4864
rect 19190 4660 19196 4724
rect 19260 4722 19266 4724
rect 20805 4722 20871 4725
rect 19260 4720 20871 4722
rect 19260 4664 20810 4720
rect 20866 4664 20871 4720
rect 19260 4662 20871 4664
rect 19260 4660 19266 4662
rect 20805 4659 20871 4662
rect 23013 4722 23079 4725
rect 23800 4722 24600 4752
rect 23013 4720 24600 4722
rect 23013 4664 23018 4720
rect 23074 4664 24600 4720
rect 23013 4662 24600 4664
rect 23013 4659 23079 4662
rect 23800 4632 24600 4662
rect 19006 4524 19012 4588
rect 19076 4586 19082 4588
rect 20253 4586 20319 4589
rect 19076 4584 20319 4586
rect 19076 4528 20258 4584
rect 20314 4528 20319 4584
rect 19076 4526 20319 4528
rect 19076 4524 19082 4526
rect 20253 4523 20319 4526
rect 6544 4384 6860 4385
rect 6544 4320 6550 4384
rect 6614 4320 6630 4384
rect 6694 4320 6710 4384
rect 6774 4320 6790 4384
rect 6854 4320 6860 4384
rect 6544 4319 6860 4320
rect 12142 4384 12458 4385
rect 12142 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12458 4384
rect 12142 4319 12458 4320
rect 17740 4384 18056 4385
rect 17740 4320 17746 4384
rect 17810 4320 17826 4384
rect 17890 4320 17906 4384
rect 17970 4320 17986 4384
rect 18050 4320 18056 4384
rect 17740 4319 18056 4320
rect 17166 4116 17172 4180
rect 17236 4178 17242 4180
rect 19241 4178 19307 4181
rect 22553 4178 22619 4181
rect 17236 4176 22619 4178
rect 17236 4120 19246 4176
rect 19302 4120 22558 4176
rect 22614 4120 22619 4176
rect 17236 4118 22619 4120
rect 17236 4116 17242 4118
rect 19241 4115 19307 4118
rect 21222 4045 21282 4118
rect 22553 4115 22619 4118
rect 23105 4178 23171 4181
rect 23800 4178 24600 4208
rect 23105 4176 24600 4178
rect 23105 4120 23110 4176
rect 23166 4120 24600 4176
rect 23105 4118 24600 4120
rect 23105 4115 23171 4118
rect 23800 4088 24600 4118
rect 16665 4044 16731 4045
rect 16614 3980 16620 4044
rect 16684 4042 16731 4044
rect 16684 4040 16776 4042
rect 16726 3984 16776 4040
rect 16684 3982 16776 3984
rect 21222 4040 21331 4045
rect 21222 3984 21270 4040
rect 21326 3984 21331 4040
rect 21222 3982 21331 3984
rect 16684 3980 16731 3982
rect 16665 3979 16731 3980
rect 21265 3979 21331 3982
rect 3745 3840 4061 3841
rect 3745 3776 3751 3840
rect 3815 3776 3831 3840
rect 3895 3776 3911 3840
rect 3975 3776 3991 3840
rect 4055 3776 4061 3840
rect 3745 3775 4061 3776
rect 9343 3840 9659 3841
rect 9343 3776 9349 3840
rect 9413 3776 9429 3840
rect 9493 3776 9509 3840
rect 9573 3776 9589 3840
rect 9653 3776 9659 3840
rect 9343 3775 9659 3776
rect 14941 3840 15257 3841
rect 14941 3776 14947 3840
rect 15011 3776 15027 3840
rect 15091 3776 15107 3840
rect 15171 3776 15187 3840
rect 15251 3776 15257 3840
rect 14941 3775 15257 3776
rect 20539 3840 20855 3841
rect 20539 3776 20545 3840
rect 20609 3776 20625 3840
rect 20689 3776 20705 3840
rect 20769 3776 20785 3840
rect 20849 3776 20855 3840
rect 20539 3775 20855 3776
rect 21030 3708 21036 3772
rect 21100 3770 21106 3772
rect 22737 3770 22803 3773
rect 21100 3768 22803 3770
rect 21100 3712 22742 3768
rect 22798 3712 22803 3768
rect 21100 3710 22803 3712
rect 21100 3708 21106 3710
rect 19517 3634 19583 3637
rect 21038 3634 21098 3708
rect 22737 3707 22803 3710
rect 19517 3632 21098 3634
rect 19517 3576 19522 3632
rect 19578 3576 21098 3632
rect 19517 3574 21098 3576
rect 21541 3634 21607 3637
rect 23800 3634 24600 3664
rect 21541 3632 24600 3634
rect 21541 3576 21546 3632
rect 21602 3576 24600 3632
rect 21541 3574 24600 3576
rect 19517 3571 19583 3574
rect 21541 3571 21607 3574
rect 23800 3544 24600 3574
rect 18505 3362 18571 3365
rect 22461 3362 22527 3365
rect 18505 3360 22527 3362
rect 18505 3304 18510 3360
rect 18566 3304 22466 3360
rect 22522 3304 22527 3360
rect 18505 3302 22527 3304
rect 18505 3299 18571 3302
rect 22461 3299 22527 3302
rect 6544 3296 6860 3297
rect 6544 3232 6550 3296
rect 6614 3232 6630 3296
rect 6694 3232 6710 3296
rect 6774 3232 6790 3296
rect 6854 3232 6860 3296
rect 6544 3231 6860 3232
rect 12142 3296 12458 3297
rect 12142 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12458 3296
rect 12142 3231 12458 3232
rect 17740 3296 18056 3297
rect 17740 3232 17746 3296
rect 17810 3232 17826 3296
rect 17890 3232 17906 3296
rect 17970 3232 17986 3296
rect 18050 3232 18056 3296
rect 17740 3231 18056 3232
rect 0 3090 800 3120
rect 1393 3090 1459 3093
rect 0 3088 1459 3090
rect 0 3032 1398 3088
rect 1454 3032 1459 3088
rect 0 3030 1459 3032
rect 0 3000 800 3030
rect 1393 3027 1459 3030
rect 23013 3090 23079 3093
rect 23800 3090 24600 3120
rect 23013 3088 24600 3090
rect 23013 3032 23018 3088
rect 23074 3032 24600 3088
rect 23013 3030 24600 3032
rect 23013 3027 23079 3030
rect 23800 3000 24600 3030
rect 19517 2954 19583 2957
rect 21725 2954 21791 2957
rect 19517 2952 21791 2954
rect 19517 2896 19522 2952
rect 19578 2896 21730 2952
rect 21786 2896 21791 2952
rect 19517 2894 21791 2896
rect 19517 2891 19583 2894
rect 21725 2891 21791 2894
rect 3745 2752 4061 2753
rect 3745 2688 3751 2752
rect 3815 2688 3831 2752
rect 3895 2688 3911 2752
rect 3975 2688 3991 2752
rect 4055 2688 4061 2752
rect 3745 2687 4061 2688
rect 9343 2752 9659 2753
rect 9343 2688 9349 2752
rect 9413 2688 9429 2752
rect 9493 2688 9509 2752
rect 9573 2688 9589 2752
rect 9653 2688 9659 2752
rect 9343 2687 9659 2688
rect 14941 2752 15257 2753
rect 14941 2688 14947 2752
rect 15011 2688 15027 2752
rect 15091 2688 15107 2752
rect 15171 2688 15187 2752
rect 15251 2688 15257 2752
rect 14941 2687 15257 2688
rect 20539 2752 20855 2753
rect 20539 2688 20545 2752
rect 20609 2688 20625 2752
rect 20689 2688 20705 2752
rect 20769 2688 20785 2752
rect 20849 2688 20855 2752
rect 20539 2687 20855 2688
rect 22645 2546 22711 2549
rect 23800 2546 24600 2576
rect 22645 2544 24600 2546
rect 22645 2488 22650 2544
rect 22706 2488 24600 2544
rect 22645 2486 24600 2488
rect 22645 2483 22711 2486
rect 23800 2456 24600 2486
rect 6544 2208 6860 2209
rect 6544 2144 6550 2208
rect 6614 2144 6630 2208
rect 6694 2144 6710 2208
rect 6774 2144 6790 2208
rect 6854 2144 6860 2208
rect 6544 2143 6860 2144
rect 12142 2208 12458 2209
rect 12142 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12458 2208
rect 12142 2143 12458 2144
rect 17740 2208 18056 2209
rect 17740 2144 17746 2208
rect 17810 2144 17826 2208
rect 17890 2144 17906 2208
rect 17970 2144 17986 2208
rect 18050 2144 18056 2208
rect 17740 2143 18056 2144
<< via3 >>
rect 3751 22332 3815 22336
rect 3751 22276 3755 22332
rect 3755 22276 3811 22332
rect 3811 22276 3815 22332
rect 3751 22272 3815 22276
rect 3831 22332 3895 22336
rect 3831 22276 3835 22332
rect 3835 22276 3891 22332
rect 3891 22276 3895 22332
rect 3831 22272 3895 22276
rect 3911 22332 3975 22336
rect 3911 22276 3915 22332
rect 3915 22276 3971 22332
rect 3971 22276 3975 22332
rect 3911 22272 3975 22276
rect 3991 22332 4055 22336
rect 3991 22276 3995 22332
rect 3995 22276 4051 22332
rect 4051 22276 4055 22332
rect 3991 22272 4055 22276
rect 9349 22332 9413 22336
rect 9349 22276 9353 22332
rect 9353 22276 9409 22332
rect 9409 22276 9413 22332
rect 9349 22272 9413 22276
rect 9429 22332 9493 22336
rect 9429 22276 9433 22332
rect 9433 22276 9489 22332
rect 9489 22276 9493 22332
rect 9429 22272 9493 22276
rect 9509 22332 9573 22336
rect 9509 22276 9513 22332
rect 9513 22276 9569 22332
rect 9569 22276 9573 22332
rect 9509 22272 9573 22276
rect 9589 22332 9653 22336
rect 9589 22276 9593 22332
rect 9593 22276 9649 22332
rect 9649 22276 9653 22332
rect 9589 22272 9653 22276
rect 14947 22332 15011 22336
rect 14947 22276 14951 22332
rect 14951 22276 15007 22332
rect 15007 22276 15011 22332
rect 14947 22272 15011 22276
rect 15027 22332 15091 22336
rect 15027 22276 15031 22332
rect 15031 22276 15087 22332
rect 15087 22276 15091 22332
rect 15027 22272 15091 22276
rect 15107 22332 15171 22336
rect 15107 22276 15111 22332
rect 15111 22276 15167 22332
rect 15167 22276 15171 22332
rect 15107 22272 15171 22276
rect 15187 22332 15251 22336
rect 15187 22276 15191 22332
rect 15191 22276 15247 22332
rect 15247 22276 15251 22332
rect 15187 22272 15251 22276
rect 20545 22332 20609 22336
rect 20545 22276 20549 22332
rect 20549 22276 20605 22332
rect 20605 22276 20609 22332
rect 20545 22272 20609 22276
rect 20625 22332 20689 22336
rect 20625 22276 20629 22332
rect 20629 22276 20685 22332
rect 20685 22276 20689 22332
rect 20625 22272 20689 22276
rect 20705 22332 20769 22336
rect 20705 22276 20709 22332
rect 20709 22276 20765 22332
rect 20765 22276 20769 22332
rect 20705 22272 20769 22276
rect 20785 22332 20849 22336
rect 20785 22276 20789 22332
rect 20789 22276 20845 22332
rect 20845 22276 20849 22332
rect 20785 22272 20849 22276
rect 5580 21932 5644 21996
rect 13308 21856 13372 21860
rect 13308 21800 13322 21856
rect 13322 21800 13372 21856
rect 13308 21796 13372 21800
rect 18276 21856 18340 21860
rect 18276 21800 18290 21856
rect 18290 21800 18340 21856
rect 18276 21796 18340 21800
rect 6550 21788 6614 21792
rect 6550 21732 6554 21788
rect 6554 21732 6610 21788
rect 6610 21732 6614 21788
rect 6550 21728 6614 21732
rect 6630 21788 6694 21792
rect 6630 21732 6634 21788
rect 6634 21732 6690 21788
rect 6690 21732 6694 21788
rect 6630 21728 6694 21732
rect 6710 21788 6774 21792
rect 6710 21732 6714 21788
rect 6714 21732 6770 21788
rect 6770 21732 6774 21788
rect 6710 21728 6774 21732
rect 6790 21788 6854 21792
rect 6790 21732 6794 21788
rect 6794 21732 6850 21788
rect 6850 21732 6854 21788
rect 6790 21728 6854 21732
rect 12148 21788 12212 21792
rect 12148 21732 12152 21788
rect 12152 21732 12208 21788
rect 12208 21732 12212 21788
rect 12148 21728 12212 21732
rect 12228 21788 12292 21792
rect 12228 21732 12232 21788
rect 12232 21732 12288 21788
rect 12288 21732 12292 21788
rect 12228 21728 12292 21732
rect 12308 21788 12372 21792
rect 12308 21732 12312 21788
rect 12312 21732 12368 21788
rect 12368 21732 12372 21788
rect 12308 21728 12372 21732
rect 12388 21788 12452 21792
rect 12388 21732 12392 21788
rect 12392 21732 12448 21788
rect 12448 21732 12452 21788
rect 12388 21728 12452 21732
rect 17746 21788 17810 21792
rect 17746 21732 17750 21788
rect 17750 21732 17806 21788
rect 17806 21732 17810 21788
rect 17746 21728 17810 21732
rect 17826 21788 17890 21792
rect 17826 21732 17830 21788
rect 17830 21732 17886 21788
rect 17886 21732 17890 21788
rect 17826 21728 17890 21732
rect 17906 21788 17970 21792
rect 17906 21732 17910 21788
rect 17910 21732 17966 21788
rect 17966 21732 17970 21788
rect 17906 21728 17970 21732
rect 17986 21788 18050 21792
rect 17986 21732 17990 21788
rect 17990 21732 18046 21788
rect 18046 21732 18050 21788
rect 17986 21728 18050 21732
rect 15332 21660 15396 21724
rect 3751 21244 3815 21248
rect 3751 21188 3755 21244
rect 3755 21188 3811 21244
rect 3811 21188 3815 21244
rect 3751 21184 3815 21188
rect 3831 21244 3895 21248
rect 3831 21188 3835 21244
rect 3835 21188 3891 21244
rect 3891 21188 3895 21244
rect 3831 21184 3895 21188
rect 3911 21244 3975 21248
rect 3911 21188 3915 21244
rect 3915 21188 3971 21244
rect 3971 21188 3975 21244
rect 3911 21184 3975 21188
rect 3991 21244 4055 21248
rect 3991 21188 3995 21244
rect 3995 21188 4051 21244
rect 4051 21188 4055 21244
rect 3991 21184 4055 21188
rect 9349 21244 9413 21248
rect 9349 21188 9353 21244
rect 9353 21188 9409 21244
rect 9409 21188 9413 21244
rect 9349 21184 9413 21188
rect 9429 21244 9493 21248
rect 9429 21188 9433 21244
rect 9433 21188 9489 21244
rect 9489 21188 9493 21244
rect 9429 21184 9493 21188
rect 9509 21244 9573 21248
rect 9509 21188 9513 21244
rect 9513 21188 9569 21244
rect 9569 21188 9573 21244
rect 9509 21184 9573 21188
rect 9589 21244 9653 21248
rect 9589 21188 9593 21244
rect 9593 21188 9649 21244
rect 9649 21188 9653 21244
rect 9589 21184 9653 21188
rect 14947 21244 15011 21248
rect 14947 21188 14951 21244
rect 14951 21188 15007 21244
rect 15007 21188 15011 21244
rect 14947 21184 15011 21188
rect 15027 21244 15091 21248
rect 15027 21188 15031 21244
rect 15031 21188 15087 21244
rect 15087 21188 15091 21244
rect 15027 21184 15091 21188
rect 15107 21244 15171 21248
rect 15107 21188 15111 21244
rect 15111 21188 15167 21244
rect 15167 21188 15171 21244
rect 15107 21184 15171 21188
rect 15187 21244 15251 21248
rect 15187 21188 15191 21244
rect 15191 21188 15247 21244
rect 15247 21188 15251 21244
rect 15187 21184 15251 21188
rect 12572 20980 12636 21044
rect 20545 21244 20609 21248
rect 20545 21188 20549 21244
rect 20549 21188 20605 21244
rect 20605 21188 20609 21244
rect 20545 21184 20609 21188
rect 20625 21244 20689 21248
rect 20625 21188 20629 21244
rect 20629 21188 20685 21244
rect 20685 21188 20689 21244
rect 20625 21184 20689 21188
rect 20705 21244 20769 21248
rect 20705 21188 20709 21244
rect 20709 21188 20765 21244
rect 20765 21188 20769 21244
rect 20705 21184 20769 21188
rect 20785 21244 20849 21248
rect 20785 21188 20789 21244
rect 20789 21188 20845 21244
rect 20845 21188 20849 21244
rect 20785 21184 20849 21188
rect 4844 20844 4908 20908
rect 6316 20844 6380 20908
rect 6550 20700 6614 20704
rect 6550 20644 6554 20700
rect 6554 20644 6610 20700
rect 6610 20644 6614 20700
rect 6550 20640 6614 20644
rect 6630 20700 6694 20704
rect 6630 20644 6634 20700
rect 6634 20644 6690 20700
rect 6690 20644 6694 20700
rect 6630 20640 6694 20644
rect 6710 20700 6774 20704
rect 6710 20644 6714 20700
rect 6714 20644 6770 20700
rect 6770 20644 6774 20700
rect 6710 20640 6774 20644
rect 6790 20700 6854 20704
rect 6790 20644 6794 20700
rect 6794 20644 6850 20700
rect 6850 20644 6854 20700
rect 6790 20640 6854 20644
rect 12148 20700 12212 20704
rect 12148 20644 12152 20700
rect 12152 20644 12208 20700
rect 12208 20644 12212 20700
rect 12148 20640 12212 20644
rect 12228 20700 12292 20704
rect 12228 20644 12232 20700
rect 12232 20644 12288 20700
rect 12288 20644 12292 20700
rect 12228 20640 12292 20644
rect 12308 20700 12372 20704
rect 12308 20644 12312 20700
rect 12312 20644 12368 20700
rect 12368 20644 12372 20700
rect 12308 20640 12372 20644
rect 12388 20700 12452 20704
rect 12388 20644 12392 20700
rect 12392 20644 12448 20700
rect 12448 20644 12452 20700
rect 12388 20640 12452 20644
rect 17746 20700 17810 20704
rect 17746 20644 17750 20700
rect 17750 20644 17806 20700
rect 17806 20644 17810 20700
rect 17746 20640 17810 20644
rect 17826 20700 17890 20704
rect 17826 20644 17830 20700
rect 17830 20644 17886 20700
rect 17886 20644 17890 20700
rect 17826 20640 17890 20644
rect 17906 20700 17970 20704
rect 17906 20644 17910 20700
rect 17910 20644 17966 20700
rect 17966 20644 17970 20700
rect 17906 20640 17970 20644
rect 17986 20700 18050 20704
rect 17986 20644 17990 20700
rect 17990 20644 18046 20700
rect 18046 20644 18050 20700
rect 17986 20640 18050 20644
rect 16988 20496 17052 20500
rect 16988 20440 17002 20496
rect 17002 20440 17052 20496
rect 16988 20436 17052 20440
rect 3751 20156 3815 20160
rect 3751 20100 3755 20156
rect 3755 20100 3811 20156
rect 3811 20100 3815 20156
rect 3751 20096 3815 20100
rect 3831 20156 3895 20160
rect 3831 20100 3835 20156
rect 3835 20100 3891 20156
rect 3891 20100 3895 20156
rect 3831 20096 3895 20100
rect 3911 20156 3975 20160
rect 3911 20100 3915 20156
rect 3915 20100 3971 20156
rect 3971 20100 3975 20156
rect 3911 20096 3975 20100
rect 3991 20156 4055 20160
rect 3991 20100 3995 20156
rect 3995 20100 4051 20156
rect 4051 20100 4055 20156
rect 3991 20096 4055 20100
rect 9349 20156 9413 20160
rect 9349 20100 9353 20156
rect 9353 20100 9409 20156
rect 9409 20100 9413 20156
rect 9349 20096 9413 20100
rect 9429 20156 9493 20160
rect 9429 20100 9433 20156
rect 9433 20100 9489 20156
rect 9489 20100 9493 20156
rect 9429 20096 9493 20100
rect 9509 20156 9573 20160
rect 9509 20100 9513 20156
rect 9513 20100 9569 20156
rect 9569 20100 9573 20156
rect 9509 20096 9573 20100
rect 9589 20156 9653 20160
rect 9589 20100 9593 20156
rect 9593 20100 9649 20156
rect 9649 20100 9653 20156
rect 9589 20096 9653 20100
rect 14947 20156 15011 20160
rect 14947 20100 14951 20156
rect 14951 20100 15007 20156
rect 15007 20100 15011 20156
rect 14947 20096 15011 20100
rect 15027 20156 15091 20160
rect 15027 20100 15031 20156
rect 15031 20100 15087 20156
rect 15087 20100 15091 20156
rect 15027 20096 15091 20100
rect 15107 20156 15171 20160
rect 15107 20100 15111 20156
rect 15111 20100 15167 20156
rect 15167 20100 15171 20156
rect 15107 20096 15171 20100
rect 15187 20156 15251 20160
rect 15187 20100 15191 20156
rect 15191 20100 15247 20156
rect 15247 20100 15251 20156
rect 15187 20096 15251 20100
rect 20545 20156 20609 20160
rect 20545 20100 20549 20156
rect 20549 20100 20605 20156
rect 20605 20100 20609 20156
rect 20545 20096 20609 20100
rect 20625 20156 20689 20160
rect 20625 20100 20629 20156
rect 20629 20100 20685 20156
rect 20685 20100 20689 20156
rect 20625 20096 20689 20100
rect 20705 20156 20769 20160
rect 20705 20100 20709 20156
rect 20709 20100 20765 20156
rect 20765 20100 20769 20156
rect 20705 20096 20769 20100
rect 20785 20156 20849 20160
rect 20785 20100 20789 20156
rect 20789 20100 20845 20156
rect 20845 20100 20849 20156
rect 20785 20096 20849 20100
rect 16436 20028 16500 20092
rect 6550 19612 6614 19616
rect 6550 19556 6554 19612
rect 6554 19556 6610 19612
rect 6610 19556 6614 19612
rect 6550 19552 6614 19556
rect 6630 19612 6694 19616
rect 6630 19556 6634 19612
rect 6634 19556 6690 19612
rect 6690 19556 6694 19612
rect 6630 19552 6694 19556
rect 6710 19612 6774 19616
rect 6710 19556 6714 19612
rect 6714 19556 6770 19612
rect 6770 19556 6774 19612
rect 6710 19552 6774 19556
rect 6790 19612 6854 19616
rect 6790 19556 6794 19612
rect 6794 19556 6850 19612
rect 6850 19556 6854 19612
rect 6790 19552 6854 19556
rect 12148 19612 12212 19616
rect 12148 19556 12152 19612
rect 12152 19556 12208 19612
rect 12208 19556 12212 19612
rect 12148 19552 12212 19556
rect 12228 19612 12292 19616
rect 12228 19556 12232 19612
rect 12232 19556 12288 19612
rect 12288 19556 12292 19612
rect 12228 19552 12292 19556
rect 12308 19612 12372 19616
rect 12308 19556 12312 19612
rect 12312 19556 12368 19612
rect 12368 19556 12372 19612
rect 12308 19552 12372 19556
rect 12388 19612 12452 19616
rect 12388 19556 12392 19612
rect 12392 19556 12448 19612
rect 12448 19556 12452 19612
rect 12388 19552 12452 19556
rect 17746 19612 17810 19616
rect 17746 19556 17750 19612
rect 17750 19556 17806 19612
rect 17806 19556 17810 19612
rect 17746 19552 17810 19556
rect 17826 19612 17890 19616
rect 17826 19556 17830 19612
rect 17830 19556 17886 19612
rect 17886 19556 17890 19612
rect 17826 19552 17890 19556
rect 17906 19612 17970 19616
rect 17906 19556 17910 19612
rect 17910 19556 17966 19612
rect 17966 19556 17970 19612
rect 17906 19552 17970 19556
rect 17986 19612 18050 19616
rect 17986 19556 17990 19612
rect 17990 19556 18046 19612
rect 18046 19556 18050 19612
rect 17986 19552 18050 19556
rect 16436 19544 16500 19548
rect 16436 19488 16486 19544
rect 16486 19488 16500 19544
rect 16436 19484 16500 19488
rect 18460 19484 18524 19548
rect 16620 19408 16684 19412
rect 16620 19352 16634 19408
rect 16634 19352 16684 19408
rect 16620 19348 16684 19352
rect 16988 19348 17052 19412
rect 3751 19068 3815 19072
rect 3751 19012 3755 19068
rect 3755 19012 3811 19068
rect 3811 19012 3815 19068
rect 3751 19008 3815 19012
rect 3831 19068 3895 19072
rect 3831 19012 3835 19068
rect 3835 19012 3891 19068
rect 3891 19012 3895 19068
rect 3831 19008 3895 19012
rect 3911 19068 3975 19072
rect 3911 19012 3915 19068
rect 3915 19012 3971 19068
rect 3971 19012 3975 19068
rect 3911 19008 3975 19012
rect 3991 19068 4055 19072
rect 3991 19012 3995 19068
rect 3995 19012 4051 19068
rect 4051 19012 4055 19068
rect 3991 19008 4055 19012
rect 9349 19068 9413 19072
rect 9349 19012 9353 19068
rect 9353 19012 9409 19068
rect 9409 19012 9413 19068
rect 9349 19008 9413 19012
rect 9429 19068 9493 19072
rect 9429 19012 9433 19068
rect 9433 19012 9489 19068
rect 9489 19012 9493 19068
rect 9429 19008 9493 19012
rect 9509 19068 9573 19072
rect 9509 19012 9513 19068
rect 9513 19012 9569 19068
rect 9569 19012 9573 19068
rect 9509 19008 9573 19012
rect 9589 19068 9653 19072
rect 9589 19012 9593 19068
rect 9593 19012 9649 19068
rect 9649 19012 9653 19068
rect 9589 19008 9653 19012
rect 14947 19068 15011 19072
rect 14947 19012 14951 19068
rect 14951 19012 15007 19068
rect 15007 19012 15011 19068
rect 14947 19008 15011 19012
rect 15027 19068 15091 19072
rect 15027 19012 15031 19068
rect 15031 19012 15087 19068
rect 15087 19012 15091 19068
rect 15027 19008 15091 19012
rect 15107 19068 15171 19072
rect 15107 19012 15111 19068
rect 15111 19012 15167 19068
rect 15167 19012 15171 19068
rect 15107 19008 15171 19012
rect 15187 19068 15251 19072
rect 15187 19012 15191 19068
rect 15191 19012 15247 19068
rect 15247 19012 15251 19068
rect 15187 19008 15251 19012
rect 20545 19068 20609 19072
rect 20545 19012 20549 19068
rect 20549 19012 20605 19068
rect 20605 19012 20609 19068
rect 20545 19008 20609 19012
rect 20625 19068 20689 19072
rect 20625 19012 20629 19068
rect 20629 19012 20685 19068
rect 20685 19012 20689 19068
rect 20625 19008 20689 19012
rect 20705 19068 20769 19072
rect 20705 19012 20709 19068
rect 20709 19012 20765 19068
rect 20765 19012 20769 19068
rect 20705 19008 20769 19012
rect 20785 19068 20849 19072
rect 20785 19012 20789 19068
rect 20789 19012 20845 19068
rect 20845 19012 20849 19068
rect 20785 19008 20849 19012
rect 13308 18804 13372 18868
rect 19932 18804 19996 18868
rect 6550 18524 6614 18528
rect 6550 18468 6554 18524
rect 6554 18468 6610 18524
rect 6610 18468 6614 18524
rect 6550 18464 6614 18468
rect 6630 18524 6694 18528
rect 6630 18468 6634 18524
rect 6634 18468 6690 18524
rect 6690 18468 6694 18524
rect 6630 18464 6694 18468
rect 6710 18524 6774 18528
rect 6710 18468 6714 18524
rect 6714 18468 6770 18524
rect 6770 18468 6774 18524
rect 6710 18464 6774 18468
rect 6790 18524 6854 18528
rect 6790 18468 6794 18524
rect 6794 18468 6850 18524
rect 6850 18468 6854 18524
rect 6790 18464 6854 18468
rect 12148 18524 12212 18528
rect 12148 18468 12152 18524
rect 12152 18468 12208 18524
rect 12208 18468 12212 18524
rect 12148 18464 12212 18468
rect 12228 18524 12292 18528
rect 12228 18468 12232 18524
rect 12232 18468 12288 18524
rect 12288 18468 12292 18524
rect 12228 18464 12292 18468
rect 12308 18524 12372 18528
rect 12308 18468 12312 18524
rect 12312 18468 12368 18524
rect 12368 18468 12372 18524
rect 12308 18464 12372 18468
rect 12388 18524 12452 18528
rect 12388 18468 12392 18524
rect 12392 18468 12448 18524
rect 12448 18468 12452 18524
rect 12388 18464 12452 18468
rect 17746 18524 17810 18528
rect 17746 18468 17750 18524
rect 17750 18468 17806 18524
rect 17806 18468 17810 18524
rect 17746 18464 17810 18468
rect 17826 18524 17890 18528
rect 17826 18468 17830 18524
rect 17830 18468 17886 18524
rect 17886 18468 17890 18524
rect 17826 18464 17890 18468
rect 17906 18524 17970 18528
rect 17906 18468 17910 18524
rect 17910 18468 17966 18524
rect 17966 18468 17970 18524
rect 17906 18464 17970 18468
rect 17986 18524 18050 18528
rect 17986 18468 17990 18524
rect 17990 18468 18046 18524
rect 18046 18468 18050 18524
rect 17986 18464 18050 18468
rect 3751 17980 3815 17984
rect 3751 17924 3755 17980
rect 3755 17924 3811 17980
rect 3811 17924 3815 17980
rect 3751 17920 3815 17924
rect 3831 17980 3895 17984
rect 3831 17924 3835 17980
rect 3835 17924 3891 17980
rect 3891 17924 3895 17980
rect 3831 17920 3895 17924
rect 3911 17980 3975 17984
rect 3911 17924 3915 17980
rect 3915 17924 3971 17980
rect 3971 17924 3975 17980
rect 3911 17920 3975 17924
rect 3991 17980 4055 17984
rect 3991 17924 3995 17980
rect 3995 17924 4051 17980
rect 4051 17924 4055 17980
rect 3991 17920 4055 17924
rect 9349 17980 9413 17984
rect 9349 17924 9353 17980
rect 9353 17924 9409 17980
rect 9409 17924 9413 17980
rect 9349 17920 9413 17924
rect 9429 17980 9493 17984
rect 9429 17924 9433 17980
rect 9433 17924 9489 17980
rect 9489 17924 9493 17980
rect 9429 17920 9493 17924
rect 9509 17980 9573 17984
rect 9509 17924 9513 17980
rect 9513 17924 9569 17980
rect 9569 17924 9573 17980
rect 9509 17920 9573 17924
rect 9589 17980 9653 17984
rect 9589 17924 9593 17980
rect 9593 17924 9649 17980
rect 9649 17924 9653 17980
rect 9589 17920 9653 17924
rect 14947 17980 15011 17984
rect 14947 17924 14951 17980
rect 14951 17924 15007 17980
rect 15007 17924 15011 17980
rect 14947 17920 15011 17924
rect 15027 17980 15091 17984
rect 15027 17924 15031 17980
rect 15031 17924 15087 17980
rect 15087 17924 15091 17980
rect 15027 17920 15091 17924
rect 15107 17980 15171 17984
rect 15107 17924 15111 17980
rect 15111 17924 15167 17980
rect 15167 17924 15171 17980
rect 15107 17920 15171 17924
rect 15187 17980 15251 17984
rect 15187 17924 15191 17980
rect 15191 17924 15247 17980
rect 15247 17924 15251 17980
rect 15187 17920 15251 17924
rect 20545 17980 20609 17984
rect 20545 17924 20549 17980
rect 20549 17924 20605 17980
rect 20605 17924 20609 17980
rect 20545 17920 20609 17924
rect 20625 17980 20689 17984
rect 20625 17924 20629 17980
rect 20629 17924 20685 17980
rect 20685 17924 20689 17980
rect 20625 17920 20689 17924
rect 20705 17980 20769 17984
rect 20705 17924 20709 17980
rect 20709 17924 20765 17980
rect 20765 17924 20769 17980
rect 20705 17920 20769 17924
rect 20785 17980 20849 17984
rect 20785 17924 20789 17980
rect 20789 17924 20845 17980
rect 20845 17924 20849 17980
rect 20785 17920 20849 17924
rect 15332 17580 15396 17644
rect 6550 17436 6614 17440
rect 6550 17380 6554 17436
rect 6554 17380 6610 17436
rect 6610 17380 6614 17436
rect 6550 17376 6614 17380
rect 6630 17436 6694 17440
rect 6630 17380 6634 17436
rect 6634 17380 6690 17436
rect 6690 17380 6694 17436
rect 6630 17376 6694 17380
rect 6710 17436 6774 17440
rect 6710 17380 6714 17436
rect 6714 17380 6770 17436
rect 6770 17380 6774 17436
rect 6710 17376 6774 17380
rect 6790 17436 6854 17440
rect 6790 17380 6794 17436
rect 6794 17380 6850 17436
rect 6850 17380 6854 17436
rect 6790 17376 6854 17380
rect 12148 17436 12212 17440
rect 12148 17380 12152 17436
rect 12152 17380 12208 17436
rect 12208 17380 12212 17436
rect 12148 17376 12212 17380
rect 12228 17436 12292 17440
rect 12228 17380 12232 17436
rect 12232 17380 12288 17436
rect 12288 17380 12292 17436
rect 12228 17376 12292 17380
rect 12308 17436 12372 17440
rect 12308 17380 12312 17436
rect 12312 17380 12368 17436
rect 12368 17380 12372 17436
rect 12308 17376 12372 17380
rect 12388 17436 12452 17440
rect 12388 17380 12392 17436
rect 12392 17380 12448 17436
rect 12448 17380 12452 17436
rect 12388 17376 12452 17380
rect 17746 17436 17810 17440
rect 17746 17380 17750 17436
rect 17750 17380 17806 17436
rect 17806 17380 17810 17436
rect 17746 17376 17810 17380
rect 17826 17436 17890 17440
rect 17826 17380 17830 17436
rect 17830 17380 17886 17436
rect 17886 17380 17890 17436
rect 17826 17376 17890 17380
rect 17906 17436 17970 17440
rect 17906 17380 17910 17436
rect 17910 17380 17966 17436
rect 17966 17380 17970 17436
rect 17906 17376 17970 17380
rect 17986 17436 18050 17440
rect 17986 17380 17990 17436
rect 17990 17380 18046 17436
rect 18046 17380 18050 17436
rect 17986 17376 18050 17380
rect 3751 16892 3815 16896
rect 3751 16836 3755 16892
rect 3755 16836 3811 16892
rect 3811 16836 3815 16892
rect 3751 16832 3815 16836
rect 3831 16892 3895 16896
rect 3831 16836 3835 16892
rect 3835 16836 3891 16892
rect 3891 16836 3895 16892
rect 3831 16832 3895 16836
rect 3911 16892 3975 16896
rect 3911 16836 3915 16892
rect 3915 16836 3971 16892
rect 3971 16836 3975 16892
rect 3911 16832 3975 16836
rect 3991 16892 4055 16896
rect 3991 16836 3995 16892
rect 3995 16836 4051 16892
rect 4051 16836 4055 16892
rect 3991 16832 4055 16836
rect 9349 16892 9413 16896
rect 9349 16836 9353 16892
rect 9353 16836 9409 16892
rect 9409 16836 9413 16892
rect 9349 16832 9413 16836
rect 9429 16892 9493 16896
rect 9429 16836 9433 16892
rect 9433 16836 9489 16892
rect 9489 16836 9493 16892
rect 9429 16832 9493 16836
rect 9509 16892 9573 16896
rect 9509 16836 9513 16892
rect 9513 16836 9569 16892
rect 9569 16836 9573 16892
rect 9509 16832 9573 16836
rect 9589 16892 9653 16896
rect 9589 16836 9593 16892
rect 9593 16836 9649 16892
rect 9649 16836 9653 16892
rect 9589 16832 9653 16836
rect 14947 16892 15011 16896
rect 14947 16836 14951 16892
rect 14951 16836 15007 16892
rect 15007 16836 15011 16892
rect 14947 16832 15011 16836
rect 15027 16892 15091 16896
rect 15027 16836 15031 16892
rect 15031 16836 15087 16892
rect 15087 16836 15091 16892
rect 15027 16832 15091 16836
rect 15107 16892 15171 16896
rect 15107 16836 15111 16892
rect 15111 16836 15167 16892
rect 15167 16836 15171 16892
rect 15107 16832 15171 16836
rect 15187 16892 15251 16896
rect 15187 16836 15191 16892
rect 15191 16836 15247 16892
rect 15247 16836 15251 16892
rect 15187 16832 15251 16836
rect 20545 16892 20609 16896
rect 20545 16836 20549 16892
rect 20549 16836 20605 16892
rect 20605 16836 20609 16892
rect 20545 16832 20609 16836
rect 20625 16892 20689 16896
rect 20625 16836 20629 16892
rect 20629 16836 20685 16892
rect 20685 16836 20689 16892
rect 20625 16832 20689 16836
rect 20705 16892 20769 16896
rect 20705 16836 20709 16892
rect 20709 16836 20765 16892
rect 20765 16836 20769 16892
rect 20705 16832 20769 16836
rect 20785 16892 20849 16896
rect 20785 16836 20789 16892
rect 20789 16836 20845 16892
rect 20845 16836 20849 16892
rect 20785 16832 20849 16836
rect 12572 16492 12636 16556
rect 6550 16348 6614 16352
rect 6550 16292 6554 16348
rect 6554 16292 6610 16348
rect 6610 16292 6614 16348
rect 6550 16288 6614 16292
rect 6630 16348 6694 16352
rect 6630 16292 6634 16348
rect 6634 16292 6690 16348
rect 6690 16292 6694 16348
rect 6630 16288 6694 16292
rect 6710 16348 6774 16352
rect 6710 16292 6714 16348
rect 6714 16292 6770 16348
rect 6770 16292 6774 16348
rect 6710 16288 6774 16292
rect 6790 16348 6854 16352
rect 6790 16292 6794 16348
rect 6794 16292 6850 16348
rect 6850 16292 6854 16348
rect 6790 16288 6854 16292
rect 12148 16348 12212 16352
rect 12148 16292 12152 16348
rect 12152 16292 12208 16348
rect 12208 16292 12212 16348
rect 12148 16288 12212 16292
rect 12228 16348 12292 16352
rect 12228 16292 12232 16348
rect 12232 16292 12288 16348
rect 12288 16292 12292 16348
rect 12228 16288 12292 16292
rect 12308 16348 12372 16352
rect 12308 16292 12312 16348
rect 12312 16292 12368 16348
rect 12368 16292 12372 16348
rect 12308 16288 12372 16292
rect 12388 16348 12452 16352
rect 12388 16292 12392 16348
rect 12392 16292 12448 16348
rect 12448 16292 12452 16348
rect 12388 16288 12452 16292
rect 17746 16348 17810 16352
rect 17746 16292 17750 16348
rect 17750 16292 17806 16348
rect 17806 16292 17810 16348
rect 17746 16288 17810 16292
rect 17826 16348 17890 16352
rect 17826 16292 17830 16348
rect 17830 16292 17886 16348
rect 17886 16292 17890 16348
rect 17826 16288 17890 16292
rect 17906 16348 17970 16352
rect 17906 16292 17910 16348
rect 17910 16292 17966 16348
rect 17966 16292 17970 16348
rect 17906 16288 17970 16292
rect 17986 16348 18050 16352
rect 17986 16292 17990 16348
rect 17990 16292 18046 16348
rect 18046 16292 18050 16348
rect 17986 16288 18050 16292
rect 3751 15804 3815 15808
rect 3751 15748 3755 15804
rect 3755 15748 3811 15804
rect 3811 15748 3815 15804
rect 3751 15744 3815 15748
rect 3831 15804 3895 15808
rect 3831 15748 3835 15804
rect 3835 15748 3891 15804
rect 3891 15748 3895 15804
rect 3831 15744 3895 15748
rect 3911 15804 3975 15808
rect 3911 15748 3915 15804
rect 3915 15748 3971 15804
rect 3971 15748 3975 15804
rect 3911 15744 3975 15748
rect 3991 15804 4055 15808
rect 3991 15748 3995 15804
rect 3995 15748 4051 15804
rect 4051 15748 4055 15804
rect 3991 15744 4055 15748
rect 9349 15804 9413 15808
rect 9349 15748 9353 15804
rect 9353 15748 9409 15804
rect 9409 15748 9413 15804
rect 9349 15744 9413 15748
rect 9429 15804 9493 15808
rect 9429 15748 9433 15804
rect 9433 15748 9489 15804
rect 9489 15748 9493 15804
rect 9429 15744 9493 15748
rect 9509 15804 9573 15808
rect 9509 15748 9513 15804
rect 9513 15748 9569 15804
rect 9569 15748 9573 15804
rect 9509 15744 9573 15748
rect 9589 15804 9653 15808
rect 9589 15748 9593 15804
rect 9593 15748 9649 15804
rect 9649 15748 9653 15804
rect 9589 15744 9653 15748
rect 14947 15804 15011 15808
rect 14947 15748 14951 15804
rect 14951 15748 15007 15804
rect 15007 15748 15011 15804
rect 14947 15744 15011 15748
rect 15027 15804 15091 15808
rect 15027 15748 15031 15804
rect 15031 15748 15087 15804
rect 15087 15748 15091 15804
rect 15027 15744 15091 15748
rect 15107 15804 15171 15808
rect 15107 15748 15111 15804
rect 15111 15748 15167 15804
rect 15167 15748 15171 15804
rect 15107 15744 15171 15748
rect 15187 15804 15251 15808
rect 15187 15748 15191 15804
rect 15191 15748 15247 15804
rect 15247 15748 15251 15804
rect 15187 15744 15251 15748
rect 20545 15804 20609 15808
rect 20545 15748 20549 15804
rect 20549 15748 20605 15804
rect 20605 15748 20609 15804
rect 20545 15744 20609 15748
rect 20625 15804 20689 15808
rect 20625 15748 20629 15804
rect 20629 15748 20685 15804
rect 20685 15748 20689 15804
rect 20625 15744 20689 15748
rect 20705 15804 20769 15808
rect 20705 15748 20709 15804
rect 20709 15748 20765 15804
rect 20765 15748 20769 15804
rect 20705 15744 20769 15748
rect 20785 15804 20849 15808
rect 20785 15748 20789 15804
rect 20789 15748 20845 15804
rect 20845 15748 20849 15804
rect 20785 15744 20849 15748
rect 4292 15328 4356 15332
rect 4292 15272 4306 15328
rect 4306 15272 4356 15328
rect 4292 15268 4356 15272
rect 6550 15260 6614 15264
rect 6550 15204 6554 15260
rect 6554 15204 6610 15260
rect 6610 15204 6614 15260
rect 6550 15200 6614 15204
rect 6630 15260 6694 15264
rect 6630 15204 6634 15260
rect 6634 15204 6690 15260
rect 6690 15204 6694 15260
rect 6630 15200 6694 15204
rect 6710 15260 6774 15264
rect 6710 15204 6714 15260
rect 6714 15204 6770 15260
rect 6770 15204 6774 15260
rect 6710 15200 6774 15204
rect 6790 15260 6854 15264
rect 6790 15204 6794 15260
rect 6794 15204 6850 15260
rect 6850 15204 6854 15260
rect 6790 15200 6854 15204
rect 12148 15260 12212 15264
rect 12148 15204 12152 15260
rect 12152 15204 12208 15260
rect 12208 15204 12212 15260
rect 12148 15200 12212 15204
rect 12228 15260 12292 15264
rect 12228 15204 12232 15260
rect 12232 15204 12288 15260
rect 12288 15204 12292 15260
rect 12228 15200 12292 15204
rect 12308 15260 12372 15264
rect 12308 15204 12312 15260
rect 12312 15204 12368 15260
rect 12368 15204 12372 15260
rect 12308 15200 12372 15204
rect 12388 15260 12452 15264
rect 12388 15204 12392 15260
rect 12392 15204 12448 15260
rect 12448 15204 12452 15260
rect 12388 15200 12452 15204
rect 17746 15260 17810 15264
rect 17746 15204 17750 15260
rect 17750 15204 17806 15260
rect 17806 15204 17810 15260
rect 17746 15200 17810 15204
rect 17826 15260 17890 15264
rect 17826 15204 17830 15260
rect 17830 15204 17886 15260
rect 17886 15204 17890 15260
rect 17826 15200 17890 15204
rect 17906 15260 17970 15264
rect 17906 15204 17910 15260
rect 17910 15204 17966 15260
rect 17966 15204 17970 15260
rect 17906 15200 17970 15204
rect 17986 15260 18050 15264
rect 17986 15204 17990 15260
rect 17990 15204 18046 15260
rect 18046 15204 18050 15260
rect 17986 15200 18050 15204
rect 16620 15192 16684 15196
rect 16620 15136 16634 15192
rect 16634 15136 16684 15192
rect 16620 15132 16684 15136
rect 4844 15056 4908 15060
rect 4844 15000 4894 15056
rect 4894 15000 4908 15056
rect 4844 14996 4908 15000
rect 3751 14716 3815 14720
rect 3751 14660 3755 14716
rect 3755 14660 3811 14716
rect 3811 14660 3815 14716
rect 3751 14656 3815 14660
rect 3831 14716 3895 14720
rect 3831 14660 3835 14716
rect 3835 14660 3891 14716
rect 3891 14660 3895 14716
rect 3831 14656 3895 14660
rect 3911 14716 3975 14720
rect 3911 14660 3915 14716
rect 3915 14660 3971 14716
rect 3971 14660 3975 14716
rect 3911 14656 3975 14660
rect 3991 14716 4055 14720
rect 3991 14660 3995 14716
rect 3995 14660 4051 14716
rect 4051 14660 4055 14716
rect 3991 14656 4055 14660
rect 9349 14716 9413 14720
rect 9349 14660 9353 14716
rect 9353 14660 9409 14716
rect 9409 14660 9413 14716
rect 9349 14656 9413 14660
rect 9429 14716 9493 14720
rect 9429 14660 9433 14716
rect 9433 14660 9489 14716
rect 9489 14660 9493 14716
rect 9429 14656 9493 14660
rect 9509 14716 9573 14720
rect 9509 14660 9513 14716
rect 9513 14660 9569 14716
rect 9569 14660 9573 14716
rect 9509 14656 9573 14660
rect 9589 14716 9653 14720
rect 9589 14660 9593 14716
rect 9593 14660 9649 14716
rect 9649 14660 9653 14716
rect 9589 14656 9653 14660
rect 14947 14716 15011 14720
rect 14947 14660 14951 14716
rect 14951 14660 15007 14716
rect 15007 14660 15011 14716
rect 14947 14656 15011 14660
rect 15027 14716 15091 14720
rect 15027 14660 15031 14716
rect 15031 14660 15087 14716
rect 15087 14660 15091 14716
rect 15027 14656 15091 14660
rect 15107 14716 15171 14720
rect 15107 14660 15111 14716
rect 15111 14660 15167 14716
rect 15167 14660 15171 14716
rect 15107 14656 15171 14660
rect 15187 14716 15251 14720
rect 15187 14660 15191 14716
rect 15191 14660 15247 14716
rect 15247 14660 15251 14716
rect 15187 14656 15251 14660
rect 20545 14716 20609 14720
rect 20545 14660 20549 14716
rect 20549 14660 20605 14716
rect 20605 14660 20609 14716
rect 20545 14656 20609 14660
rect 20625 14716 20689 14720
rect 20625 14660 20629 14716
rect 20629 14660 20685 14716
rect 20685 14660 20689 14716
rect 20625 14656 20689 14660
rect 20705 14716 20769 14720
rect 20705 14660 20709 14716
rect 20709 14660 20765 14716
rect 20765 14660 20769 14716
rect 20705 14656 20769 14660
rect 20785 14716 20849 14720
rect 20785 14660 20789 14716
rect 20789 14660 20845 14716
rect 20845 14660 20849 14716
rect 20785 14656 20849 14660
rect 17172 14180 17236 14244
rect 6550 14172 6614 14176
rect 6550 14116 6554 14172
rect 6554 14116 6610 14172
rect 6610 14116 6614 14172
rect 6550 14112 6614 14116
rect 6630 14172 6694 14176
rect 6630 14116 6634 14172
rect 6634 14116 6690 14172
rect 6690 14116 6694 14172
rect 6630 14112 6694 14116
rect 6710 14172 6774 14176
rect 6710 14116 6714 14172
rect 6714 14116 6770 14172
rect 6770 14116 6774 14172
rect 6710 14112 6774 14116
rect 6790 14172 6854 14176
rect 6790 14116 6794 14172
rect 6794 14116 6850 14172
rect 6850 14116 6854 14172
rect 6790 14112 6854 14116
rect 12148 14172 12212 14176
rect 12148 14116 12152 14172
rect 12152 14116 12208 14172
rect 12208 14116 12212 14172
rect 12148 14112 12212 14116
rect 12228 14172 12292 14176
rect 12228 14116 12232 14172
rect 12232 14116 12288 14172
rect 12288 14116 12292 14172
rect 12228 14112 12292 14116
rect 12308 14172 12372 14176
rect 12308 14116 12312 14172
rect 12312 14116 12368 14172
rect 12368 14116 12372 14172
rect 12308 14112 12372 14116
rect 12388 14172 12452 14176
rect 12388 14116 12392 14172
rect 12392 14116 12448 14172
rect 12448 14116 12452 14172
rect 12388 14112 12452 14116
rect 17746 14172 17810 14176
rect 17746 14116 17750 14172
rect 17750 14116 17806 14172
rect 17806 14116 17810 14172
rect 17746 14112 17810 14116
rect 17826 14172 17890 14176
rect 17826 14116 17830 14172
rect 17830 14116 17886 14172
rect 17886 14116 17890 14172
rect 17826 14112 17890 14116
rect 17906 14172 17970 14176
rect 17906 14116 17910 14172
rect 17910 14116 17966 14172
rect 17966 14116 17970 14172
rect 17906 14112 17970 14116
rect 17986 14172 18050 14176
rect 17986 14116 17990 14172
rect 17990 14116 18046 14172
rect 18046 14116 18050 14172
rect 17986 14112 18050 14116
rect 3751 13628 3815 13632
rect 3751 13572 3755 13628
rect 3755 13572 3811 13628
rect 3811 13572 3815 13628
rect 3751 13568 3815 13572
rect 3831 13628 3895 13632
rect 3831 13572 3835 13628
rect 3835 13572 3891 13628
rect 3891 13572 3895 13628
rect 3831 13568 3895 13572
rect 3911 13628 3975 13632
rect 3911 13572 3915 13628
rect 3915 13572 3971 13628
rect 3971 13572 3975 13628
rect 3911 13568 3975 13572
rect 3991 13628 4055 13632
rect 3991 13572 3995 13628
rect 3995 13572 4051 13628
rect 4051 13572 4055 13628
rect 3991 13568 4055 13572
rect 9349 13628 9413 13632
rect 9349 13572 9353 13628
rect 9353 13572 9409 13628
rect 9409 13572 9413 13628
rect 9349 13568 9413 13572
rect 9429 13628 9493 13632
rect 9429 13572 9433 13628
rect 9433 13572 9489 13628
rect 9489 13572 9493 13628
rect 9429 13568 9493 13572
rect 9509 13628 9573 13632
rect 9509 13572 9513 13628
rect 9513 13572 9569 13628
rect 9569 13572 9573 13628
rect 9509 13568 9573 13572
rect 9589 13628 9653 13632
rect 9589 13572 9593 13628
rect 9593 13572 9649 13628
rect 9649 13572 9653 13628
rect 9589 13568 9653 13572
rect 14947 13628 15011 13632
rect 14947 13572 14951 13628
rect 14951 13572 15007 13628
rect 15007 13572 15011 13628
rect 14947 13568 15011 13572
rect 15027 13628 15091 13632
rect 15027 13572 15031 13628
rect 15031 13572 15087 13628
rect 15087 13572 15091 13628
rect 15027 13568 15091 13572
rect 15107 13628 15171 13632
rect 15107 13572 15111 13628
rect 15111 13572 15167 13628
rect 15167 13572 15171 13628
rect 15107 13568 15171 13572
rect 15187 13628 15251 13632
rect 15187 13572 15191 13628
rect 15191 13572 15247 13628
rect 15247 13572 15251 13628
rect 15187 13568 15251 13572
rect 20545 13628 20609 13632
rect 20545 13572 20549 13628
rect 20549 13572 20605 13628
rect 20605 13572 20609 13628
rect 20545 13568 20609 13572
rect 20625 13628 20689 13632
rect 20625 13572 20629 13628
rect 20629 13572 20685 13628
rect 20685 13572 20689 13628
rect 20625 13568 20689 13572
rect 20705 13628 20769 13632
rect 20705 13572 20709 13628
rect 20709 13572 20765 13628
rect 20765 13572 20769 13628
rect 20705 13568 20769 13572
rect 20785 13628 20849 13632
rect 20785 13572 20789 13628
rect 20789 13572 20845 13628
rect 20845 13572 20849 13628
rect 20785 13568 20849 13572
rect 5580 13364 5644 13428
rect 18276 13364 18340 13428
rect 6550 13084 6614 13088
rect 6550 13028 6554 13084
rect 6554 13028 6610 13084
rect 6610 13028 6614 13084
rect 6550 13024 6614 13028
rect 6630 13084 6694 13088
rect 6630 13028 6634 13084
rect 6634 13028 6690 13084
rect 6690 13028 6694 13084
rect 6630 13024 6694 13028
rect 6710 13084 6774 13088
rect 6710 13028 6714 13084
rect 6714 13028 6770 13084
rect 6770 13028 6774 13084
rect 6710 13024 6774 13028
rect 6790 13084 6854 13088
rect 6790 13028 6794 13084
rect 6794 13028 6850 13084
rect 6850 13028 6854 13084
rect 6790 13024 6854 13028
rect 12148 13084 12212 13088
rect 12148 13028 12152 13084
rect 12152 13028 12208 13084
rect 12208 13028 12212 13084
rect 12148 13024 12212 13028
rect 12228 13084 12292 13088
rect 12228 13028 12232 13084
rect 12232 13028 12288 13084
rect 12288 13028 12292 13084
rect 12228 13024 12292 13028
rect 12308 13084 12372 13088
rect 12308 13028 12312 13084
rect 12312 13028 12368 13084
rect 12368 13028 12372 13084
rect 12308 13024 12372 13028
rect 12388 13084 12452 13088
rect 12388 13028 12392 13084
rect 12392 13028 12448 13084
rect 12448 13028 12452 13084
rect 12388 13024 12452 13028
rect 17746 13084 17810 13088
rect 17746 13028 17750 13084
rect 17750 13028 17806 13084
rect 17806 13028 17810 13084
rect 17746 13024 17810 13028
rect 17826 13084 17890 13088
rect 17826 13028 17830 13084
rect 17830 13028 17886 13084
rect 17886 13028 17890 13084
rect 17826 13024 17890 13028
rect 17906 13084 17970 13088
rect 17906 13028 17910 13084
rect 17910 13028 17966 13084
rect 17966 13028 17970 13084
rect 17906 13024 17970 13028
rect 17986 13084 18050 13088
rect 17986 13028 17990 13084
rect 17990 13028 18046 13084
rect 18046 13028 18050 13084
rect 17986 13024 18050 13028
rect 4292 12820 4356 12884
rect 18828 12684 18892 12748
rect 3751 12540 3815 12544
rect 3751 12484 3755 12540
rect 3755 12484 3811 12540
rect 3811 12484 3815 12540
rect 3751 12480 3815 12484
rect 3831 12540 3895 12544
rect 3831 12484 3835 12540
rect 3835 12484 3891 12540
rect 3891 12484 3895 12540
rect 3831 12480 3895 12484
rect 3911 12540 3975 12544
rect 3911 12484 3915 12540
rect 3915 12484 3971 12540
rect 3971 12484 3975 12540
rect 3911 12480 3975 12484
rect 3991 12540 4055 12544
rect 3991 12484 3995 12540
rect 3995 12484 4051 12540
rect 4051 12484 4055 12540
rect 3991 12480 4055 12484
rect 9349 12540 9413 12544
rect 9349 12484 9353 12540
rect 9353 12484 9409 12540
rect 9409 12484 9413 12540
rect 9349 12480 9413 12484
rect 9429 12540 9493 12544
rect 9429 12484 9433 12540
rect 9433 12484 9489 12540
rect 9489 12484 9493 12540
rect 9429 12480 9493 12484
rect 9509 12540 9573 12544
rect 9509 12484 9513 12540
rect 9513 12484 9569 12540
rect 9569 12484 9573 12540
rect 9509 12480 9573 12484
rect 9589 12540 9653 12544
rect 9589 12484 9593 12540
rect 9593 12484 9649 12540
rect 9649 12484 9653 12540
rect 9589 12480 9653 12484
rect 14947 12540 15011 12544
rect 14947 12484 14951 12540
rect 14951 12484 15007 12540
rect 15007 12484 15011 12540
rect 14947 12480 15011 12484
rect 15027 12540 15091 12544
rect 15027 12484 15031 12540
rect 15031 12484 15087 12540
rect 15087 12484 15091 12540
rect 15027 12480 15091 12484
rect 15107 12540 15171 12544
rect 15107 12484 15111 12540
rect 15111 12484 15167 12540
rect 15167 12484 15171 12540
rect 15107 12480 15171 12484
rect 15187 12540 15251 12544
rect 15187 12484 15191 12540
rect 15191 12484 15247 12540
rect 15247 12484 15251 12540
rect 15187 12480 15251 12484
rect 20545 12540 20609 12544
rect 20545 12484 20549 12540
rect 20549 12484 20605 12540
rect 20605 12484 20609 12540
rect 20545 12480 20609 12484
rect 20625 12540 20689 12544
rect 20625 12484 20629 12540
rect 20629 12484 20685 12540
rect 20685 12484 20689 12540
rect 20625 12480 20689 12484
rect 20705 12540 20769 12544
rect 20705 12484 20709 12540
rect 20709 12484 20765 12540
rect 20765 12484 20769 12540
rect 20705 12480 20769 12484
rect 20785 12540 20849 12544
rect 20785 12484 20789 12540
rect 20789 12484 20845 12540
rect 20845 12484 20849 12540
rect 20785 12480 20849 12484
rect 18460 12276 18524 12340
rect 6550 11996 6614 12000
rect 6550 11940 6554 11996
rect 6554 11940 6610 11996
rect 6610 11940 6614 11996
rect 6550 11936 6614 11940
rect 6630 11996 6694 12000
rect 6630 11940 6634 11996
rect 6634 11940 6690 11996
rect 6690 11940 6694 11996
rect 6630 11936 6694 11940
rect 6710 11996 6774 12000
rect 6710 11940 6714 11996
rect 6714 11940 6770 11996
rect 6770 11940 6774 11996
rect 6710 11936 6774 11940
rect 6790 11996 6854 12000
rect 6790 11940 6794 11996
rect 6794 11940 6850 11996
rect 6850 11940 6854 11996
rect 6790 11936 6854 11940
rect 12148 11996 12212 12000
rect 12148 11940 12152 11996
rect 12152 11940 12208 11996
rect 12208 11940 12212 11996
rect 12148 11936 12212 11940
rect 12228 11996 12292 12000
rect 12228 11940 12232 11996
rect 12232 11940 12288 11996
rect 12288 11940 12292 11996
rect 12228 11936 12292 11940
rect 12308 11996 12372 12000
rect 12308 11940 12312 11996
rect 12312 11940 12368 11996
rect 12368 11940 12372 11996
rect 12308 11936 12372 11940
rect 12388 11996 12452 12000
rect 12388 11940 12392 11996
rect 12392 11940 12448 11996
rect 12448 11940 12452 11996
rect 12388 11936 12452 11940
rect 17746 11996 17810 12000
rect 17746 11940 17750 11996
rect 17750 11940 17806 11996
rect 17806 11940 17810 11996
rect 17746 11936 17810 11940
rect 17826 11996 17890 12000
rect 17826 11940 17830 11996
rect 17830 11940 17886 11996
rect 17886 11940 17890 11996
rect 17826 11936 17890 11940
rect 17906 11996 17970 12000
rect 17906 11940 17910 11996
rect 17910 11940 17966 11996
rect 17966 11940 17970 11996
rect 17906 11936 17970 11940
rect 17986 11996 18050 12000
rect 17986 11940 17990 11996
rect 17990 11940 18046 11996
rect 18046 11940 18050 11996
rect 17986 11936 18050 11940
rect 6316 11732 6380 11796
rect 3751 11452 3815 11456
rect 3751 11396 3755 11452
rect 3755 11396 3811 11452
rect 3811 11396 3815 11452
rect 3751 11392 3815 11396
rect 3831 11452 3895 11456
rect 3831 11396 3835 11452
rect 3835 11396 3891 11452
rect 3891 11396 3895 11452
rect 3831 11392 3895 11396
rect 3911 11452 3975 11456
rect 3911 11396 3915 11452
rect 3915 11396 3971 11452
rect 3971 11396 3975 11452
rect 3911 11392 3975 11396
rect 3991 11452 4055 11456
rect 3991 11396 3995 11452
rect 3995 11396 4051 11452
rect 4051 11396 4055 11452
rect 3991 11392 4055 11396
rect 9349 11452 9413 11456
rect 9349 11396 9353 11452
rect 9353 11396 9409 11452
rect 9409 11396 9413 11452
rect 9349 11392 9413 11396
rect 9429 11452 9493 11456
rect 9429 11396 9433 11452
rect 9433 11396 9489 11452
rect 9489 11396 9493 11452
rect 9429 11392 9493 11396
rect 9509 11452 9573 11456
rect 9509 11396 9513 11452
rect 9513 11396 9569 11452
rect 9569 11396 9573 11452
rect 9509 11392 9573 11396
rect 9589 11452 9653 11456
rect 9589 11396 9593 11452
rect 9593 11396 9649 11452
rect 9649 11396 9653 11452
rect 9589 11392 9653 11396
rect 14947 11452 15011 11456
rect 14947 11396 14951 11452
rect 14951 11396 15007 11452
rect 15007 11396 15011 11452
rect 14947 11392 15011 11396
rect 15027 11452 15091 11456
rect 15027 11396 15031 11452
rect 15031 11396 15087 11452
rect 15087 11396 15091 11452
rect 15027 11392 15091 11396
rect 15107 11452 15171 11456
rect 15107 11396 15111 11452
rect 15111 11396 15167 11452
rect 15167 11396 15171 11452
rect 15107 11392 15171 11396
rect 15187 11452 15251 11456
rect 15187 11396 15191 11452
rect 15191 11396 15247 11452
rect 15247 11396 15251 11452
rect 15187 11392 15251 11396
rect 20545 11452 20609 11456
rect 20545 11396 20549 11452
rect 20549 11396 20605 11452
rect 20605 11396 20609 11452
rect 20545 11392 20609 11396
rect 20625 11452 20689 11456
rect 20625 11396 20629 11452
rect 20629 11396 20685 11452
rect 20685 11396 20689 11452
rect 20625 11392 20689 11396
rect 20705 11452 20769 11456
rect 20705 11396 20709 11452
rect 20709 11396 20765 11452
rect 20765 11396 20769 11452
rect 20705 11392 20769 11396
rect 20785 11452 20849 11456
rect 20785 11396 20789 11452
rect 20789 11396 20845 11452
rect 20845 11396 20849 11452
rect 20785 11392 20849 11396
rect 19196 11188 19260 11252
rect 6550 10908 6614 10912
rect 6550 10852 6554 10908
rect 6554 10852 6610 10908
rect 6610 10852 6614 10908
rect 6550 10848 6614 10852
rect 6630 10908 6694 10912
rect 6630 10852 6634 10908
rect 6634 10852 6690 10908
rect 6690 10852 6694 10908
rect 6630 10848 6694 10852
rect 6710 10908 6774 10912
rect 6710 10852 6714 10908
rect 6714 10852 6770 10908
rect 6770 10852 6774 10908
rect 6710 10848 6774 10852
rect 6790 10908 6854 10912
rect 6790 10852 6794 10908
rect 6794 10852 6850 10908
rect 6850 10852 6854 10908
rect 6790 10848 6854 10852
rect 12148 10908 12212 10912
rect 12148 10852 12152 10908
rect 12152 10852 12208 10908
rect 12208 10852 12212 10908
rect 12148 10848 12212 10852
rect 12228 10908 12292 10912
rect 12228 10852 12232 10908
rect 12232 10852 12288 10908
rect 12288 10852 12292 10908
rect 12228 10848 12292 10852
rect 12308 10908 12372 10912
rect 12308 10852 12312 10908
rect 12312 10852 12368 10908
rect 12368 10852 12372 10908
rect 12308 10848 12372 10852
rect 12388 10908 12452 10912
rect 12388 10852 12392 10908
rect 12392 10852 12448 10908
rect 12448 10852 12452 10908
rect 12388 10848 12452 10852
rect 17746 10908 17810 10912
rect 17746 10852 17750 10908
rect 17750 10852 17806 10908
rect 17806 10852 17810 10908
rect 17746 10848 17810 10852
rect 17826 10908 17890 10912
rect 17826 10852 17830 10908
rect 17830 10852 17886 10908
rect 17886 10852 17890 10908
rect 17826 10848 17890 10852
rect 17906 10908 17970 10912
rect 17906 10852 17910 10908
rect 17910 10852 17966 10908
rect 17966 10852 17970 10908
rect 17906 10848 17970 10852
rect 17986 10908 18050 10912
rect 17986 10852 17990 10908
rect 17990 10852 18046 10908
rect 18046 10852 18050 10908
rect 17986 10848 18050 10852
rect 3751 10364 3815 10368
rect 3751 10308 3755 10364
rect 3755 10308 3811 10364
rect 3811 10308 3815 10364
rect 3751 10304 3815 10308
rect 3831 10364 3895 10368
rect 3831 10308 3835 10364
rect 3835 10308 3891 10364
rect 3891 10308 3895 10364
rect 3831 10304 3895 10308
rect 3911 10364 3975 10368
rect 3911 10308 3915 10364
rect 3915 10308 3971 10364
rect 3971 10308 3975 10364
rect 3911 10304 3975 10308
rect 3991 10364 4055 10368
rect 3991 10308 3995 10364
rect 3995 10308 4051 10364
rect 4051 10308 4055 10364
rect 3991 10304 4055 10308
rect 9349 10364 9413 10368
rect 9349 10308 9353 10364
rect 9353 10308 9409 10364
rect 9409 10308 9413 10364
rect 9349 10304 9413 10308
rect 9429 10364 9493 10368
rect 9429 10308 9433 10364
rect 9433 10308 9489 10364
rect 9489 10308 9493 10364
rect 9429 10304 9493 10308
rect 9509 10364 9573 10368
rect 9509 10308 9513 10364
rect 9513 10308 9569 10364
rect 9569 10308 9573 10364
rect 9509 10304 9573 10308
rect 9589 10364 9653 10368
rect 9589 10308 9593 10364
rect 9593 10308 9649 10364
rect 9649 10308 9653 10364
rect 9589 10304 9653 10308
rect 14947 10364 15011 10368
rect 14947 10308 14951 10364
rect 14951 10308 15007 10364
rect 15007 10308 15011 10364
rect 14947 10304 15011 10308
rect 15027 10364 15091 10368
rect 15027 10308 15031 10364
rect 15031 10308 15087 10364
rect 15087 10308 15091 10364
rect 15027 10304 15091 10308
rect 15107 10364 15171 10368
rect 15107 10308 15111 10364
rect 15111 10308 15167 10364
rect 15167 10308 15171 10364
rect 15107 10304 15171 10308
rect 15187 10364 15251 10368
rect 15187 10308 15191 10364
rect 15191 10308 15247 10364
rect 15247 10308 15251 10364
rect 15187 10304 15251 10308
rect 20545 10364 20609 10368
rect 20545 10308 20549 10364
rect 20549 10308 20605 10364
rect 20605 10308 20609 10364
rect 20545 10304 20609 10308
rect 20625 10364 20689 10368
rect 20625 10308 20629 10364
rect 20629 10308 20685 10364
rect 20685 10308 20689 10364
rect 20625 10304 20689 10308
rect 20705 10364 20769 10368
rect 20705 10308 20709 10364
rect 20709 10308 20765 10364
rect 20765 10308 20769 10364
rect 20705 10304 20769 10308
rect 20785 10364 20849 10368
rect 20785 10308 20789 10364
rect 20789 10308 20845 10364
rect 20845 10308 20849 10364
rect 20785 10304 20849 10308
rect 6550 9820 6614 9824
rect 6550 9764 6554 9820
rect 6554 9764 6610 9820
rect 6610 9764 6614 9820
rect 6550 9760 6614 9764
rect 6630 9820 6694 9824
rect 6630 9764 6634 9820
rect 6634 9764 6690 9820
rect 6690 9764 6694 9820
rect 6630 9760 6694 9764
rect 6710 9820 6774 9824
rect 6710 9764 6714 9820
rect 6714 9764 6770 9820
rect 6770 9764 6774 9820
rect 6710 9760 6774 9764
rect 6790 9820 6854 9824
rect 6790 9764 6794 9820
rect 6794 9764 6850 9820
rect 6850 9764 6854 9820
rect 6790 9760 6854 9764
rect 12148 9820 12212 9824
rect 12148 9764 12152 9820
rect 12152 9764 12208 9820
rect 12208 9764 12212 9820
rect 12148 9760 12212 9764
rect 12228 9820 12292 9824
rect 12228 9764 12232 9820
rect 12232 9764 12288 9820
rect 12288 9764 12292 9820
rect 12228 9760 12292 9764
rect 12308 9820 12372 9824
rect 12308 9764 12312 9820
rect 12312 9764 12368 9820
rect 12368 9764 12372 9820
rect 12308 9760 12372 9764
rect 12388 9820 12452 9824
rect 12388 9764 12392 9820
rect 12392 9764 12448 9820
rect 12448 9764 12452 9820
rect 12388 9760 12452 9764
rect 17746 9820 17810 9824
rect 17746 9764 17750 9820
rect 17750 9764 17806 9820
rect 17806 9764 17810 9820
rect 17746 9760 17810 9764
rect 17826 9820 17890 9824
rect 17826 9764 17830 9820
rect 17830 9764 17886 9820
rect 17886 9764 17890 9820
rect 17826 9760 17890 9764
rect 17906 9820 17970 9824
rect 17906 9764 17910 9820
rect 17910 9764 17966 9820
rect 17966 9764 17970 9820
rect 17906 9760 17970 9764
rect 17986 9820 18050 9824
rect 17986 9764 17990 9820
rect 17990 9764 18046 9820
rect 18046 9764 18050 9820
rect 17986 9760 18050 9764
rect 3751 9276 3815 9280
rect 3751 9220 3755 9276
rect 3755 9220 3811 9276
rect 3811 9220 3815 9276
rect 3751 9216 3815 9220
rect 3831 9276 3895 9280
rect 3831 9220 3835 9276
rect 3835 9220 3891 9276
rect 3891 9220 3895 9276
rect 3831 9216 3895 9220
rect 3911 9276 3975 9280
rect 3911 9220 3915 9276
rect 3915 9220 3971 9276
rect 3971 9220 3975 9276
rect 3911 9216 3975 9220
rect 3991 9276 4055 9280
rect 3991 9220 3995 9276
rect 3995 9220 4051 9276
rect 4051 9220 4055 9276
rect 3991 9216 4055 9220
rect 9349 9276 9413 9280
rect 9349 9220 9353 9276
rect 9353 9220 9409 9276
rect 9409 9220 9413 9276
rect 9349 9216 9413 9220
rect 9429 9276 9493 9280
rect 9429 9220 9433 9276
rect 9433 9220 9489 9276
rect 9489 9220 9493 9276
rect 9429 9216 9493 9220
rect 9509 9276 9573 9280
rect 9509 9220 9513 9276
rect 9513 9220 9569 9276
rect 9569 9220 9573 9276
rect 9509 9216 9573 9220
rect 9589 9276 9653 9280
rect 9589 9220 9593 9276
rect 9593 9220 9649 9276
rect 9649 9220 9653 9276
rect 9589 9216 9653 9220
rect 14947 9276 15011 9280
rect 14947 9220 14951 9276
rect 14951 9220 15007 9276
rect 15007 9220 15011 9276
rect 14947 9216 15011 9220
rect 15027 9276 15091 9280
rect 15027 9220 15031 9276
rect 15031 9220 15087 9276
rect 15087 9220 15091 9276
rect 15027 9216 15091 9220
rect 15107 9276 15171 9280
rect 15107 9220 15111 9276
rect 15111 9220 15167 9276
rect 15167 9220 15171 9276
rect 15107 9216 15171 9220
rect 15187 9276 15251 9280
rect 15187 9220 15191 9276
rect 15191 9220 15247 9276
rect 15247 9220 15251 9276
rect 15187 9216 15251 9220
rect 20545 9276 20609 9280
rect 20545 9220 20549 9276
rect 20549 9220 20605 9276
rect 20605 9220 20609 9276
rect 20545 9216 20609 9220
rect 20625 9276 20689 9280
rect 20625 9220 20629 9276
rect 20629 9220 20685 9276
rect 20685 9220 20689 9276
rect 20625 9216 20689 9220
rect 20705 9276 20769 9280
rect 20705 9220 20709 9276
rect 20709 9220 20765 9276
rect 20765 9220 20769 9276
rect 20705 9216 20769 9220
rect 20785 9276 20849 9280
rect 20785 9220 20789 9276
rect 20789 9220 20845 9276
rect 20845 9220 20849 9276
rect 20785 9216 20849 9220
rect 19012 8740 19076 8804
rect 6550 8732 6614 8736
rect 6550 8676 6554 8732
rect 6554 8676 6610 8732
rect 6610 8676 6614 8732
rect 6550 8672 6614 8676
rect 6630 8732 6694 8736
rect 6630 8676 6634 8732
rect 6634 8676 6690 8732
rect 6690 8676 6694 8732
rect 6630 8672 6694 8676
rect 6710 8732 6774 8736
rect 6710 8676 6714 8732
rect 6714 8676 6770 8732
rect 6770 8676 6774 8732
rect 6710 8672 6774 8676
rect 6790 8732 6854 8736
rect 6790 8676 6794 8732
rect 6794 8676 6850 8732
rect 6850 8676 6854 8732
rect 6790 8672 6854 8676
rect 12148 8732 12212 8736
rect 12148 8676 12152 8732
rect 12152 8676 12208 8732
rect 12208 8676 12212 8732
rect 12148 8672 12212 8676
rect 12228 8732 12292 8736
rect 12228 8676 12232 8732
rect 12232 8676 12288 8732
rect 12288 8676 12292 8732
rect 12228 8672 12292 8676
rect 12308 8732 12372 8736
rect 12308 8676 12312 8732
rect 12312 8676 12368 8732
rect 12368 8676 12372 8732
rect 12308 8672 12372 8676
rect 12388 8732 12452 8736
rect 12388 8676 12392 8732
rect 12392 8676 12448 8732
rect 12448 8676 12452 8732
rect 12388 8672 12452 8676
rect 17746 8732 17810 8736
rect 17746 8676 17750 8732
rect 17750 8676 17806 8732
rect 17806 8676 17810 8732
rect 17746 8672 17810 8676
rect 17826 8732 17890 8736
rect 17826 8676 17830 8732
rect 17830 8676 17886 8732
rect 17886 8676 17890 8732
rect 17826 8672 17890 8676
rect 17906 8732 17970 8736
rect 17906 8676 17910 8732
rect 17910 8676 17966 8732
rect 17966 8676 17970 8732
rect 17906 8672 17970 8676
rect 17986 8732 18050 8736
rect 17986 8676 17990 8732
rect 17990 8676 18046 8732
rect 18046 8676 18050 8732
rect 17986 8672 18050 8676
rect 16620 8332 16684 8396
rect 3751 8188 3815 8192
rect 3751 8132 3755 8188
rect 3755 8132 3811 8188
rect 3811 8132 3815 8188
rect 3751 8128 3815 8132
rect 3831 8188 3895 8192
rect 3831 8132 3835 8188
rect 3835 8132 3891 8188
rect 3891 8132 3895 8188
rect 3831 8128 3895 8132
rect 3911 8188 3975 8192
rect 3911 8132 3915 8188
rect 3915 8132 3971 8188
rect 3971 8132 3975 8188
rect 3911 8128 3975 8132
rect 3991 8188 4055 8192
rect 3991 8132 3995 8188
rect 3995 8132 4051 8188
rect 4051 8132 4055 8188
rect 3991 8128 4055 8132
rect 9349 8188 9413 8192
rect 9349 8132 9353 8188
rect 9353 8132 9409 8188
rect 9409 8132 9413 8188
rect 9349 8128 9413 8132
rect 9429 8188 9493 8192
rect 9429 8132 9433 8188
rect 9433 8132 9489 8188
rect 9489 8132 9493 8188
rect 9429 8128 9493 8132
rect 9509 8188 9573 8192
rect 9509 8132 9513 8188
rect 9513 8132 9569 8188
rect 9569 8132 9573 8188
rect 9509 8128 9573 8132
rect 9589 8188 9653 8192
rect 9589 8132 9593 8188
rect 9593 8132 9649 8188
rect 9649 8132 9653 8188
rect 9589 8128 9653 8132
rect 14947 8188 15011 8192
rect 14947 8132 14951 8188
rect 14951 8132 15007 8188
rect 15007 8132 15011 8188
rect 14947 8128 15011 8132
rect 15027 8188 15091 8192
rect 15027 8132 15031 8188
rect 15031 8132 15087 8188
rect 15087 8132 15091 8188
rect 15027 8128 15091 8132
rect 15107 8188 15171 8192
rect 15107 8132 15111 8188
rect 15111 8132 15167 8188
rect 15167 8132 15171 8188
rect 15107 8128 15171 8132
rect 15187 8188 15251 8192
rect 15187 8132 15191 8188
rect 15191 8132 15247 8188
rect 15247 8132 15251 8188
rect 15187 8128 15251 8132
rect 20545 8188 20609 8192
rect 20545 8132 20549 8188
rect 20549 8132 20605 8188
rect 20605 8132 20609 8188
rect 20545 8128 20609 8132
rect 20625 8188 20689 8192
rect 20625 8132 20629 8188
rect 20629 8132 20685 8188
rect 20685 8132 20689 8188
rect 20625 8128 20689 8132
rect 20705 8188 20769 8192
rect 20705 8132 20709 8188
rect 20709 8132 20765 8188
rect 20765 8132 20769 8188
rect 20705 8128 20769 8132
rect 20785 8188 20849 8192
rect 20785 8132 20789 8188
rect 20789 8132 20845 8188
rect 20845 8132 20849 8188
rect 20785 8128 20849 8132
rect 20300 7788 20364 7852
rect 21036 7652 21100 7716
rect 6550 7644 6614 7648
rect 6550 7588 6554 7644
rect 6554 7588 6610 7644
rect 6610 7588 6614 7644
rect 6550 7584 6614 7588
rect 6630 7644 6694 7648
rect 6630 7588 6634 7644
rect 6634 7588 6690 7644
rect 6690 7588 6694 7644
rect 6630 7584 6694 7588
rect 6710 7644 6774 7648
rect 6710 7588 6714 7644
rect 6714 7588 6770 7644
rect 6770 7588 6774 7644
rect 6710 7584 6774 7588
rect 6790 7644 6854 7648
rect 6790 7588 6794 7644
rect 6794 7588 6850 7644
rect 6850 7588 6854 7644
rect 6790 7584 6854 7588
rect 12148 7644 12212 7648
rect 12148 7588 12152 7644
rect 12152 7588 12208 7644
rect 12208 7588 12212 7644
rect 12148 7584 12212 7588
rect 12228 7644 12292 7648
rect 12228 7588 12232 7644
rect 12232 7588 12288 7644
rect 12288 7588 12292 7644
rect 12228 7584 12292 7588
rect 12308 7644 12372 7648
rect 12308 7588 12312 7644
rect 12312 7588 12368 7644
rect 12368 7588 12372 7644
rect 12308 7584 12372 7588
rect 12388 7644 12452 7648
rect 12388 7588 12392 7644
rect 12392 7588 12448 7644
rect 12448 7588 12452 7644
rect 12388 7584 12452 7588
rect 17746 7644 17810 7648
rect 17746 7588 17750 7644
rect 17750 7588 17806 7644
rect 17806 7588 17810 7644
rect 17746 7584 17810 7588
rect 17826 7644 17890 7648
rect 17826 7588 17830 7644
rect 17830 7588 17886 7644
rect 17886 7588 17890 7644
rect 17826 7584 17890 7588
rect 17906 7644 17970 7648
rect 17906 7588 17910 7644
rect 17910 7588 17966 7644
rect 17966 7588 17970 7644
rect 17906 7584 17970 7588
rect 17986 7644 18050 7648
rect 17986 7588 17990 7644
rect 17990 7588 18046 7644
rect 18046 7588 18050 7644
rect 17986 7584 18050 7588
rect 21404 7168 21468 7172
rect 21404 7112 21454 7168
rect 21454 7112 21468 7168
rect 21404 7108 21468 7112
rect 3751 7100 3815 7104
rect 3751 7044 3755 7100
rect 3755 7044 3811 7100
rect 3811 7044 3815 7100
rect 3751 7040 3815 7044
rect 3831 7100 3895 7104
rect 3831 7044 3835 7100
rect 3835 7044 3891 7100
rect 3891 7044 3895 7100
rect 3831 7040 3895 7044
rect 3911 7100 3975 7104
rect 3911 7044 3915 7100
rect 3915 7044 3971 7100
rect 3971 7044 3975 7100
rect 3911 7040 3975 7044
rect 3991 7100 4055 7104
rect 3991 7044 3995 7100
rect 3995 7044 4051 7100
rect 4051 7044 4055 7100
rect 3991 7040 4055 7044
rect 9349 7100 9413 7104
rect 9349 7044 9353 7100
rect 9353 7044 9409 7100
rect 9409 7044 9413 7100
rect 9349 7040 9413 7044
rect 9429 7100 9493 7104
rect 9429 7044 9433 7100
rect 9433 7044 9489 7100
rect 9489 7044 9493 7100
rect 9429 7040 9493 7044
rect 9509 7100 9573 7104
rect 9509 7044 9513 7100
rect 9513 7044 9569 7100
rect 9569 7044 9573 7100
rect 9509 7040 9573 7044
rect 9589 7100 9653 7104
rect 9589 7044 9593 7100
rect 9593 7044 9649 7100
rect 9649 7044 9653 7100
rect 9589 7040 9653 7044
rect 14947 7100 15011 7104
rect 14947 7044 14951 7100
rect 14951 7044 15007 7100
rect 15007 7044 15011 7100
rect 14947 7040 15011 7044
rect 15027 7100 15091 7104
rect 15027 7044 15031 7100
rect 15031 7044 15087 7100
rect 15087 7044 15091 7100
rect 15027 7040 15091 7044
rect 15107 7100 15171 7104
rect 15107 7044 15111 7100
rect 15111 7044 15167 7100
rect 15167 7044 15171 7100
rect 15107 7040 15171 7044
rect 15187 7100 15251 7104
rect 15187 7044 15191 7100
rect 15191 7044 15247 7100
rect 15247 7044 15251 7100
rect 15187 7040 15251 7044
rect 20545 7100 20609 7104
rect 20545 7044 20549 7100
rect 20549 7044 20605 7100
rect 20605 7044 20609 7100
rect 20545 7040 20609 7044
rect 20625 7100 20689 7104
rect 20625 7044 20629 7100
rect 20629 7044 20685 7100
rect 20685 7044 20689 7100
rect 20625 7040 20689 7044
rect 20705 7100 20769 7104
rect 20705 7044 20709 7100
rect 20709 7044 20765 7100
rect 20765 7044 20769 7100
rect 20705 7040 20769 7044
rect 20785 7100 20849 7104
rect 20785 7044 20789 7100
rect 20789 7044 20845 7100
rect 20845 7044 20849 7100
rect 20785 7040 20849 7044
rect 18644 6972 18708 7036
rect 22140 6972 22204 7036
rect 6550 6556 6614 6560
rect 6550 6500 6554 6556
rect 6554 6500 6610 6556
rect 6610 6500 6614 6556
rect 6550 6496 6614 6500
rect 6630 6556 6694 6560
rect 6630 6500 6634 6556
rect 6634 6500 6690 6556
rect 6690 6500 6694 6556
rect 6630 6496 6694 6500
rect 6710 6556 6774 6560
rect 6710 6500 6714 6556
rect 6714 6500 6770 6556
rect 6770 6500 6774 6556
rect 6710 6496 6774 6500
rect 6790 6556 6854 6560
rect 6790 6500 6794 6556
rect 6794 6500 6850 6556
rect 6850 6500 6854 6556
rect 6790 6496 6854 6500
rect 12148 6556 12212 6560
rect 12148 6500 12152 6556
rect 12152 6500 12208 6556
rect 12208 6500 12212 6556
rect 12148 6496 12212 6500
rect 12228 6556 12292 6560
rect 12228 6500 12232 6556
rect 12232 6500 12288 6556
rect 12288 6500 12292 6556
rect 12228 6496 12292 6500
rect 12308 6556 12372 6560
rect 12308 6500 12312 6556
rect 12312 6500 12368 6556
rect 12368 6500 12372 6556
rect 12308 6496 12372 6500
rect 12388 6556 12452 6560
rect 12388 6500 12392 6556
rect 12392 6500 12448 6556
rect 12448 6500 12452 6556
rect 12388 6496 12452 6500
rect 17746 6556 17810 6560
rect 17746 6500 17750 6556
rect 17750 6500 17806 6556
rect 17806 6500 17810 6556
rect 17746 6496 17810 6500
rect 17826 6556 17890 6560
rect 17826 6500 17830 6556
rect 17830 6500 17886 6556
rect 17886 6500 17890 6556
rect 17826 6496 17890 6500
rect 17906 6556 17970 6560
rect 17906 6500 17910 6556
rect 17910 6500 17966 6556
rect 17966 6500 17970 6556
rect 17906 6496 17970 6500
rect 17986 6556 18050 6560
rect 17986 6500 17990 6556
rect 17990 6500 18046 6556
rect 18046 6500 18050 6556
rect 17986 6496 18050 6500
rect 20300 6428 20364 6492
rect 21404 6292 21468 6356
rect 3751 6012 3815 6016
rect 3751 5956 3755 6012
rect 3755 5956 3811 6012
rect 3811 5956 3815 6012
rect 3751 5952 3815 5956
rect 3831 6012 3895 6016
rect 3831 5956 3835 6012
rect 3835 5956 3891 6012
rect 3891 5956 3895 6012
rect 3831 5952 3895 5956
rect 3911 6012 3975 6016
rect 3911 5956 3915 6012
rect 3915 5956 3971 6012
rect 3971 5956 3975 6012
rect 3911 5952 3975 5956
rect 3991 6012 4055 6016
rect 3991 5956 3995 6012
rect 3995 5956 4051 6012
rect 4051 5956 4055 6012
rect 3991 5952 4055 5956
rect 9349 6012 9413 6016
rect 9349 5956 9353 6012
rect 9353 5956 9409 6012
rect 9409 5956 9413 6012
rect 9349 5952 9413 5956
rect 9429 6012 9493 6016
rect 9429 5956 9433 6012
rect 9433 5956 9489 6012
rect 9489 5956 9493 6012
rect 9429 5952 9493 5956
rect 9509 6012 9573 6016
rect 9509 5956 9513 6012
rect 9513 5956 9569 6012
rect 9569 5956 9573 6012
rect 9509 5952 9573 5956
rect 9589 6012 9653 6016
rect 9589 5956 9593 6012
rect 9593 5956 9649 6012
rect 9649 5956 9653 6012
rect 9589 5952 9653 5956
rect 14947 6012 15011 6016
rect 14947 5956 14951 6012
rect 14951 5956 15007 6012
rect 15007 5956 15011 6012
rect 14947 5952 15011 5956
rect 15027 6012 15091 6016
rect 15027 5956 15031 6012
rect 15031 5956 15087 6012
rect 15087 5956 15091 6012
rect 15027 5952 15091 5956
rect 15107 6012 15171 6016
rect 15107 5956 15111 6012
rect 15111 5956 15167 6012
rect 15167 5956 15171 6012
rect 15107 5952 15171 5956
rect 15187 6012 15251 6016
rect 15187 5956 15191 6012
rect 15191 5956 15247 6012
rect 15247 5956 15251 6012
rect 15187 5952 15251 5956
rect 20545 6012 20609 6016
rect 20545 5956 20549 6012
rect 20549 5956 20605 6012
rect 20605 5956 20609 6012
rect 20545 5952 20609 5956
rect 20625 6012 20689 6016
rect 20625 5956 20629 6012
rect 20629 5956 20685 6012
rect 20685 5956 20689 6012
rect 20625 5952 20689 5956
rect 20705 6012 20769 6016
rect 20705 5956 20709 6012
rect 20709 5956 20765 6012
rect 20765 5956 20769 6012
rect 20705 5952 20769 5956
rect 20785 6012 20849 6016
rect 20785 5956 20789 6012
rect 20789 5956 20845 6012
rect 20845 5956 20849 6012
rect 20785 5952 20849 5956
rect 18644 5884 18708 5948
rect 22140 5884 22204 5948
rect 6550 5468 6614 5472
rect 6550 5412 6554 5468
rect 6554 5412 6610 5468
rect 6610 5412 6614 5468
rect 6550 5408 6614 5412
rect 6630 5468 6694 5472
rect 6630 5412 6634 5468
rect 6634 5412 6690 5468
rect 6690 5412 6694 5468
rect 6630 5408 6694 5412
rect 6710 5468 6774 5472
rect 6710 5412 6714 5468
rect 6714 5412 6770 5468
rect 6770 5412 6774 5468
rect 6710 5408 6774 5412
rect 6790 5468 6854 5472
rect 6790 5412 6794 5468
rect 6794 5412 6850 5468
rect 6850 5412 6854 5468
rect 6790 5408 6854 5412
rect 12148 5468 12212 5472
rect 12148 5412 12152 5468
rect 12152 5412 12208 5468
rect 12208 5412 12212 5468
rect 12148 5408 12212 5412
rect 12228 5468 12292 5472
rect 12228 5412 12232 5468
rect 12232 5412 12288 5468
rect 12288 5412 12292 5468
rect 12228 5408 12292 5412
rect 12308 5468 12372 5472
rect 12308 5412 12312 5468
rect 12312 5412 12368 5468
rect 12368 5412 12372 5468
rect 12308 5408 12372 5412
rect 12388 5468 12452 5472
rect 12388 5412 12392 5468
rect 12392 5412 12448 5468
rect 12448 5412 12452 5468
rect 12388 5408 12452 5412
rect 17746 5468 17810 5472
rect 17746 5412 17750 5468
rect 17750 5412 17806 5468
rect 17806 5412 17810 5468
rect 17746 5408 17810 5412
rect 17826 5468 17890 5472
rect 17826 5412 17830 5468
rect 17830 5412 17886 5468
rect 17886 5412 17890 5468
rect 17826 5408 17890 5412
rect 17906 5468 17970 5472
rect 17906 5412 17910 5468
rect 17910 5412 17966 5468
rect 17966 5412 17970 5468
rect 17906 5408 17970 5412
rect 17986 5468 18050 5472
rect 17986 5412 17990 5468
rect 17990 5412 18046 5468
rect 18046 5412 18050 5468
rect 17986 5408 18050 5412
rect 18828 5068 18892 5132
rect 3751 4924 3815 4928
rect 3751 4868 3755 4924
rect 3755 4868 3811 4924
rect 3811 4868 3815 4924
rect 3751 4864 3815 4868
rect 3831 4924 3895 4928
rect 3831 4868 3835 4924
rect 3835 4868 3891 4924
rect 3891 4868 3895 4924
rect 3831 4864 3895 4868
rect 3911 4924 3975 4928
rect 3911 4868 3915 4924
rect 3915 4868 3971 4924
rect 3971 4868 3975 4924
rect 3911 4864 3975 4868
rect 3991 4924 4055 4928
rect 3991 4868 3995 4924
rect 3995 4868 4051 4924
rect 4051 4868 4055 4924
rect 3991 4864 4055 4868
rect 9349 4924 9413 4928
rect 9349 4868 9353 4924
rect 9353 4868 9409 4924
rect 9409 4868 9413 4924
rect 9349 4864 9413 4868
rect 9429 4924 9493 4928
rect 9429 4868 9433 4924
rect 9433 4868 9489 4924
rect 9489 4868 9493 4924
rect 9429 4864 9493 4868
rect 9509 4924 9573 4928
rect 9509 4868 9513 4924
rect 9513 4868 9569 4924
rect 9569 4868 9573 4924
rect 9509 4864 9573 4868
rect 9589 4924 9653 4928
rect 9589 4868 9593 4924
rect 9593 4868 9649 4924
rect 9649 4868 9653 4924
rect 9589 4864 9653 4868
rect 14947 4924 15011 4928
rect 14947 4868 14951 4924
rect 14951 4868 15007 4924
rect 15007 4868 15011 4924
rect 14947 4864 15011 4868
rect 15027 4924 15091 4928
rect 15027 4868 15031 4924
rect 15031 4868 15087 4924
rect 15087 4868 15091 4924
rect 15027 4864 15091 4868
rect 15107 4924 15171 4928
rect 15107 4868 15111 4924
rect 15111 4868 15167 4924
rect 15167 4868 15171 4924
rect 15107 4864 15171 4868
rect 15187 4924 15251 4928
rect 15187 4868 15191 4924
rect 15191 4868 15247 4924
rect 15247 4868 15251 4924
rect 15187 4864 15251 4868
rect 20545 4924 20609 4928
rect 20545 4868 20549 4924
rect 20549 4868 20605 4924
rect 20605 4868 20609 4924
rect 20545 4864 20609 4868
rect 20625 4924 20689 4928
rect 20625 4868 20629 4924
rect 20629 4868 20685 4924
rect 20685 4868 20689 4924
rect 20625 4864 20689 4868
rect 20705 4924 20769 4928
rect 20705 4868 20709 4924
rect 20709 4868 20765 4924
rect 20765 4868 20769 4924
rect 20705 4864 20769 4868
rect 20785 4924 20849 4928
rect 20785 4868 20789 4924
rect 20789 4868 20845 4924
rect 20845 4868 20849 4924
rect 20785 4864 20849 4868
rect 19196 4660 19260 4724
rect 19012 4524 19076 4588
rect 6550 4380 6614 4384
rect 6550 4324 6554 4380
rect 6554 4324 6610 4380
rect 6610 4324 6614 4380
rect 6550 4320 6614 4324
rect 6630 4380 6694 4384
rect 6630 4324 6634 4380
rect 6634 4324 6690 4380
rect 6690 4324 6694 4380
rect 6630 4320 6694 4324
rect 6710 4380 6774 4384
rect 6710 4324 6714 4380
rect 6714 4324 6770 4380
rect 6770 4324 6774 4380
rect 6710 4320 6774 4324
rect 6790 4380 6854 4384
rect 6790 4324 6794 4380
rect 6794 4324 6850 4380
rect 6850 4324 6854 4380
rect 6790 4320 6854 4324
rect 12148 4380 12212 4384
rect 12148 4324 12152 4380
rect 12152 4324 12208 4380
rect 12208 4324 12212 4380
rect 12148 4320 12212 4324
rect 12228 4380 12292 4384
rect 12228 4324 12232 4380
rect 12232 4324 12288 4380
rect 12288 4324 12292 4380
rect 12228 4320 12292 4324
rect 12308 4380 12372 4384
rect 12308 4324 12312 4380
rect 12312 4324 12368 4380
rect 12368 4324 12372 4380
rect 12308 4320 12372 4324
rect 12388 4380 12452 4384
rect 12388 4324 12392 4380
rect 12392 4324 12448 4380
rect 12448 4324 12452 4380
rect 12388 4320 12452 4324
rect 17746 4380 17810 4384
rect 17746 4324 17750 4380
rect 17750 4324 17806 4380
rect 17806 4324 17810 4380
rect 17746 4320 17810 4324
rect 17826 4380 17890 4384
rect 17826 4324 17830 4380
rect 17830 4324 17886 4380
rect 17886 4324 17890 4380
rect 17826 4320 17890 4324
rect 17906 4380 17970 4384
rect 17906 4324 17910 4380
rect 17910 4324 17966 4380
rect 17966 4324 17970 4380
rect 17906 4320 17970 4324
rect 17986 4380 18050 4384
rect 17986 4324 17990 4380
rect 17990 4324 18046 4380
rect 18046 4324 18050 4380
rect 17986 4320 18050 4324
rect 17172 4116 17236 4180
rect 16620 4040 16684 4044
rect 16620 3984 16670 4040
rect 16670 3984 16684 4040
rect 16620 3980 16684 3984
rect 3751 3836 3815 3840
rect 3751 3780 3755 3836
rect 3755 3780 3811 3836
rect 3811 3780 3815 3836
rect 3751 3776 3815 3780
rect 3831 3836 3895 3840
rect 3831 3780 3835 3836
rect 3835 3780 3891 3836
rect 3891 3780 3895 3836
rect 3831 3776 3895 3780
rect 3911 3836 3975 3840
rect 3911 3780 3915 3836
rect 3915 3780 3971 3836
rect 3971 3780 3975 3836
rect 3911 3776 3975 3780
rect 3991 3836 4055 3840
rect 3991 3780 3995 3836
rect 3995 3780 4051 3836
rect 4051 3780 4055 3836
rect 3991 3776 4055 3780
rect 9349 3836 9413 3840
rect 9349 3780 9353 3836
rect 9353 3780 9409 3836
rect 9409 3780 9413 3836
rect 9349 3776 9413 3780
rect 9429 3836 9493 3840
rect 9429 3780 9433 3836
rect 9433 3780 9489 3836
rect 9489 3780 9493 3836
rect 9429 3776 9493 3780
rect 9509 3836 9573 3840
rect 9509 3780 9513 3836
rect 9513 3780 9569 3836
rect 9569 3780 9573 3836
rect 9509 3776 9573 3780
rect 9589 3836 9653 3840
rect 9589 3780 9593 3836
rect 9593 3780 9649 3836
rect 9649 3780 9653 3836
rect 9589 3776 9653 3780
rect 14947 3836 15011 3840
rect 14947 3780 14951 3836
rect 14951 3780 15007 3836
rect 15007 3780 15011 3836
rect 14947 3776 15011 3780
rect 15027 3836 15091 3840
rect 15027 3780 15031 3836
rect 15031 3780 15087 3836
rect 15087 3780 15091 3836
rect 15027 3776 15091 3780
rect 15107 3836 15171 3840
rect 15107 3780 15111 3836
rect 15111 3780 15167 3836
rect 15167 3780 15171 3836
rect 15107 3776 15171 3780
rect 15187 3836 15251 3840
rect 15187 3780 15191 3836
rect 15191 3780 15247 3836
rect 15247 3780 15251 3836
rect 15187 3776 15251 3780
rect 20545 3836 20609 3840
rect 20545 3780 20549 3836
rect 20549 3780 20605 3836
rect 20605 3780 20609 3836
rect 20545 3776 20609 3780
rect 20625 3836 20689 3840
rect 20625 3780 20629 3836
rect 20629 3780 20685 3836
rect 20685 3780 20689 3836
rect 20625 3776 20689 3780
rect 20705 3836 20769 3840
rect 20705 3780 20709 3836
rect 20709 3780 20765 3836
rect 20765 3780 20769 3836
rect 20705 3776 20769 3780
rect 20785 3836 20849 3840
rect 20785 3780 20789 3836
rect 20789 3780 20845 3836
rect 20845 3780 20849 3836
rect 20785 3776 20849 3780
rect 21036 3708 21100 3772
rect 6550 3292 6614 3296
rect 6550 3236 6554 3292
rect 6554 3236 6610 3292
rect 6610 3236 6614 3292
rect 6550 3232 6614 3236
rect 6630 3292 6694 3296
rect 6630 3236 6634 3292
rect 6634 3236 6690 3292
rect 6690 3236 6694 3292
rect 6630 3232 6694 3236
rect 6710 3292 6774 3296
rect 6710 3236 6714 3292
rect 6714 3236 6770 3292
rect 6770 3236 6774 3292
rect 6710 3232 6774 3236
rect 6790 3292 6854 3296
rect 6790 3236 6794 3292
rect 6794 3236 6850 3292
rect 6850 3236 6854 3292
rect 6790 3232 6854 3236
rect 12148 3292 12212 3296
rect 12148 3236 12152 3292
rect 12152 3236 12208 3292
rect 12208 3236 12212 3292
rect 12148 3232 12212 3236
rect 12228 3292 12292 3296
rect 12228 3236 12232 3292
rect 12232 3236 12288 3292
rect 12288 3236 12292 3292
rect 12228 3232 12292 3236
rect 12308 3292 12372 3296
rect 12308 3236 12312 3292
rect 12312 3236 12368 3292
rect 12368 3236 12372 3292
rect 12308 3232 12372 3236
rect 12388 3292 12452 3296
rect 12388 3236 12392 3292
rect 12392 3236 12448 3292
rect 12448 3236 12452 3292
rect 12388 3232 12452 3236
rect 17746 3292 17810 3296
rect 17746 3236 17750 3292
rect 17750 3236 17806 3292
rect 17806 3236 17810 3292
rect 17746 3232 17810 3236
rect 17826 3292 17890 3296
rect 17826 3236 17830 3292
rect 17830 3236 17886 3292
rect 17886 3236 17890 3292
rect 17826 3232 17890 3236
rect 17906 3292 17970 3296
rect 17906 3236 17910 3292
rect 17910 3236 17966 3292
rect 17966 3236 17970 3292
rect 17906 3232 17970 3236
rect 17986 3292 18050 3296
rect 17986 3236 17990 3292
rect 17990 3236 18046 3292
rect 18046 3236 18050 3292
rect 17986 3232 18050 3236
rect 3751 2748 3815 2752
rect 3751 2692 3755 2748
rect 3755 2692 3811 2748
rect 3811 2692 3815 2748
rect 3751 2688 3815 2692
rect 3831 2748 3895 2752
rect 3831 2692 3835 2748
rect 3835 2692 3891 2748
rect 3891 2692 3895 2748
rect 3831 2688 3895 2692
rect 3911 2748 3975 2752
rect 3911 2692 3915 2748
rect 3915 2692 3971 2748
rect 3971 2692 3975 2748
rect 3911 2688 3975 2692
rect 3991 2748 4055 2752
rect 3991 2692 3995 2748
rect 3995 2692 4051 2748
rect 4051 2692 4055 2748
rect 3991 2688 4055 2692
rect 9349 2748 9413 2752
rect 9349 2692 9353 2748
rect 9353 2692 9409 2748
rect 9409 2692 9413 2748
rect 9349 2688 9413 2692
rect 9429 2748 9493 2752
rect 9429 2692 9433 2748
rect 9433 2692 9489 2748
rect 9489 2692 9493 2748
rect 9429 2688 9493 2692
rect 9509 2748 9573 2752
rect 9509 2692 9513 2748
rect 9513 2692 9569 2748
rect 9569 2692 9573 2748
rect 9509 2688 9573 2692
rect 9589 2748 9653 2752
rect 9589 2692 9593 2748
rect 9593 2692 9649 2748
rect 9649 2692 9653 2748
rect 9589 2688 9653 2692
rect 14947 2748 15011 2752
rect 14947 2692 14951 2748
rect 14951 2692 15007 2748
rect 15007 2692 15011 2748
rect 14947 2688 15011 2692
rect 15027 2748 15091 2752
rect 15027 2692 15031 2748
rect 15031 2692 15087 2748
rect 15087 2692 15091 2748
rect 15027 2688 15091 2692
rect 15107 2748 15171 2752
rect 15107 2692 15111 2748
rect 15111 2692 15167 2748
rect 15167 2692 15171 2748
rect 15107 2688 15171 2692
rect 15187 2748 15251 2752
rect 15187 2692 15191 2748
rect 15191 2692 15247 2748
rect 15247 2692 15251 2748
rect 15187 2688 15251 2692
rect 20545 2748 20609 2752
rect 20545 2692 20549 2748
rect 20549 2692 20605 2748
rect 20605 2692 20609 2748
rect 20545 2688 20609 2692
rect 20625 2748 20689 2752
rect 20625 2692 20629 2748
rect 20629 2692 20685 2748
rect 20685 2692 20689 2748
rect 20625 2688 20689 2692
rect 20705 2748 20769 2752
rect 20705 2692 20709 2748
rect 20709 2692 20765 2748
rect 20765 2692 20769 2748
rect 20705 2688 20769 2692
rect 20785 2748 20849 2752
rect 20785 2692 20789 2748
rect 20789 2692 20845 2748
rect 20845 2692 20849 2748
rect 20785 2688 20849 2692
rect 6550 2204 6614 2208
rect 6550 2148 6554 2204
rect 6554 2148 6610 2204
rect 6610 2148 6614 2204
rect 6550 2144 6614 2148
rect 6630 2204 6694 2208
rect 6630 2148 6634 2204
rect 6634 2148 6690 2204
rect 6690 2148 6694 2204
rect 6630 2144 6694 2148
rect 6710 2204 6774 2208
rect 6710 2148 6714 2204
rect 6714 2148 6770 2204
rect 6770 2148 6774 2204
rect 6710 2144 6774 2148
rect 6790 2204 6854 2208
rect 6790 2148 6794 2204
rect 6794 2148 6850 2204
rect 6850 2148 6854 2204
rect 6790 2144 6854 2148
rect 12148 2204 12212 2208
rect 12148 2148 12152 2204
rect 12152 2148 12208 2204
rect 12208 2148 12212 2204
rect 12148 2144 12212 2148
rect 12228 2204 12292 2208
rect 12228 2148 12232 2204
rect 12232 2148 12288 2204
rect 12288 2148 12292 2204
rect 12228 2144 12292 2148
rect 12308 2204 12372 2208
rect 12308 2148 12312 2204
rect 12312 2148 12368 2204
rect 12368 2148 12372 2204
rect 12308 2144 12372 2148
rect 12388 2204 12452 2208
rect 12388 2148 12392 2204
rect 12392 2148 12448 2204
rect 12448 2148 12452 2204
rect 12388 2144 12452 2148
rect 17746 2204 17810 2208
rect 17746 2148 17750 2204
rect 17750 2148 17806 2204
rect 17806 2148 17810 2204
rect 17746 2144 17810 2148
rect 17826 2204 17890 2208
rect 17826 2148 17830 2204
rect 17830 2148 17886 2204
rect 17886 2148 17890 2204
rect 17826 2144 17890 2148
rect 17906 2204 17970 2208
rect 17906 2148 17910 2204
rect 17910 2148 17966 2204
rect 17966 2148 17970 2204
rect 17906 2144 17970 2148
rect 17986 2204 18050 2208
rect 17986 2148 17990 2204
rect 17990 2148 18046 2204
rect 18046 2148 18050 2204
rect 17986 2144 18050 2148
<< metal4 >>
rect 3743 22336 4063 22352
rect 3743 22272 3751 22336
rect 3815 22272 3831 22336
rect 3895 22272 3911 22336
rect 3975 22272 3991 22336
rect 4055 22272 4063 22336
rect 3743 21248 4063 22272
rect 5579 21996 5645 21997
rect 5579 21932 5580 21996
rect 5644 21932 5645 21996
rect 5579 21931 5645 21932
rect 3743 21184 3751 21248
rect 3815 21184 3831 21248
rect 3895 21184 3911 21248
rect 3975 21184 3991 21248
rect 4055 21184 4063 21248
rect 3743 20160 4063 21184
rect 4843 20908 4909 20909
rect 4843 20844 4844 20908
rect 4908 20844 4909 20908
rect 4843 20843 4909 20844
rect 3743 20096 3751 20160
rect 3815 20096 3831 20160
rect 3895 20096 3911 20160
rect 3975 20096 3991 20160
rect 4055 20096 4063 20160
rect 3743 19072 4063 20096
rect 3743 19008 3751 19072
rect 3815 19008 3831 19072
rect 3895 19008 3911 19072
rect 3975 19008 3991 19072
rect 4055 19008 4063 19072
rect 3743 17984 4063 19008
rect 3743 17920 3751 17984
rect 3815 17920 3831 17984
rect 3895 17920 3911 17984
rect 3975 17920 3991 17984
rect 4055 17920 4063 17984
rect 3743 16896 4063 17920
rect 3743 16832 3751 16896
rect 3815 16832 3831 16896
rect 3895 16832 3911 16896
rect 3975 16832 3991 16896
rect 4055 16832 4063 16896
rect 3743 15808 4063 16832
rect 3743 15744 3751 15808
rect 3815 15744 3831 15808
rect 3895 15744 3911 15808
rect 3975 15744 3991 15808
rect 4055 15744 4063 15808
rect 3743 14720 4063 15744
rect 4291 15332 4357 15333
rect 4291 15268 4292 15332
rect 4356 15268 4357 15332
rect 4291 15267 4357 15268
rect 3743 14656 3751 14720
rect 3815 14656 3831 14720
rect 3895 14656 3911 14720
rect 3975 14656 3991 14720
rect 4055 14656 4063 14720
rect 3743 13632 4063 14656
rect 3743 13568 3751 13632
rect 3815 13568 3831 13632
rect 3895 13568 3911 13632
rect 3975 13568 3991 13632
rect 4055 13568 4063 13632
rect 3743 12544 4063 13568
rect 4294 12885 4354 15267
rect 4846 15061 4906 20843
rect 4843 15060 4909 15061
rect 4843 14996 4844 15060
rect 4908 14996 4909 15060
rect 4843 14995 4909 14996
rect 5582 13429 5642 21931
rect 6542 21792 6862 22352
rect 6542 21728 6550 21792
rect 6614 21728 6630 21792
rect 6694 21728 6710 21792
rect 6774 21728 6790 21792
rect 6854 21728 6862 21792
rect 6315 20908 6381 20909
rect 6315 20844 6316 20908
rect 6380 20844 6381 20908
rect 6315 20843 6381 20844
rect 5579 13428 5645 13429
rect 5579 13364 5580 13428
rect 5644 13364 5645 13428
rect 5579 13363 5645 13364
rect 4291 12884 4357 12885
rect 4291 12820 4292 12884
rect 4356 12820 4357 12884
rect 4291 12819 4357 12820
rect 3743 12480 3751 12544
rect 3815 12480 3831 12544
rect 3895 12480 3911 12544
rect 3975 12480 3991 12544
rect 4055 12480 4063 12544
rect 3743 11456 4063 12480
rect 6318 11797 6378 20843
rect 6542 20704 6862 21728
rect 6542 20640 6550 20704
rect 6614 20640 6630 20704
rect 6694 20640 6710 20704
rect 6774 20640 6790 20704
rect 6854 20640 6862 20704
rect 6542 19616 6862 20640
rect 6542 19552 6550 19616
rect 6614 19552 6630 19616
rect 6694 19552 6710 19616
rect 6774 19552 6790 19616
rect 6854 19552 6862 19616
rect 6542 18528 6862 19552
rect 6542 18464 6550 18528
rect 6614 18464 6630 18528
rect 6694 18464 6710 18528
rect 6774 18464 6790 18528
rect 6854 18464 6862 18528
rect 6542 17440 6862 18464
rect 6542 17376 6550 17440
rect 6614 17376 6630 17440
rect 6694 17376 6710 17440
rect 6774 17376 6790 17440
rect 6854 17376 6862 17440
rect 6542 16352 6862 17376
rect 6542 16288 6550 16352
rect 6614 16288 6630 16352
rect 6694 16288 6710 16352
rect 6774 16288 6790 16352
rect 6854 16288 6862 16352
rect 6542 15264 6862 16288
rect 6542 15200 6550 15264
rect 6614 15200 6630 15264
rect 6694 15200 6710 15264
rect 6774 15200 6790 15264
rect 6854 15200 6862 15264
rect 6542 14176 6862 15200
rect 6542 14112 6550 14176
rect 6614 14112 6630 14176
rect 6694 14112 6710 14176
rect 6774 14112 6790 14176
rect 6854 14112 6862 14176
rect 6542 13088 6862 14112
rect 6542 13024 6550 13088
rect 6614 13024 6630 13088
rect 6694 13024 6710 13088
rect 6774 13024 6790 13088
rect 6854 13024 6862 13088
rect 6542 12000 6862 13024
rect 6542 11936 6550 12000
rect 6614 11936 6630 12000
rect 6694 11936 6710 12000
rect 6774 11936 6790 12000
rect 6854 11936 6862 12000
rect 6315 11796 6381 11797
rect 6315 11732 6316 11796
rect 6380 11732 6381 11796
rect 6315 11731 6381 11732
rect 3743 11392 3751 11456
rect 3815 11392 3831 11456
rect 3895 11392 3911 11456
rect 3975 11392 3991 11456
rect 4055 11392 4063 11456
rect 3743 10368 4063 11392
rect 3743 10304 3751 10368
rect 3815 10304 3831 10368
rect 3895 10304 3911 10368
rect 3975 10304 3991 10368
rect 4055 10304 4063 10368
rect 3743 9280 4063 10304
rect 3743 9216 3751 9280
rect 3815 9216 3831 9280
rect 3895 9216 3911 9280
rect 3975 9216 3991 9280
rect 4055 9216 4063 9280
rect 3743 8192 4063 9216
rect 3743 8128 3751 8192
rect 3815 8128 3831 8192
rect 3895 8128 3911 8192
rect 3975 8128 3991 8192
rect 4055 8128 4063 8192
rect 3743 7104 4063 8128
rect 3743 7040 3751 7104
rect 3815 7040 3831 7104
rect 3895 7040 3911 7104
rect 3975 7040 3991 7104
rect 4055 7040 4063 7104
rect 3743 6016 4063 7040
rect 3743 5952 3751 6016
rect 3815 5952 3831 6016
rect 3895 5952 3911 6016
rect 3975 5952 3991 6016
rect 4055 5952 4063 6016
rect 3743 4928 4063 5952
rect 3743 4864 3751 4928
rect 3815 4864 3831 4928
rect 3895 4864 3911 4928
rect 3975 4864 3991 4928
rect 4055 4864 4063 4928
rect 3743 3840 4063 4864
rect 3743 3776 3751 3840
rect 3815 3776 3831 3840
rect 3895 3776 3911 3840
rect 3975 3776 3991 3840
rect 4055 3776 4063 3840
rect 3743 2752 4063 3776
rect 3743 2688 3751 2752
rect 3815 2688 3831 2752
rect 3895 2688 3911 2752
rect 3975 2688 3991 2752
rect 4055 2688 4063 2752
rect 3743 2128 4063 2688
rect 6542 10912 6862 11936
rect 6542 10848 6550 10912
rect 6614 10848 6630 10912
rect 6694 10848 6710 10912
rect 6774 10848 6790 10912
rect 6854 10848 6862 10912
rect 6542 9824 6862 10848
rect 6542 9760 6550 9824
rect 6614 9760 6630 9824
rect 6694 9760 6710 9824
rect 6774 9760 6790 9824
rect 6854 9760 6862 9824
rect 6542 8736 6862 9760
rect 6542 8672 6550 8736
rect 6614 8672 6630 8736
rect 6694 8672 6710 8736
rect 6774 8672 6790 8736
rect 6854 8672 6862 8736
rect 6542 7648 6862 8672
rect 6542 7584 6550 7648
rect 6614 7584 6630 7648
rect 6694 7584 6710 7648
rect 6774 7584 6790 7648
rect 6854 7584 6862 7648
rect 6542 6560 6862 7584
rect 6542 6496 6550 6560
rect 6614 6496 6630 6560
rect 6694 6496 6710 6560
rect 6774 6496 6790 6560
rect 6854 6496 6862 6560
rect 6542 5472 6862 6496
rect 6542 5408 6550 5472
rect 6614 5408 6630 5472
rect 6694 5408 6710 5472
rect 6774 5408 6790 5472
rect 6854 5408 6862 5472
rect 6542 4384 6862 5408
rect 6542 4320 6550 4384
rect 6614 4320 6630 4384
rect 6694 4320 6710 4384
rect 6774 4320 6790 4384
rect 6854 4320 6862 4384
rect 6542 3296 6862 4320
rect 6542 3232 6550 3296
rect 6614 3232 6630 3296
rect 6694 3232 6710 3296
rect 6774 3232 6790 3296
rect 6854 3232 6862 3296
rect 6542 2208 6862 3232
rect 6542 2144 6550 2208
rect 6614 2144 6630 2208
rect 6694 2144 6710 2208
rect 6774 2144 6790 2208
rect 6854 2144 6862 2208
rect 6542 2128 6862 2144
rect 9341 22336 9661 22352
rect 9341 22272 9349 22336
rect 9413 22272 9429 22336
rect 9493 22272 9509 22336
rect 9573 22272 9589 22336
rect 9653 22272 9661 22336
rect 9341 21248 9661 22272
rect 9341 21184 9349 21248
rect 9413 21184 9429 21248
rect 9493 21184 9509 21248
rect 9573 21184 9589 21248
rect 9653 21184 9661 21248
rect 9341 20160 9661 21184
rect 9341 20096 9349 20160
rect 9413 20096 9429 20160
rect 9493 20096 9509 20160
rect 9573 20096 9589 20160
rect 9653 20096 9661 20160
rect 9341 19072 9661 20096
rect 9341 19008 9349 19072
rect 9413 19008 9429 19072
rect 9493 19008 9509 19072
rect 9573 19008 9589 19072
rect 9653 19008 9661 19072
rect 9341 17984 9661 19008
rect 9341 17920 9349 17984
rect 9413 17920 9429 17984
rect 9493 17920 9509 17984
rect 9573 17920 9589 17984
rect 9653 17920 9661 17984
rect 9341 16896 9661 17920
rect 9341 16832 9349 16896
rect 9413 16832 9429 16896
rect 9493 16832 9509 16896
rect 9573 16832 9589 16896
rect 9653 16832 9661 16896
rect 9341 15808 9661 16832
rect 9341 15744 9349 15808
rect 9413 15744 9429 15808
rect 9493 15744 9509 15808
rect 9573 15744 9589 15808
rect 9653 15744 9661 15808
rect 9341 14720 9661 15744
rect 9341 14656 9349 14720
rect 9413 14656 9429 14720
rect 9493 14656 9509 14720
rect 9573 14656 9589 14720
rect 9653 14656 9661 14720
rect 9341 13632 9661 14656
rect 9341 13568 9349 13632
rect 9413 13568 9429 13632
rect 9493 13568 9509 13632
rect 9573 13568 9589 13632
rect 9653 13568 9661 13632
rect 9341 12544 9661 13568
rect 9341 12480 9349 12544
rect 9413 12480 9429 12544
rect 9493 12480 9509 12544
rect 9573 12480 9589 12544
rect 9653 12480 9661 12544
rect 9341 11456 9661 12480
rect 9341 11392 9349 11456
rect 9413 11392 9429 11456
rect 9493 11392 9509 11456
rect 9573 11392 9589 11456
rect 9653 11392 9661 11456
rect 9341 10368 9661 11392
rect 9341 10304 9349 10368
rect 9413 10304 9429 10368
rect 9493 10304 9509 10368
rect 9573 10304 9589 10368
rect 9653 10304 9661 10368
rect 9341 9280 9661 10304
rect 9341 9216 9349 9280
rect 9413 9216 9429 9280
rect 9493 9216 9509 9280
rect 9573 9216 9589 9280
rect 9653 9216 9661 9280
rect 9341 8192 9661 9216
rect 9341 8128 9349 8192
rect 9413 8128 9429 8192
rect 9493 8128 9509 8192
rect 9573 8128 9589 8192
rect 9653 8128 9661 8192
rect 9341 7104 9661 8128
rect 9341 7040 9349 7104
rect 9413 7040 9429 7104
rect 9493 7040 9509 7104
rect 9573 7040 9589 7104
rect 9653 7040 9661 7104
rect 9341 6016 9661 7040
rect 9341 5952 9349 6016
rect 9413 5952 9429 6016
rect 9493 5952 9509 6016
rect 9573 5952 9589 6016
rect 9653 5952 9661 6016
rect 9341 4928 9661 5952
rect 9341 4864 9349 4928
rect 9413 4864 9429 4928
rect 9493 4864 9509 4928
rect 9573 4864 9589 4928
rect 9653 4864 9661 4928
rect 9341 3840 9661 4864
rect 9341 3776 9349 3840
rect 9413 3776 9429 3840
rect 9493 3776 9509 3840
rect 9573 3776 9589 3840
rect 9653 3776 9661 3840
rect 9341 2752 9661 3776
rect 9341 2688 9349 2752
rect 9413 2688 9429 2752
rect 9493 2688 9509 2752
rect 9573 2688 9589 2752
rect 9653 2688 9661 2752
rect 9341 2128 9661 2688
rect 12140 21792 12460 22352
rect 14939 22336 15259 22352
rect 14939 22272 14947 22336
rect 15011 22272 15027 22336
rect 15091 22272 15107 22336
rect 15171 22272 15187 22336
rect 15251 22272 15259 22336
rect 13307 21860 13373 21861
rect 13307 21796 13308 21860
rect 13372 21796 13373 21860
rect 13307 21795 13373 21796
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 20704 12460 21728
rect 12571 21044 12637 21045
rect 12571 20980 12572 21044
rect 12636 20980 12637 21044
rect 12571 20979 12637 20980
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 19616 12460 20640
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 18528 12460 19552
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 17440 12460 18464
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 16352 12460 17376
rect 12574 16557 12634 20979
rect 13310 18869 13370 21795
rect 14939 21248 15259 22272
rect 17738 21792 18058 22352
rect 20537 22336 20857 22352
rect 20537 22272 20545 22336
rect 20609 22272 20625 22336
rect 20689 22272 20705 22336
rect 20769 22272 20785 22336
rect 20849 22272 20857 22336
rect 18275 21860 18341 21861
rect 18275 21796 18276 21860
rect 18340 21796 18341 21860
rect 18275 21795 18341 21796
rect 17738 21728 17746 21792
rect 17810 21728 17826 21792
rect 17890 21728 17906 21792
rect 17970 21728 17986 21792
rect 18050 21728 18058 21792
rect 15331 21724 15397 21725
rect 15331 21660 15332 21724
rect 15396 21660 15397 21724
rect 15331 21659 15397 21660
rect 14939 21184 14947 21248
rect 15011 21184 15027 21248
rect 15091 21184 15107 21248
rect 15171 21184 15187 21248
rect 15251 21184 15259 21248
rect 14939 20160 15259 21184
rect 14939 20096 14947 20160
rect 15011 20096 15027 20160
rect 15091 20096 15107 20160
rect 15171 20096 15187 20160
rect 15251 20096 15259 20160
rect 14939 19072 15259 20096
rect 14939 19008 14947 19072
rect 15011 19008 15027 19072
rect 15091 19008 15107 19072
rect 15171 19008 15187 19072
rect 15251 19008 15259 19072
rect 13307 18868 13373 18869
rect 13307 18804 13308 18868
rect 13372 18804 13373 18868
rect 13307 18803 13373 18804
rect 14939 17984 15259 19008
rect 14939 17920 14947 17984
rect 15011 17920 15027 17984
rect 15091 17920 15107 17984
rect 15171 17920 15187 17984
rect 15251 17920 15259 17984
rect 14939 16896 15259 17920
rect 15334 17645 15394 21659
rect 17738 20704 18058 21728
rect 17738 20640 17746 20704
rect 17810 20640 17826 20704
rect 17890 20640 17906 20704
rect 17970 20640 17986 20704
rect 18050 20640 18058 20704
rect 16987 20500 17053 20501
rect 16987 20436 16988 20500
rect 17052 20436 17053 20500
rect 16987 20435 17053 20436
rect 16435 20092 16501 20093
rect 16435 20028 16436 20092
rect 16500 20028 16501 20092
rect 16435 20027 16501 20028
rect 16438 19549 16498 20027
rect 16435 19548 16501 19549
rect 16435 19484 16436 19548
rect 16500 19484 16501 19548
rect 16435 19483 16501 19484
rect 16990 19413 17050 20435
rect 17738 19616 18058 20640
rect 17738 19552 17746 19616
rect 17810 19552 17826 19616
rect 17890 19552 17906 19616
rect 17970 19552 17986 19616
rect 18050 19552 18058 19616
rect 16619 19412 16685 19413
rect 16619 19348 16620 19412
rect 16684 19348 16685 19412
rect 16619 19347 16685 19348
rect 16987 19412 17053 19413
rect 16987 19348 16988 19412
rect 17052 19348 17053 19412
rect 16987 19347 17053 19348
rect 15331 17644 15397 17645
rect 15331 17580 15332 17644
rect 15396 17580 15397 17644
rect 15331 17579 15397 17580
rect 14939 16832 14947 16896
rect 15011 16832 15027 16896
rect 15091 16832 15107 16896
rect 15171 16832 15187 16896
rect 15251 16832 15259 16896
rect 12571 16556 12637 16557
rect 12571 16492 12572 16556
rect 12636 16492 12637 16556
rect 12571 16491 12637 16492
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 15264 12460 16288
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 14176 12460 15200
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 13088 12460 14112
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 12000 12460 13024
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 10912 12460 11936
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 9824 12460 10848
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 8736 12460 9760
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 7648 12460 8672
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 6560 12460 7584
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 5472 12460 6496
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 4384 12460 5408
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 3296 12460 4320
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 2208 12460 3232
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2128 12460 2144
rect 14939 15808 15259 16832
rect 14939 15744 14947 15808
rect 15011 15744 15027 15808
rect 15091 15744 15107 15808
rect 15171 15744 15187 15808
rect 15251 15744 15259 15808
rect 14939 14720 15259 15744
rect 16622 15197 16682 19347
rect 17738 18528 18058 19552
rect 17738 18464 17746 18528
rect 17810 18464 17826 18528
rect 17890 18464 17906 18528
rect 17970 18464 17986 18528
rect 18050 18464 18058 18528
rect 17738 17440 18058 18464
rect 17738 17376 17746 17440
rect 17810 17376 17826 17440
rect 17890 17376 17906 17440
rect 17970 17376 17986 17440
rect 18050 17376 18058 17440
rect 17738 16352 18058 17376
rect 17738 16288 17746 16352
rect 17810 16288 17826 16352
rect 17890 16288 17906 16352
rect 17970 16288 17986 16352
rect 18050 16288 18058 16352
rect 17738 15264 18058 16288
rect 17738 15200 17746 15264
rect 17810 15200 17826 15264
rect 17890 15200 17906 15264
rect 17970 15200 17986 15264
rect 18050 15200 18058 15264
rect 16619 15196 16685 15197
rect 16619 15132 16620 15196
rect 16684 15132 16685 15196
rect 16619 15131 16685 15132
rect 14939 14656 14947 14720
rect 15011 14656 15027 14720
rect 15091 14656 15107 14720
rect 15171 14656 15187 14720
rect 15251 14656 15259 14720
rect 14939 13632 15259 14656
rect 17171 14244 17237 14245
rect 17171 14180 17172 14244
rect 17236 14180 17237 14244
rect 17171 14179 17237 14180
rect 14939 13568 14947 13632
rect 15011 13568 15027 13632
rect 15091 13568 15107 13632
rect 15171 13568 15187 13632
rect 15251 13568 15259 13632
rect 14939 12544 15259 13568
rect 14939 12480 14947 12544
rect 15011 12480 15027 12544
rect 15091 12480 15107 12544
rect 15171 12480 15187 12544
rect 15251 12480 15259 12544
rect 14939 11456 15259 12480
rect 14939 11392 14947 11456
rect 15011 11392 15027 11456
rect 15091 11392 15107 11456
rect 15171 11392 15187 11456
rect 15251 11392 15259 11456
rect 14939 10368 15259 11392
rect 14939 10304 14947 10368
rect 15011 10304 15027 10368
rect 15091 10304 15107 10368
rect 15171 10304 15187 10368
rect 15251 10304 15259 10368
rect 14939 9280 15259 10304
rect 14939 9216 14947 9280
rect 15011 9216 15027 9280
rect 15091 9216 15107 9280
rect 15171 9216 15187 9280
rect 15251 9216 15259 9280
rect 14939 8192 15259 9216
rect 16619 8396 16685 8397
rect 16619 8332 16620 8396
rect 16684 8332 16685 8396
rect 16619 8331 16685 8332
rect 14939 8128 14947 8192
rect 15011 8128 15027 8192
rect 15091 8128 15107 8192
rect 15171 8128 15187 8192
rect 15251 8128 15259 8192
rect 14939 7104 15259 8128
rect 14939 7040 14947 7104
rect 15011 7040 15027 7104
rect 15091 7040 15107 7104
rect 15171 7040 15187 7104
rect 15251 7040 15259 7104
rect 14939 6016 15259 7040
rect 14939 5952 14947 6016
rect 15011 5952 15027 6016
rect 15091 5952 15107 6016
rect 15171 5952 15187 6016
rect 15251 5952 15259 6016
rect 14939 4928 15259 5952
rect 14939 4864 14947 4928
rect 15011 4864 15027 4928
rect 15091 4864 15107 4928
rect 15171 4864 15187 4928
rect 15251 4864 15259 4928
rect 14939 3840 15259 4864
rect 16622 4045 16682 8331
rect 17174 4181 17234 14179
rect 17738 14176 18058 15200
rect 17738 14112 17746 14176
rect 17810 14112 17826 14176
rect 17890 14112 17906 14176
rect 17970 14112 17986 14176
rect 18050 14112 18058 14176
rect 17738 13088 18058 14112
rect 18278 13429 18338 21795
rect 20537 21248 20857 22272
rect 20537 21184 20545 21248
rect 20609 21184 20625 21248
rect 20689 21184 20705 21248
rect 20769 21184 20785 21248
rect 20849 21184 20857 21248
rect 20537 20160 20857 21184
rect 20537 20096 20545 20160
rect 20609 20096 20625 20160
rect 20689 20096 20705 20160
rect 20769 20096 20785 20160
rect 20849 20096 20857 20160
rect 18459 19548 18525 19549
rect 18459 19484 18460 19548
rect 18524 19484 18525 19548
rect 18459 19483 18525 19484
rect 18275 13428 18341 13429
rect 18275 13364 18276 13428
rect 18340 13364 18341 13428
rect 18275 13363 18341 13364
rect 17738 13024 17746 13088
rect 17810 13024 17826 13088
rect 17890 13024 17906 13088
rect 17970 13024 17986 13088
rect 18050 13024 18058 13088
rect 17738 12000 18058 13024
rect 18462 12341 18522 19483
rect 20537 19072 20857 20096
rect 20537 19008 20545 19072
rect 20609 19008 20625 19072
rect 20689 19008 20705 19072
rect 20769 19008 20785 19072
rect 20849 19008 20857 19072
rect 19931 18868 19997 18869
rect 19931 18804 19932 18868
rect 19996 18804 19997 18868
rect 19931 18803 19997 18804
rect 18827 12748 18893 12749
rect 18827 12684 18828 12748
rect 18892 12684 18893 12748
rect 18827 12683 18893 12684
rect 18459 12340 18525 12341
rect 18459 12276 18460 12340
rect 18524 12276 18525 12340
rect 18459 12275 18525 12276
rect 17738 11936 17746 12000
rect 17810 11936 17826 12000
rect 17890 11936 17906 12000
rect 17970 11936 17986 12000
rect 18050 11936 18058 12000
rect 17738 10912 18058 11936
rect 17738 10848 17746 10912
rect 17810 10848 17826 10912
rect 17890 10848 17906 10912
rect 17970 10848 17986 10912
rect 18050 10848 18058 10912
rect 17738 9824 18058 10848
rect 17738 9760 17746 9824
rect 17810 9760 17826 9824
rect 17890 9760 17906 9824
rect 17970 9760 17986 9824
rect 18050 9760 18058 9824
rect 17738 8736 18058 9760
rect 17738 8672 17746 8736
rect 17810 8672 17826 8736
rect 17890 8672 17906 8736
rect 17970 8672 17986 8736
rect 18050 8672 18058 8736
rect 17738 7648 18058 8672
rect 17738 7584 17746 7648
rect 17810 7584 17826 7648
rect 17890 7584 17906 7648
rect 17970 7584 17986 7648
rect 18050 7584 18058 7648
rect 17738 6560 18058 7584
rect 18643 7036 18709 7037
rect 18643 6972 18644 7036
rect 18708 6972 18709 7036
rect 18643 6971 18709 6972
rect 17738 6496 17746 6560
rect 17810 6496 17826 6560
rect 17890 6496 17906 6560
rect 17970 6496 17986 6560
rect 18050 6496 18058 6560
rect 17738 5472 18058 6496
rect 18646 5949 18706 6971
rect 18643 5948 18709 5949
rect 18643 5884 18644 5948
rect 18708 5884 18709 5948
rect 18643 5883 18709 5884
rect 17738 5408 17746 5472
rect 17810 5408 17826 5472
rect 17890 5408 17906 5472
rect 17970 5408 17986 5472
rect 18050 5408 18058 5472
rect 17738 4384 18058 5408
rect 18830 5133 18890 12683
rect 19934 12450 19994 18803
rect 20537 17984 20857 19008
rect 20537 17920 20545 17984
rect 20609 17920 20625 17984
rect 20689 17920 20705 17984
rect 20769 17920 20785 17984
rect 20849 17920 20857 17984
rect 20537 16896 20857 17920
rect 20537 16832 20545 16896
rect 20609 16832 20625 16896
rect 20689 16832 20705 16896
rect 20769 16832 20785 16896
rect 20849 16832 20857 16896
rect 20537 15808 20857 16832
rect 20537 15744 20545 15808
rect 20609 15744 20625 15808
rect 20689 15744 20705 15808
rect 20769 15744 20785 15808
rect 20849 15744 20857 15808
rect 20537 14720 20857 15744
rect 20537 14656 20545 14720
rect 20609 14656 20625 14720
rect 20689 14656 20705 14720
rect 20769 14656 20785 14720
rect 20849 14656 20857 14720
rect 20537 13632 20857 14656
rect 20537 13568 20545 13632
rect 20609 13568 20625 13632
rect 20689 13568 20705 13632
rect 20769 13568 20785 13632
rect 20849 13568 20857 13632
rect 20537 12544 20857 13568
rect 20537 12480 20545 12544
rect 20609 12480 20625 12544
rect 20689 12480 20705 12544
rect 20769 12480 20785 12544
rect 20849 12480 20857 12544
rect 19934 12390 20362 12450
rect 19195 11252 19261 11253
rect 19195 11188 19196 11252
rect 19260 11188 19261 11252
rect 19195 11187 19261 11188
rect 19011 8804 19077 8805
rect 19011 8740 19012 8804
rect 19076 8740 19077 8804
rect 19011 8739 19077 8740
rect 18827 5132 18893 5133
rect 18827 5068 18828 5132
rect 18892 5068 18893 5132
rect 18827 5067 18893 5068
rect 19014 4589 19074 8739
rect 19198 4725 19258 11187
rect 20302 7853 20362 12390
rect 20537 11456 20857 12480
rect 20537 11392 20545 11456
rect 20609 11392 20625 11456
rect 20689 11392 20705 11456
rect 20769 11392 20785 11456
rect 20849 11392 20857 11456
rect 20537 10368 20857 11392
rect 20537 10304 20545 10368
rect 20609 10304 20625 10368
rect 20689 10304 20705 10368
rect 20769 10304 20785 10368
rect 20849 10304 20857 10368
rect 20537 9280 20857 10304
rect 20537 9216 20545 9280
rect 20609 9216 20625 9280
rect 20689 9216 20705 9280
rect 20769 9216 20785 9280
rect 20849 9216 20857 9280
rect 20537 8192 20857 9216
rect 20537 8128 20545 8192
rect 20609 8128 20625 8192
rect 20689 8128 20705 8192
rect 20769 8128 20785 8192
rect 20849 8128 20857 8192
rect 20299 7852 20365 7853
rect 20299 7788 20300 7852
rect 20364 7788 20365 7852
rect 20299 7787 20365 7788
rect 20302 6493 20362 7787
rect 20537 7104 20857 8128
rect 21035 7716 21101 7717
rect 21035 7652 21036 7716
rect 21100 7652 21101 7716
rect 21035 7651 21101 7652
rect 20537 7040 20545 7104
rect 20609 7040 20625 7104
rect 20689 7040 20705 7104
rect 20769 7040 20785 7104
rect 20849 7040 20857 7104
rect 20299 6492 20365 6493
rect 20299 6428 20300 6492
rect 20364 6428 20365 6492
rect 20299 6427 20365 6428
rect 20537 6016 20857 7040
rect 20537 5952 20545 6016
rect 20609 5952 20625 6016
rect 20689 5952 20705 6016
rect 20769 5952 20785 6016
rect 20849 5952 20857 6016
rect 20537 4928 20857 5952
rect 20537 4864 20545 4928
rect 20609 4864 20625 4928
rect 20689 4864 20705 4928
rect 20769 4864 20785 4928
rect 20849 4864 20857 4928
rect 19195 4724 19261 4725
rect 19195 4660 19196 4724
rect 19260 4660 19261 4724
rect 19195 4659 19261 4660
rect 19011 4588 19077 4589
rect 19011 4524 19012 4588
rect 19076 4524 19077 4588
rect 19011 4523 19077 4524
rect 17738 4320 17746 4384
rect 17810 4320 17826 4384
rect 17890 4320 17906 4384
rect 17970 4320 17986 4384
rect 18050 4320 18058 4384
rect 17171 4180 17237 4181
rect 17171 4116 17172 4180
rect 17236 4116 17237 4180
rect 17171 4115 17237 4116
rect 16619 4044 16685 4045
rect 16619 3980 16620 4044
rect 16684 3980 16685 4044
rect 16619 3979 16685 3980
rect 14939 3776 14947 3840
rect 15011 3776 15027 3840
rect 15091 3776 15107 3840
rect 15171 3776 15187 3840
rect 15251 3776 15259 3840
rect 14939 2752 15259 3776
rect 14939 2688 14947 2752
rect 15011 2688 15027 2752
rect 15091 2688 15107 2752
rect 15171 2688 15187 2752
rect 15251 2688 15259 2752
rect 14939 2128 15259 2688
rect 17738 3296 18058 4320
rect 17738 3232 17746 3296
rect 17810 3232 17826 3296
rect 17890 3232 17906 3296
rect 17970 3232 17986 3296
rect 18050 3232 18058 3296
rect 17738 2208 18058 3232
rect 17738 2144 17746 2208
rect 17810 2144 17826 2208
rect 17890 2144 17906 2208
rect 17970 2144 17986 2208
rect 18050 2144 18058 2208
rect 17738 2128 18058 2144
rect 20537 3840 20857 4864
rect 20537 3776 20545 3840
rect 20609 3776 20625 3840
rect 20689 3776 20705 3840
rect 20769 3776 20785 3840
rect 20849 3776 20857 3840
rect 20537 2752 20857 3776
rect 21038 3773 21098 7651
rect 21403 7172 21469 7173
rect 21403 7108 21404 7172
rect 21468 7108 21469 7172
rect 21403 7107 21469 7108
rect 21406 6357 21466 7107
rect 22139 7036 22205 7037
rect 22139 6972 22140 7036
rect 22204 6972 22205 7036
rect 22139 6971 22205 6972
rect 21403 6356 21469 6357
rect 21403 6292 21404 6356
rect 21468 6292 21469 6356
rect 21403 6291 21469 6292
rect 22142 5949 22202 6971
rect 22139 5948 22205 5949
rect 22139 5884 22140 5948
rect 22204 5884 22205 5948
rect 22139 5883 22205 5884
rect 21035 3772 21101 3773
rect 21035 3708 21036 3772
rect 21100 3708 21101 3772
rect 21035 3707 21101 3708
rect 20537 2688 20545 2752
rect 20609 2688 20625 2752
rect 20689 2688 20705 2752
rect 20769 2688 20785 2752
rect 20849 2688 20857 2752
rect 20537 2128 20857 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_FTB00_A
timestamp 1649977179
transform 1 0 10948 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform -1 0 10856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 16560 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 16192 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform 1 0 14536 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform -1 0 2576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform -1 0 2116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform -1 0 2300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform -1 0 2944 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform -1 0 3128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1649977179
transform -1 0 2852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1649977179
transform -1 0 2484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1649977179
transform -1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 23184 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 17940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 13984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 12328 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 12880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 23184 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 23184 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 2668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 11316 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 10304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 5428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 3036 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 3312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform 1 0 16008 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 3220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 2300 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 3404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 2852 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 2944 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 5980 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6624 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7820 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9476 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11868 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1649977179
transform -1 0 6532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 9568 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 5520 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12052 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5244 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 5060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 8096 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 14168 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 2576 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 9108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 10580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15824 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 18032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 17848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 23000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 23000 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 23000 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14536 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14168 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 4692 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1649977179
transform -1 0 16100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 8556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 8464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 10948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 7360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf_A
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 9568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 23000 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 17756 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1649977179
transform -1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1649977179
transform -1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16192 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 23000 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 14352 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 15364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 23000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 10948 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 14352 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 11960 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 13432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 23000 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output38_A
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output50_A
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1649977179
transform -1 0 19596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 1649977179
transform -1 0 19964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1649977179
transform -1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1649977179
transform -1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1649977179
transform -1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1649977179
transform -1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform -1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform -1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1649977179
transform -1 0 11408 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform -1 0 13432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1649977179
transform -1 0 15088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_E_FTB01_A
timestamp 1649977179
transform -1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 22632 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1649977179
transform -1 0 12972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater98_A
timestamp 1649977179
transform -1 0 14628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater99_A
timestamp 1649977179
transform -1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater102_A
timestamp 1649977179
transform -1 0 3680 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater104_A
timestamp 1649977179
transform -1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60
timestamp 1649977179
transform 1 0 6624 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_62
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_74
timestamp 1649977179
transform 1 0 7912 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_86
timestamp 1649977179
transform 1 0 9016 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_98
timestamp 1649977179
transform 1 0 10120 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_196
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_216
timestamp 1649977179
transform 1 0 20976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_228
timestamp 1649977179
transform 1 0 22080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_235
timestamp 1649977179
transform 1 0 22724 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_65
timestamp 1649977179
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_68
timestamp 1649977179
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_92
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_100
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_104
timestamp 1649977179
transform 1 0 10672 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1649977179
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_102
timestamp 1649977179
transform 1 0 10488 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_114
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_126
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_92
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1649977179
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 1649977179
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_190
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_239
timestamp 1649977179
transform 1 0 23092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_70
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1649977179
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_113
timestamp 1649977179
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_119
timestamp 1649977179
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_123
timestamp 1649977179
transform 1 0 12420 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_171
timestamp 1649977179
transform 1 0 16836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_12
timestamp 1649977179
transform 1 0 2208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_186
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_239
timestamp 1649977179
transform 1 0 23092 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_79
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp 1649977179
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_123
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_36
timestamp 1649977179
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_49
timestamp 1649977179
transform 1 0 5612 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_55
timestamp 1649977179
transform 1 0 6164 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_74
timestamp 1649977179
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1649977179
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_20
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_96
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1649977179
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_105
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1649977179
transform 1 0 12420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 1649977179
transform 1 0 10304 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_239
timestamp 1649977179
transform 1 0 23092 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_117
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 1649977179
transform 1 0 3036 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_80
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_92
timestamp 1649977179
transform 1 0 9568 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_149
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_186
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_45
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1649977179
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_165
timestamp 1649977179
transform 1 0 16284 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1649977179
transform 1 0 3220 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_47
timestamp 1649977179
transform 1 0 5428 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_75
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_124
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1649977179
transform 1 0 13064 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_143
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_13
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_25
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_37
timestamp 1649977179
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_130
timestamp 1649977179
transform 1 0 13064 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_226
timestamp 1649977179
transform 1 0 21896 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_44
timestamp 1649977179
transform 1 0 5152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_78
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_88
timestamp 1649977179
transform 1 0 9200 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_122
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1649977179
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1649977179
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_107
timestamp 1649977179
transform 1 0 10948 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_164
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_36
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_132
timestamp 1649977179
transform 1 0 13248 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_32
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_111
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_173
timestamp 1649977179
transform 1 0 17020 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_75
timestamp 1649977179
transform 1 0 8004 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_191
timestamp 1649977179
transform 1 0 18676 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_129
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1649977179
transform 1 0 3220 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_34
timestamp 1649977179
transform 1 0 4232 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_120
timestamp 1649977179
transform 1 0 12144 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_127
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_222
timestamp 1649977179
transform 1 0 21528 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_11
timestamp 1649977179
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_16
timestamp 1649977179
transform 1 0 2576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_44
timestamp 1649977179
transform 1 0 5152 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_73
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_152
timestamp 1649977179
transform 1 0 15088 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_231
timestamp 1649977179
transform 1 0 22356 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_22
timestamp 1649977179
transform 1 0 3128 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_10
timestamp 1649977179
transform 1 0 2024 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1649977179
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 1649977179
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_113
timestamp 1649977179
transform 1 0 11500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 23460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 23460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 23460 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 23460 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 23460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 23460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 23460 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 23460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 23460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 23460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 23460 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 23460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 23460 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 23460 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 23460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 23460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  Test_en_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_W_FTB01
timestamp 1649977179
transform 1 0 1840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 13432 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 23000 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 16744 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 16560 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform -1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform -1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 2392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform 1 0 3220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform 1 0 3496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform -1 0 4048 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform -1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  clk_0_FTB00
timestamp 1649977179
transform -1 0 15088 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  grid_clb_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1649977179
transform -1 0 18400 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1649977179
transform -1 0 21712 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1649977179
transform -1 0 17388 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1649977179
transform -1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1649977179
transform -1 0 16652 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 18400 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 18400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 19136 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 22080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 22908 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 18676 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 18676 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 9016 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 11408 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 13156 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 13616 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 4876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 16192 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 5704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 6532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 10396 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12972 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5060 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3864 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 3588 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 4784 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 4600 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4784 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4508 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 3680 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 3956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 3956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 5152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 4508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 6992 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4416 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform -1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 7176 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 7728 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 7084 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 8280 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 8280 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 14996 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform -1 0 8188 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6624 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4876 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9016 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__127
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11040 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16100 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9016 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9476 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__128
timestamp 1649977179
transform -1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8648 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__129
timestamp 1649977179
transform -1 0 8188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11592 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__130
timestamp 1649977179
transform 1 0 12512 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 9476 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5704 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 4784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform -1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4508 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 4416 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 5428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 7176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 4968 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 4416 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform -1 0 4140 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6808 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8004 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6624 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 10856 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 10304 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 8832 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform -1 0 8280 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 7084 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 8648 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 9568 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 11408 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 8372 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform -1 0 7360 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3496 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__131
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6072 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14628 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7912 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6992 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__132
timestamp 1649977179
transform -1 0 6256 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6900 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11132 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__133
timestamp 1649977179
transform -1 0 11408 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__134
timestamp 1649977179
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 12696 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4048 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8464 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 8372 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 9200 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 3680 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 4876 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4416 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3588 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5152 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 15456 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 15732 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 12512 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 22172 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 4692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 4232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 7820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 13892 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 12420 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform 1 0 4692 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7176 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5888 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 15548 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 13984 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 13064 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 11132 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 6256 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 7636 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 9108 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13984 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__135
timestamp 1649977179
transform 1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13984 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11684 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14812 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17020 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15732 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__136
timestamp 1649977179
transform 1 0 18400 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18308 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__137
timestamp 1649977179
transform -1 0 17388 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14260 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13432 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__106
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 18216 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 19136 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13156 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13340 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14904 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 16560 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16008 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 17112 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 17204 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16468 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 17480 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 17940 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 15732 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 16192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 16008 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 16376 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 17480 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform -1 0 13156 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15824 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13064 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11132 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 18676 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 18400 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 18216 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 17020 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 18124 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 18492 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 20240 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19136 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21528 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__107
timestamp 1649977179
transform -1 0 18400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17664 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20148 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18768 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 22172 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19596 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20976 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20884 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__108
timestamp 1649977179
transform -1 0 16560 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20608 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20884 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__109
timestamp 1649977179
transform -1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20700 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__110
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 5888 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 10212 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9016 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7176 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7636 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10488 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 10672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23000 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7360 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5888 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6808 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 9752 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 4416 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 12972 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 9936 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 12880 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13616 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13064 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__111
timestamp 1649977179
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18492 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 22172 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16284 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16100 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19136 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__112
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20148 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18584 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__114
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15088 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 13156 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12420 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 11132 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 18216 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20148 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 20240 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform 1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23000 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 21160 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform -1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11684 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14904 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13156 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 13432 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 11868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 12052 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform -1 0 12328 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 11776 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 17112 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 16468 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18492 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18308 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__115
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17480 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14536 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20424 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14628 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16836 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__116
timestamp 1649977179
transform -1 0 16560 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19136 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20700 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__117
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13984 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__118
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 17204 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21620 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 21528 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 22632 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 22356 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 21528 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 22632 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform -1 0 21528 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21528 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 21528 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 22356 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform 1 0 22356 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform 1 0 22356 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 22172 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 21712 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 19136 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 18676 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 18584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 23092 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12144 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16192 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 13248 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 14904 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 18584 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 21620 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 20700 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 18676 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 21620 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 18676 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 19688 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 20056 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 22172 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__119
timestamp 1649977179
transform -1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 22172 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20148 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19596 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17756 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21712 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__120
timestamp 1649977179
transform -1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20884 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 22080 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__121
timestamp 1649977179
transform -1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__122
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22540 0 1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21528 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 22448 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 21068 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 21528 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform -1 0 21436 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 22172 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform -1 0 21068 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 22632 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 22632 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 22816 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 22724 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 22632 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 22724 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 22724 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 21712 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform 1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 13984 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 21804 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 19136 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 22448 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.delay_buf
timestamp 1649977179
transform -1 0 11500 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17020 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14720 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 20700 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 18308 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 21068 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 20700 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 20148 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 18216 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21068 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 22080 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21988 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__123
timestamp 1649977179
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20332 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21896 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__124
timestamp 1649977179
transform -1 0 19136 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20884 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__125
timestamp 1649977179
transform -1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__126
timestamp 1649977179
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output38 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform 1 0 20976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 21712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1649977179
transform -1 0 17112 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1649977179
transform -1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1649977179
transform -1 0 22448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform 1 0 22448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform 1 0 22816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 22448 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 22816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 22724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 22816 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 22080 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 2116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 2024 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 22448 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 4140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23184 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1649977179
transform -1 0 19136 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform -1 0 22724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1649977179
transform -1 0 18216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  repeater80
timestamp 1649977179
transform -1 0 21528 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater81
timestamp 1649977179
transform -1 0 23000 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater82
timestamp 1649977179
transform -1 0 21528 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater83 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21620 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater84
timestamp 1649977179
transform -1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater85
timestamp 1649977179
transform -1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater86
timestamp 1649977179
transform -1 0 11316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater87
timestamp 1649977179
transform -1 0 11408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater88
timestamp 1649977179
transform -1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater89
timestamp 1649977179
transform -1 0 16560 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater90
timestamp 1649977179
transform 1 0 5704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater91
timestamp 1649977179
transform -1 0 5520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater92
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater93
timestamp 1649977179
transform 1 0 5336 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater94
timestamp 1649977179
transform -1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater95
timestamp 1649977179
transform 1 0 4784 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater96
timestamp 1649977179
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater97
timestamp 1649977179
transform -1 0 16468 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater98
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater99
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater100
timestamp 1649977179
transform -1 0 15456 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater101
timestamp 1649977179
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater102
timestamp 1649977179
transform -1 0 10672 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater103
timestamp 1649977179
transform 1 0 16836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater104
timestamp 1649977179
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
<< labels >>
flabel metal2 s 17038 23800 17094 24600 0 FreeSans 224 90 0 0 SC_IN_TOP
port 0 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal2 s 17682 23800 17738 24600 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 2 nsew signal tristate
flabel metal3 s 23800 7896 24600 8016 0 FreeSans 480 0 0 0 Test_en_E_in
port 3 nsew signal input
flabel metal3 s 23800 7352 24600 7472 0 FreeSans 480 0 0 0 Test_en_E_out
port 4 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 Test_en_W_in
port 5 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 Test_en_W_out
port 6 nsew signal tristate
flabel metal4 s 6542 2128 6862 22352 0 FreeSans 1920 90 0 0 VGND
port 7 nsew ground bidirectional
flabel metal4 s 12140 2128 12460 22352 0 FreeSans 1920 90 0 0 VGND
port 7 nsew ground bidirectional
flabel metal4 s 17738 2128 18058 22352 0 FreeSans 1920 90 0 0 VGND
port 7 nsew ground bidirectional
flabel metal4 s 3743 2128 4063 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal4 s 9341 2128 9661 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal4 s 14939 2128 15259 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal4 s 20537 2128 20857 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_50_
port 9 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_51_
port 10 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 ccff_head
port 11 nsew signal input
flabel metal3 s 23800 6808 24600 6928 0 FreeSans 480 0 0 0 ccff_tail
port 12 nsew signal tristate
flabel metal2 s 18326 23800 18382 24600 0 FreeSans 224 90 0 0 clk_0_N_in
port 13 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 clk_0_S_in
port 14 nsew signal input
flabel metal3 s 23800 8984 24600 9104 0 FreeSans 480 0 0 0 prog_clk_0_E_out
port 15 nsew signal tristate
flabel metal3 s 23800 8440 24600 8560 0 FreeSans 480 0 0 0 prog_clk_0_N_in
port 16 nsew signal input
flabel metal2 s 18970 23800 19026 24600 0 FreeSans 224 90 0 0 prog_clk_0_N_out
port 17 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 18 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 prog_clk_0_S_out
port 19 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 prog_clk_0_W_out
port 20 nsew signal tristate
flabel metal3 s 23800 9528 24600 9648 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_16_
port 21 nsew signal input
flabel metal3 s 23800 10072 24600 10192 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_17_
port 22 nsew signal input
flabel metal3 s 23800 10616 24600 10736 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_18_
port 23 nsew signal input
flabel metal3 s 23800 11160 24600 11280 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_19_
port 24 nsew signal input
flabel metal3 s 23800 11704 24600 11824 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_20_
port 25 nsew signal input
flabel metal3 s 23800 12248 24600 12368 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_21_
port 26 nsew signal input
flabel metal3 s 23800 12792 24600 12912 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_22_
port 27 nsew signal input
flabel metal3 s 23800 13336 24600 13456 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_23_
port 28 nsew signal input
flabel metal3 s 23800 13880 24600 14000 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_24_
port 29 nsew signal input
flabel metal3 s 23800 14424 24600 14544 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_25_
port 30 nsew signal input
flabel metal3 s 23800 14968 24600 15088 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_26_
port 31 nsew signal input
flabel metal3 s 23800 15512 24600 15632 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_27_
port 32 nsew signal input
flabel metal3 s 23800 16056 24600 16176 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_28_
port 33 nsew signal input
flabel metal3 s 23800 16600 24600 16720 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_29_
port 34 nsew signal input
flabel metal3 s 23800 17144 24600 17264 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_30_
port 35 nsew signal input
flabel metal3 s 23800 17688 24600 17808 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_31_
port 36 nsew signal input
flabel metal3 s 23800 2456 24600 2576 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_42_lower
port 37 nsew signal tristate
flabel metal3 s 23800 18232 24600 18352 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_42_upper
port 38 nsew signal tristate
flabel metal3 s 23800 3000 24600 3120 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_43_lower
port 39 nsew signal tristate
flabel metal3 s 23800 18776 24600 18896 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_43_upper
port 40 nsew signal tristate
flabel metal3 s 23800 3544 24600 3664 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_44_lower
port 41 nsew signal tristate
flabel metal3 s 23800 19320 24600 19440 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_44_upper
port 42 nsew signal tristate
flabel metal3 s 23800 4088 24600 4208 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_45_lower
port 43 nsew signal tristate
flabel metal3 s 23800 19864 24600 19984 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_45_upper
port 44 nsew signal tristate
flabel metal3 s 23800 4632 24600 4752 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_46_lower
port 45 nsew signal tristate
flabel metal3 s 23800 20408 24600 20528 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_46_upper
port 46 nsew signal tristate
flabel metal3 s 23800 5176 24600 5296 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_47_lower
port 47 nsew signal tristate
flabel metal3 s 23800 20952 24600 21072 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_47_upper
port 48 nsew signal tristate
flabel metal3 s 23800 5720 24600 5840 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_48_lower
port 49 nsew signal tristate
flabel metal3 s 23800 21496 24600 21616 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_48_upper
port 50 nsew signal tristate
flabel metal3 s 23800 6264 24600 6384 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_49_lower
port 51 nsew signal tristate
flabel metal3 s 23800 22040 24600 22160 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_49_upper
port 52 nsew signal tristate
flabel metal2 s 5446 23800 5502 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_0_
port 53 nsew signal input
flabel metal2 s 11886 23800 11942 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_10_
port 54 nsew signal input
flabel metal2 s 12530 23800 12586 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_11_
port 55 nsew signal input
flabel metal2 s 13174 23800 13230 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_12_
port 56 nsew signal input
flabel metal2 s 13818 23800 13874 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_13_
port 57 nsew signal input
flabel metal2 s 14462 23800 14518 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_14_
port 58 nsew signal input
flabel metal2 s 15106 23800 15162 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_15_
port 59 nsew signal input
flabel metal2 s 6090 23800 6146 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_1_
port 60 nsew signal input
flabel metal2 s 6734 23800 6790 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_2_
port 61 nsew signal input
flabel metal2 s 15750 23800 15806 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_32_
port 62 nsew signal input
flabel metal2 s 16394 23800 16450 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_33_
port 63 nsew signal input
flabel metal2 s 19614 23800 19670 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_34_lower
port 64 nsew signal tristate
flabel metal2 s 294 23800 350 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_34_upper
port 65 nsew signal tristate
flabel metal2 s 20258 23800 20314 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_35_lower
port 66 nsew signal tristate
flabel metal2 s 938 23800 994 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_35_upper
port 67 nsew signal tristate
flabel metal2 s 20902 23800 20958 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_36_lower
port 68 nsew signal tristate
flabel metal2 s 1582 23800 1638 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_36_upper
port 69 nsew signal tristate
flabel metal2 s 21546 23800 21602 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_37_lower
port 70 nsew signal tristate
flabel metal2 s 2226 23800 2282 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_37_upper
port 71 nsew signal tristate
flabel metal2 s 22190 23800 22246 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_38_lower
port 72 nsew signal tristate
flabel metal2 s 2870 23800 2926 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_38_upper
port 73 nsew signal tristate
flabel metal2 s 22834 23800 22890 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_39_lower
port 74 nsew signal tristate
flabel metal2 s 3514 23800 3570 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_39_upper
port 75 nsew signal tristate
flabel metal2 s 7378 23800 7434 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_3_
port 76 nsew signal input
flabel metal2 s 23478 23800 23534 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_40_lower
port 77 nsew signal tristate
flabel metal2 s 4158 23800 4214 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_40_upper
port 78 nsew signal tristate
flabel metal2 s 24122 23800 24178 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_41_lower
port 79 nsew signal tristate
flabel metal2 s 4802 23800 4858 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_41_upper
port 80 nsew signal tristate
flabel metal2 s 8022 23800 8078 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_4_
port 81 nsew signal input
flabel metal2 s 8666 23800 8722 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_5_
port 82 nsew signal input
flabel metal2 s 9310 23800 9366 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_6_
port 83 nsew signal input
flabel metal2 s 9954 23800 10010 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_7_
port 84 nsew signal input
flabel metal2 s 10598 23800 10654 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_8_
port 85 nsew signal input
flabel metal2 s 11242 23800 11298 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_9_
port 86 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 24600 24600
<< end >>
